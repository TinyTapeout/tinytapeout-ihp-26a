module tt_um_SotaSoC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire \soc_inst.bus_spi_sclk ;
 wire \soc_inst.core_instr_addr[0] ;
 wire \soc_inst.core_instr_addr[10] ;
 wire \soc_inst.core_instr_addr[11] ;
 wire \soc_inst.core_instr_addr[12] ;
 wire \soc_inst.core_instr_addr[13] ;
 wire \soc_inst.core_instr_addr[14] ;
 wire \soc_inst.core_instr_addr[15] ;
 wire \soc_inst.core_instr_addr[16] ;
 wire \soc_inst.core_instr_addr[17] ;
 wire \soc_inst.core_instr_addr[18] ;
 wire \soc_inst.core_instr_addr[19] ;
 wire \soc_inst.core_instr_addr[1] ;
 wire \soc_inst.core_instr_addr[20] ;
 wire \soc_inst.core_instr_addr[21] ;
 wire \soc_inst.core_instr_addr[22] ;
 wire \soc_inst.core_instr_addr[23] ;
 wire \soc_inst.core_instr_addr[2] ;
 wire \soc_inst.core_instr_addr[3] ;
 wire \soc_inst.core_instr_addr[4] ;
 wire \soc_inst.core_instr_addr[5] ;
 wire \soc_inst.core_instr_addr[6] ;
 wire \soc_inst.core_instr_addr[7] ;
 wire \soc_inst.core_instr_addr[8] ;
 wire \soc_inst.core_instr_addr[9] ;
 wire \soc_inst.core_instr_data[0] ;
 wire \soc_inst.core_instr_data[10] ;
 wire \soc_inst.core_instr_data[11] ;
 wire \soc_inst.core_instr_data[12] ;
 wire \soc_inst.core_instr_data[13] ;
 wire \soc_inst.core_instr_data[14] ;
 wire \soc_inst.core_instr_data[15] ;
 wire \soc_inst.core_instr_data[16] ;
 wire \soc_inst.core_instr_data[17] ;
 wire \soc_inst.core_instr_data[18] ;
 wire \soc_inst.core_instr_data[19] ;
 wire \soc_inst.core_instr_data[1] ;
 wire \soc_inst.core_instr_data[20] ;
 wire \soc_inst.core_instr_data[21] ;
 wire \soc_inst.core_instr_data[22] ;
 wire \soc_inst.core_instr_data[23] ;
 wire \soc_inst.core_instr_data[24] ;
 wire \soc_inst.core_instr_data[25] ;
 wire \soc_inst.core_instr_data[26] ;
 wire \soc_inst.core_instr_data[27] ;
 wire \soc_inst.core_instr_data[28] ;
 wire \soc_inst.core_instr_data[29] ;
 wire \soc_inst.core_instr_data[2] ;
 wire \soc_inst.core_instr_data[30] ;
 wire \soc_inst.core_instr_data[31] ;
 wire \soc_inst.core_instr_data[3] ;
 wire \soc_inst.core_instr_data[4] ;
 wire \soc_inst.core_instr_data[5] ;
 wire \soc_inst.core_instr_data[6] ;
 wire \soc_inst.core_instr_data[7] ;
 wire \soc_inst.core_instr_data[8] ;
 wire \soc_inst.core_instr_data[9] ;
 wire \soc_inst.core_mem_addr[0] ;
 wire \soc_inst.core_mem_addr[10] ;
 wire \soc_inst.core_mem_addr[11] ;
 wire \soc_inst.core_mem_addr[12] ;
 wire \soc_inst.core_mem_addr[13] ;
 wire \soc_inst.core_mem_addr[14] ;
 wire \soc_inst.core_mem_addr[15] ;
 wire \soc_inst.core_mem_addr[16] ;
 wire \soc_inst.core_mem_addr[17] ;
 wire \soc_inst.core_mem_addr[18] ;
 wire \soc_inst.core_mem_addr[19] ;
 wire \soc_inst.core_mem_addr[1] ;
 wire \soc_inst.core_mem_addr[20] ;
 wire \soc_inst.core_mem_addr[21] ;
 wire \soc_inst.core_mem_addr[22] ;
 wire \soc_inst.core_mem_addr[23] ;
 wire \soc_inst.core_mem_addr[24] ;
 wire \soc_inst.core_mem_addr[25] ;
 wire \soc_inst.core_mem_addr[26] ;
 wire \soc_inst.core_mem_addr[27] ;
 wire \soc_inst.core_mem_addr[28] ;
 wire \soc_inst.core_mem_addr[29] ;
 wire \soc_inst.core_mem_addr[2] ;
 wire \soc_inst.core_mem_addr[30] ;
 wire \soc_inst.core_mem_addr[31] ;
 wire \soc_inst.core_mem_addr[3] ;
 wire \soc_inst.core_mem_addr[5] ;
 wire \soc_inst.core_mem_addr[6] ;
 wire \soc_inst.core_mem_addr[7] ;
 wire \soc_inst.core_mem_addr[8] ;
 wire \soc_inst.core_mem_addr[9] ;
 wire \soc_inst.core_mem_flag[0] ;
 wire \soc_inst.core_mem_flag[1] ;
 wire \soc_inst.core_mem_flag[2] ;
 wire \soc_inst.core_mem_rdata[0] ;
 wire \soc_inst.core_mem_rdata[10] ;
 wire \soc_inst.core_mem_rdata[11] ;
 wire \soc_inst.core_mem_rdata[12] ;
 wire \soc_inst.core_mem_rdata[13] ;
 wire \soc_inst.core_mem_rdata[14] ;
 wire \soc_inst.core_mem_rdata[15] ;
 wire \soc_inst.core_mem_rdata[16] ;
 wire \soc_inst.core_mem_rdata[17] ;
 wire \soc_inst.core_mem_rdata[18] ;
 wire \soc_inst.core_mem_rdata[19] ;
 wire \soc_inst.core_mem_rdata[1] ;
 wire \soc_inst.core_mem_rdata[20] ;
 wire \soc_inst.core_mem_rdata[21] ;
 wire \soc_inst.core_mem_rdata[22] ;
 wire \soc_inst.core_mem_rdata[23] ;
 wire \soc_inst.core_mem_rdata[24] ;
 wire \soc_inst.core_mem_rdata[25] ;
 wire \soc_inst.core_mem_rdata[26] ;
 wire \soc_inst.core_mem_rdata[27] ;
 wire \soc_inst.core_mem_rdata[28] ;
 wire \soc_inst.core_mem_rdata[29] ;
 wire \soc_inst.core_mem_rdata[2] ;
 wire \soc_inst.core_mem_rdata[30] ;
 wire \soc_inst.core_mem_rdata[31] ;
 wire \soc_inst.core_mem_rdata[3] ;
 wire \soc_inst.core_mem_rdata[4] ;
 wire \soc_inst.core_mem_rdata[5] ;
 wire \soc_inst.core_mem_rdata[6] ;
 wire \soc_inst.core_mem_rdata[7] ;
 wire \soc_inst.core_mem_rdata[8] ;
 wire \soc_inst.core_mem_rdata[9] ;
 wire \soc_inst.core_mem_re ;
 wire \soc_inst.core_mem_wdata[0] ;
 wire \soc_inst.core_mem_wdata[10] ;
 wire \soc_inst.core_mem_wdata[11] ;
 wire \soc_inst.core_mem_wdata[12] ;
 wire \soc_inst.core_mem_wdata[13] ;
 wire \soc_inst.core_mem_wdata[14] ;
 wire \soc_inst.core_mem_wdata[15] ;
 wire \soc_inst.core_mem_wdata[16] ;
 wire \soc_inst.core_mem_wdata[17] ;
 wire \soc_inst.core_mem_wdata[18] ;
 wire \soc_inst.core_mem_wdata[19] ;
 wire \soc_inst.core_mem_wdata[1] ;
 wire \soc_inst.core_mem_wdata[20] ;
 wire \soc_inst.core_mem_wdata[21] ;
 wire \soc_inst.core_mem_wdata[22] ;
 wire \soc_inst.core_mem_wdata[23] ;
 wire \soc_inst.core_mem_wdata[24] ;
 wire \soc_inst.core_mem_wdata[25] ;
 wire \soc_inst.core_mem_wdata[26] ;
 wire \soc_inst.core_mem_wdata[27] ;
 wire \soc_inst.core_mem_wdata[28] ;
 wire \soc_inst.core_mem_wdata[29] ;
 wire \soc_inst.core_mem_wdata[2] ;
 wire \soc_inst.core_mem_wdata[30] ;
 wire \soc_inst.core_mem_wdata[31] ;
 wire \soc_inst.core_mem_wdata[3] ;
 wire \soc_inst.core_mem_wdata[4] ;
 wire \soc_inst.core_mem_wdata[5] ;
 wire \soc_inst.core_mem_wdata[6] ;
 wire \soc_inst.core_mem_wdata[7] ;
 wire \soc_inst.core_mem_wdata[8] ;
 wire \soc_inst.core_mem_wdata[9] ;
 wire \soc_inst.core_mem_we ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[0] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[1] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[2] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[3] ;
 wire \soc_inst.cpu_core.alu.a[0] ;
 wire \soc_inst.cpu_core.alu.a[10] ;
 wire \soc_inst.cpu_core.alu.a[11] ;
 wire \soc_inst.cpu_core.alu.a[12] ;
 wire \soc_inst.cpu_core.alu.a[13] ;
 wire \soc_inst.cpu_core.alu.a[14] ;
 wire \soc_inst.cpu_core.alu.a[15] ;
 wire \soc_inst.cpu_core.alu.a[16] ;
 wire \soc_inst.cpu_core.alu.a[17] ;
 wire \soc_inst.cpu_core.alu.a[18] ;
 wire \soc_inst.cpu_core.alu.a[19] ;
 wire \soc_inst.cpu_core.alu.a[1] ;
 wire \soc_inst.cpu_core.alu.a[20] ;
 wire \soc_inst.cpu_core.alu.a[21] ;
 wire \soc_inst.cpu_core.alu.a[22] ;
 wire \soc_inst.cpu_core.alu.a[23] ;
 wire \soc_inst.cpu_core.alu.a[24] ;
 wire \soc_inst.cpu_core.alu.a[25] ;
 wire \soc_inst.cpu_core.alu.a[26] ;
 wire \soc_inst.cpu_core.alu.a[27] ;
 wire \soc_inst.cpu_core.alu.a[28] ;
 wire \soc_inst.cpu_core.alu.a[29] ;
 wire \soc_inst.cpu_core.alu.a[2] ;
 wire \soc_inst.cpu_core.alu.a[30] ;
 wire \soc_inst.cpu_core.alu.a[31] ;
 wire \soc_inst.cpu_core.alu.a[3] ;
 wire \soc_inst.cpu_core.alu.a[4] ;
 wire \soc_inst.cpu_core.alu.a[5] ;
 wire \soc_inst.cpu_core.alu.a[6] ;
 wire \soc_inst.cpu_core.alu.a[7] ;
 wire \soc_inst.cpu_core.alu.a[8] ;
 wire \soc_inst.cpu_core.alu.a[9] ;
 wire \soc_inst.cpu_core.alu.b[0] ;
 wire \soc_inst.cpu_core.alu.b[10] ;
 wire \soc_inst.cpu_core.alu.b[11] ;
 wire \soc_inst.cpu_core.alu.b[12] ;
 wire \soc_inst.cpu_core.alu.b[13] ;
 wire \soc_inst.cpu_core.alu.b[14] ;
 wire \soc_inst.cpu_core.alu.b[15] ;
 wire \soc_inst.cpu_core.alu.b[16] ;
 wire \soc_inst.cpu_core.alu.b[17] ;
 wire \soc_inst.cpu_core.alu.b[18] ;
 wire \soc_inst.cpu_core.alu.b[19] ;
 wire \soc_inst.cpu_core.alu.b[1] ;
 wire \soc_inst.cpu_core.alu.b[20] ;
 wire \soc_inst.cpu_core.alu.b[21] ;
 wire \soc_inst.cpu_core.alu.b[22] ;
 wire \soc_inst.cpu_core.alu.b[23] ;
 wire \soc_inst.cpu_core.alu.b[24] ;
 wire \soc_inst.cpu_core.alu.b[25] ;
 wire \soc_inst.cpu_core.alu.b[26] ;
 wire \soc_inst.cpu_core.alu.b[27] ;
 wire \soc_inst.cpu_core.alu.b[28] ;
 wire \soc_inst.cpu_core.alu.b[29] ;
 wire \soc_inst.cpu_core.alu.b[2] ;
 wire \soc_inst.cpu_core.alu.b[30] ;
 wire \soc_inst.cpu_core.alu.b[31] ;
 wire \soc_inst.cpu_core.alu.b[3] ;
 wire \soc_inst.cpu_core.alu.b[4] ;
 wire \soc_inst.cpu_core.alu.b[5] ;
 wire \soc_inst.cpu_core.alu.b[6] ;
 wire \soc_inst.cpu_core.alu.b[7] ;
 wire \soc_inst.cpu_core.alu.b[8] ;
 wire \soc_inst.cpu_core.alu.b[9] ;
 wire \soc_inst.cpu_core.alu.op[0] ;
 wire \soc_inst.cpu_core.alu.op[1] ;
 wire \soc_inst.cpu_core.alu.op[2] ;
 wire \soc_inst.cpu_core.alu.op[3] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[0] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[10] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[11] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[1] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[2] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[3] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[4] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[5] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[6] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[7] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[8] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[9] ;
 wire \soc_inst.cpu_core.csr_file.external_interrupt ;
 wire \soc_inst.cpu_core.csr_file.mcause[0] ;
 wire \soc_inst.cpu_core.csr_file.mcause[10] ;
 wire \soc_inst.cpu_core.csr_file.mcause[11] ;
 wire \soc_inst.cpu_core.csr_file.mcause[12] ;
 wire \soc_inst.cpu_core.csr_file.mcause[13] ;
 wire \soc_inst.cpu_core.csr_file.mcause[14] ;
 wire \soc_inst.cpu_core.csr_file.mcause[15] ;
 wire \soc_inst.cpu_core.csr_file.mcause[16] ;
 wire \soc_inst.cpu_core.csr_file.mcause[17] ;
 wire \soc_inst.cpu_core.csr_file.mcause[18] ;
 wire \soc_inst.cpu_core.csr_file.mcause[19] ;
 wire \soc_inst.cpu_core.csr_file.mcause[1] ;
 wire \soc_inst.cpu_core.csr_file.mcause[20] ;
 wire \soc_inst.cpu_core.csr_file.mcause[21] ;
 wire \soc_inst.cpu_core.csr_file.mcause[22] ;
 wire \soc_inst.cpu_core.csr_file.mcause[23] ;
 wire \soc_inst.cpu_core.csr_file.mcause[24] ;
 wire \soc_inst.cpu_core.csr_file.mcause[25] ;
 wire \soc_inst.cpu_core.csr_file.mcause[26] ;
 wire \soc_inst.cpu_core.csr_file.mcause[27] ;
 wire \soc_inst.cpu_core.csr_file.mcause[28] ;
 wire \soc_inst.cpu_core.csr_file.mcause[29] ;
 wire \soc_inst.cpu_core.csr_file.mcause[2] ;
 wire \soc_inst.cpu_core.csr_file.mcause[30] ;
 wire \soc_inst.cpu_core.csr_file.mcause[31] ;
 wire \soc_inst.cpu_core.csr_file.mcause[3] ;
 wire \soc_inst.cpu_core.csr_file.mcause[4] ;
 wire \soc_inst.cpu_core.csr_file.mcause[5] ;
 wire \soc_inst.cpu_core.csr_file.mcause[6] ;
 wire \soc_inst.cpu_core.csr_file.mcause[7] ;
 wire \soc_inst.cpu_core.csr_file.mcause[8] ;
 wire \soc_inst.cpu_core.csr_file.mcause[9] ;
 wire \soc_inst.cpu_core.csr_file.mepc[0] ;
 wire \soc_inst.cpu_core.csr_file.mepc[10] ;
 wire \soc_inst.cpu_core.csr_file.mepc[11] ;
 wire \soc_inst.cpu_core.csr_file.mepc[12] ;
 wire \soc_inst.cpu_core.csr_file.mepc[13] ;
 wire \soc_inst.cpu_core.csr_file.mepc[14] ;
 wire \soc_inst.cpu_core.csr_file.mepc[15] ;
 wire \soc_inst.cpu_core.csr_file.mepc[16] ;
 wire \soc_inst.cpu_core.csr_file.mepc[17] ;
 wire \soc_inst.cpu_core.csr_file.mepc[18] ;
 wire \soc_inst.cpu_core.csr_file.mepc[19] ;
 wire \soc_inst.cpu_core.csr_file.mepc[1] ;
 wire \soc_inst.cpu_core.csr_file.mepc[20] ;
 wire \soc_inst.cpu_core.csr_file.mepc[21] ;
 wire \soc_inst.cpu_core.csr_file.mepc[22] ;
 wire \soc_inst.cpu_core.csr_file.mepc[23] ;
 wire \soc_inst.cpu_core.csr_file.mepc[2] ;
 wire \soc_inst.cpu_core.csr_file.mepc[3] ;
 wire \soc_inst.cpu_core.csr_file.mepc[4] ;
 wire \soc_inst.cpu_core.csr_file.mepc[5] ;
 wire \soc_inst.cpu_core.csr_file.mepc[6] ;
 wire \soc_inst.cpu_core.csr_file.mepc[7] ;
 wire \soc_inst.cpu_core.csr_file.mepc[8] ;
 wire \soc_inst.cpu_core.csr_file.mepc[9] ;
 wire \soc_inst.cpu_core.csr_file.mie[11] ;
 wire \soc_inst.cpu_core.csr_file.mie[7] ;
 wire \soc_inst.cpu_core.csr_file.mip_eip ;
 wire \soc_inst.cpu_core.csr_file.mip_tip ;
 wire \soc_inst.cpu_core.csr_file.mret_trigger ;
 wire \soc_inst.cpu_core.csr_file.mscratch[0] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[10] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[11] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[12] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[13] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[14] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[15] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[16] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[17] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[18] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[19] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[1] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[20] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[21] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[22] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[23] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[24] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[25] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[26] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[27] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[28] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[29] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[2] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[30] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[31] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[3] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[4] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[5] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[6] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[7] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[8] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[9] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[0] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[10] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[13] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[14] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[15] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[16] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[17] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[18] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[19] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[1] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[20] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[21] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[22] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[23] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[24] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[25] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[26] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[27] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[28] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[29] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[2] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[30] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[31] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[3] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[4] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[5] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[6] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[7] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[8] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[9] ;
 wire \soc_inst.cpu_core.csr_file.mtime[0] ;
 wire \soc_inst.cpu_core.csr_file.mtime[10] ;
 wire \soc_inst.cpu_core.csr_file.mtime[11] ;
 wire \soc_inst.cpu_core.csr_file.mtime[12] ;
 wire \soc_inst.cpu_core.csr_file.mtime[13] ;
 wire \soc_inst.cpu_core.csr_file.mtime[14] ;
 wire \soc_inst.cpu_core.csr_file.mtime[15] ;
 wire \soc_inst.cpu_core.csr_file.mtime[16] ;
 wire \soc_inst.cpu_core.csr_file.mtime[17] ;
 wire \soc_inst.cpu_core.csr_file.mtime[18] ;
 wire \soc_inst.cpu_core.csr_file.mtime[19] ;
 wire \soc_inst.cpu_core.csr_file.mtime[1] ;
 wire \soc_inst.cpu_core.csr_file.mtime[20] ;
 wire \soc_inst.cpu_core.csr_file.mtime[21] ;
 wire \soc_inst.cpu_core.csr_file.mtime[22] ;
 wire \soc_inst.cpu_core.csr_file.mtime[23] ;
 wire \soc_inst.cpu_core.csr_file.mtime[24] ;
 wire \soc_inst.cpu_core.csr_file.mtime[25] ;
 wire \soc_inst.cpu_core.csr_file.mtime[26] ;
 wire \soc_inst.cpu_core.csr_file.mtime[27] ;
 wire \soc_inst.cpu_core.csr_file.mtime[28] ;
 wire \soc_inst.cpu_core.csr_file.mtime[29] ;
 wire \soc_inst.cpu_core.csr_file.mtime[2] ;
 wire \soc_inst.cpu_core.csr_file.mtime[30] ;
 wire \soc_inst.cpu_core.csr_file.mtime[31] ;
 wire \soc_inst.cpu_core.csr_file.mtime[32] ;
 wire \soc_inst.cpu_core.csr_file.mtime[33] ;
 wire \soc_inst.cpu_core.csr_file.mtime[34] ;
 wire \soc_inst.cpu_core.csr_file.mtime[35] ;
 wire \soc_inst.cpu_core.csr_file.mtime[36] ;
 wire \soc_inst.cpu_core.csr_file.mtime[37] ;
 wire \soc_inst.cpu_core.csr_file.mtime[38] ;
 wire \soc_inst.cpu_core.csr_file.mtime[39] ;
 wire \soc_inst.cpu_core.csr_file.mtime[3] ;
 wire \soc_inst.cpu_core.csr_file.mtime[40] ;
 wire \soc_inst.cpu_core.csr_file.mtime[41] ;
 wire \soc_inst.cpu_core.csr_file.mtime[42] ;
 wire \soc_inst.cpu_core.csr_file.mtime[43] ;
 wire \soc_inst.cpu_core.csr_file.mtime[44] ;
 wire \soc_inst.cpu_core.csr_file.mtime[45] ;
 wire \soc_inst.cpu_core.csr_file.mtime[46] ;
 wire \soc_inst.cpu_core.csr_file.mtime[47] ;
 wire \soc_inst.cpu_core.csr_file.mtime[4] ;
 wire \soc_inst.cpu_core.csr_file.mtime[5] ;
 wire \soc_inst.cpu_core.csr_file.mtime[6] ;
 wire \soc_inst.cpu_core.csr_file.mtime[7] ;
 wire \soc_inst.cpu_core.csr_file.mtime[8] ;
 wire \soc_inst.cpu_core.csr_file.mtime[9] ;
 wire \soc_inst.cpu_core.csr_file.mtval[0] ;
 wire \soc_inst.cpu_core.csr_file.mtval[10] ;
 wire \soc_inst.cpu_core.csr_file.mtval[11] ;
 wire \soc_inst.cpu_core.csr_file.mtval[12] ;
 wire \soc_inst.cpu_core.csr_file.mtval[13] ;
 wire \soc_inst.cpu_core.csr_file.mtval[14] ;
 wire \soc_inst.cpu_core.csr_file.mtval[15] ;
 wire \soc_inst.cpu_core.csr_file.mtval[16] ;
 wire \soc_inst.cpu_core.csr_file.mtval[17] ;
 wire \soc_inst.cpu_core.csr_file.mtval[18] ;
 wire \soc_inst.cpu_core.csr_file.mtval[19] ;
 wire \soc_inst.cpu_core.csr_file.mtval[1] ;
 wire \soc_inst.cpu_core.csr_file.mtval[20] ;
 wire \soc_inst.cpu_core.csr_file.mtval[21] ;
 wire \soc_inst.cpu_core.csr_file.mtval[22] ;
 wire \soc_inst.cpu_core.csr_file.mtval[23] ;
 wire \soc_inst.cpu_core.csr_file.mtval[24] ;
 wire \soc_inst.cpu_core.csr_file.mtval[25] ;
 wire \soc_inst.cpu_core.csr_file.mtval[26] ;
 wire \soc_inst.cpu_core.csr_file.mtval[27] ;
 wire \soc_inst.cpu_core.csr_file.mtval[28] ;
 wire \soc_inst.cpu_core.csr_file.mtval[29] ;
 wire \soc_inst.cpu_core.csr_file.mtval[2] ;
 wire \soc_inst.cpu_core.csr_file.mtval[30] ;
 wire \soc_inst.cpu_core.csr_file.mtval[31] ;
 wire \soc_inst.cpu_core.csr_file.mtval[3] ;
 wire \soc_inst.cpu_core.csr_file.mtval[4] ;
 wire \soc_inst.cpu_core.csr_file.mtval[5] ;
 wire \soc_inst.cpu_core.csr_file.mtval[6] ;
 wire \soc_inst.cpu_core.csr_file.mtval[7] ;
 wire \soc_inst.cpu_core.csr_file.mtval[8] ;
 wire \soc_inst.cpu_core.csr_file.mtval[9] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[0] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[10] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[11] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[12] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[13] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[14] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[15] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[16] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[17] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[18] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[19] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[1] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[20] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[21] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[22] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[23] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[2] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[3] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[4] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[5] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[6] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[7] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[8] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[9] ;
 wire \soc_inst.cpu_core.csr_file.timer_interrupt ;
 wire \soc_inst.cpu_core.error_flag_reg ;
 wire \soc_inst.cpu_core.ex_alu_result[0] ;
 wire \soc_inst.cpu_core.ex_alu_result[10] ;
 wire \soc_inst.cpu_core.ex_alu_result[11] ;
 wire \soc_inst.cpu_core.ex_alu_result[12] ;
 wire \soc_inst.cpu_core.ex_alu_result[13] ;
 wire \soc_inst.cpu_core.ex_alu_result[14] ;
 wire \soc_inst.cpu_core.ex_alu_result[15] ;
 wire \soc_inst.cpu_core.ex_alu_result[16] ;
 wire \soc_inst.cpu_core.ex_alu_result[17] ;
 wire \soc_inst.cpu_core.ex_alu_result[18] ;
 wire \soc_inst.cpu_core.ex_alu_result[19] ;
 wire \soc_inst.cpu_core.ex_alu_result[1] ;
 wire \soc_inst.cpu_core.ex_alu_result[20] ;
 wire \soc_inst.cpu_core.ex_alu_result[21] ;
 wire \soc_inst.cpu_core.ex_alu_result[22] ;
 wire \soc_inst.cpu_core.ex_alu_result[23] ;
 wire \soc_inst.cpu_core.ex_alu_result[24] ;
 wire \soc_inst.cpu_core.ex_alu_result[25] ;
 wire \soc_inst.cpu_core.ex_alu_result[26] ;
 wire \soc_inst.cpu_core.ex_alu_result[27] ;
 wire \soc_inst.cpu_core.ex_alu_result[28] ;
 wire \soc_inst.cpu_core.ex_alu_result[29] ;
 wire \soc_inst.cpu_core.ex_alu_result[2] ;
 wire \soc_inst.cpu_core.ex_alu_result[30] ;
 wire \soc_inst.cpu_core.ex_alu_result[31] ;
 wire \soc_inst.cpu_core.ex_alu_result[3] ;
 wire \soc_inst.cpu_core.ex_alu_result[4] ;
 wire \soc_inst.cpu_core.ex_alu_result[5] ;
 wire \soc_inst.cpu_core.ex_alu_result[6] ;
 wire \soc_inst.cpu_core.ex_alu_result[7] ;
 wire \soc_inst.cpu_core.ex_alu_result[8] ;
 wire \soc_inst.cpu_core.ex_alu_result[9] ;
 wire \soc_inst.cpu_core.ex_branch_target[0] ;
 wire \soc_inst.cpu_core.ex_branch_target[10] ;
 wire \soc_inst.cpu_core.ex_branch_target[11] ;
 wire \soc_inst.cpu_core.ex_branch_target[12] ;
 wire \soc_inst.cpu_core.ex_branch_target[13] ;
 wire \soc_inst.cpu_core.ex_branch_target[14] ;
 wire \soc_inst.cpu_core.ex_branch_target[15] ;
 wire \soc_inst.cpu_core.ex_branch_target[16] ;
 wire \soc_inst.cpu_core.ex_branch_target[17] ;
 wire \soc_inst.cpu_core.ex_branch_target[18] ;
 wire \soc_inst.cpu_core.ex_branch_target[19] ;
 wire \soc_inst.cpu_core.ex_branch_target[1] ;
 wire \soc_inst.cpu_core.ex_branch_target[20] ;
 wire \soc_inst.cpu_core.ex_branch_target[21] ;
 wire \soc_inst.cpu_core.ex_branch_target[22] ;
 wire \soc_inst.cpu_core.ex_branch_target[23] ;
 wire \soc_inst.cpu_core.ex_branch_target[24] ;
 wire \soc_inst.cpu_core.ex_branch_target[25] ;
 wire \soc_inst.cpu_core.ex_branch_target[26] ;
 wire \soc_inst.cpu_core.ex_branch_target[27] ;
 wire \soc_inst.cpu_core.ex_branch_target[28] ;
 wire \soc_inst.cpu_core.ex_branch_target[29] ;
 wire \soc_inst.cpu_core.ex_branch_target[2] ;
 wire \soc_inst.cpu_core.ex_branch_target[30] ;
 wire \soc_inst.cpu_core.ex_branch_target[31] ;
 wire \soc_inst.cpu_core.ex_branch_target[3] ;
 wire \soc_inst.cpu_core.ex_branch_target[4] ;
 wire \soc_inst.cpu_core.ex_branch_target[5] ;
 wire \soc_inst.cpu_core.ex_branch_target[6] ;
 wire \soc_inst.cpu_core.ex_branch_target[7] ;
 wire \soc_inst.cpu_core.ex_branch_target[8] ;
 wire \soc_inst.cpu_core.ex_branch_target[9] ;
 wire \soc_inst.cpu_core.ex_exception_pc[0] ;
 wire \soc_inst.cpu_core.ex_exception_pc[10] ;
 wire \soc_inst.cpu_core.ex_exception_pc[11] ;
 wire \soc_inst.cpu_core.ex_exception_pc[12] ;
 wire \soc_inst.cpu_core.ex_exception_pc[13] ;
 wire \soc_inst.cpu_core.ex_exception_pc[14] ;
 wire \soc_inst.cpu_core.ex_exception_pc[15] ;
 wire \soc_inst.cpu_core.ex_exception_pc[16] ;
 wire \soc_inst.cpu_core.ex_exception_pc[17] ;
 wire \soc_inst.cpu_core.ex_exception_pc[18] ;
 wire \soc_inst.cpu_core.ex_exception_pc[19] ;
 wire \soc_inst.cpu_core.ex_exception_pc[1] ;
 wire \soc_inst.cpu_core.ex_exception_pc[20] ;
 wire \soc_inst.cpu_core.ex_exception_pc[21] ;
 wire \soc_inst.cpu_core.ex_exception_pc[22] ;
 wire \soc_inst.cpu_core.ex_exception_pc[23] ;
 wire \soc_inst.cpu_core.ex_exception_pc[2] ;
 wire \soc_inst.cpu_core.ex_exception_pc[3] ;
 wire \soc_inst.cpu_core.ex_exception_pc[4] ;
 wire \soc_inst.cpu_core.ex_exception_pc[5] ;
 wire \soc_inst.cpu_core.ex_exception_pc[6] ;
 wire \soc_inst.cpu_core.ex_exception_pc[7] ;
 wire \soc_inst.cpu_core.ex_exception_pc[8] ;
 wire \soc_inst.cpu_core.ex_exception_pc[9] ;
 wire \soc_inst.cpu_core.ex_funct3[0] ;
 wire \soc_inst.cpu_core.ex_funct3[1] ;
 wire \soc_inst.cpu_core.ex_funct3[2] ;
 wire \soc_inst.cpu_core.ex_funct7[0] ;
 wire \soc_inst.cpu_core.ex_funct7[1] ;
 wire \soc_inst.cpu_core.ex_funct7[2] ;
 wire \soc_inst.cpu_core.ex_funct7[3] ;
 wire \soc_inst.cpu_core.ex_funct7[4] ;
 wire \soc_inst.cpu_core.ex_funct7[5] ;
 wire \soc_inst.cpu_core.ex_funct7[6] ;
 wire \soc_inst.cpu_core.ex_instr[10] ;
 wire \soc_inst.cpu_core.ex_instr[11] ;
 wire \soc_inst.cpu_core.ex_instr[15] ;
 wire \soc_inst.cpu_core.ex_instr[16] ;
 wire \soc_inst.cpu_core.ex_instr[17] ;
 wire \soc_inst.cpu_core.ex_instr[18] ;
 wire \soc_inst.cpu_core.ex_instr[19] ;
 wire \soc_inst.cpu_core.ex_instr[20] ;
 wire \soc_inst.cpu_core.ex_instr[21] ;
 wire \soc_inst.cpu_core.ex_instr[22] ;
 wire \soc_inst.cpu_core.ex_instr[23] ;
 wire \soc_inst.cpu_core.ex_instr[24] ;
 wire \soc_inst.cpu_core.ex_instr[2] ;
 wire \soc_inst.cpu_core.ex_instr[3] ;
 wire \soc_inst.cpu_core.ex_instr[5] ;
 wire \soc_inst.cpu_core.ex_instr[6] ;
 wire \soc_inst.cpu_core.ex_instr[7] ;
 wire \soc_inst.cpu_core.ex_instr[8] ;
 wire \soc_inst.cpu_core.ex_instr[9] ;
 wire \soc_inst.cpu_core.ex_is_ebreak ;
 wire \soc_inst.cpu_core.ex_is_ecall ;
 wire \soc_inst.cpu_core.ex_mem_re ;
 wire \soc_inst.cpu_core.ex_mem_we ;
 wire \soc_inst.cpu_core.ex_reg_we ;
 wire \soc_inst.cpu_core.ex_rs1_data[0] ;
 wire \soc_inst.cpu_core.ex_rs1_data[10] ;
 wire \soc_inst.cpu_core.ex_rs1_data[11] ;
 wire \soc_inst.cpu_core.ex_rs1_data[12] ;
 wire \soc_inst.cpu_core.ex_rs1_data[13] ;
 wire \soc_inst.cpu_core.ex_rs1_data[14] ;
 wire \soc_inst.cpu_core.ex_rs1_data[15] ;
 wire \soc_inst.cpu_core.ex_rs1_data[16] ;
 wire \soc_inst.cpu_core.ex_rs1_data[17] ;
 wire \soc_inst.cpu_core.ex_rs1_data[18] ;
 wire \soc_inst.cpu_core.ex_rs1_data[19] ;
 wire \soc_inst.cpu_core.ex_rs1_data[1] ;
 wire \soc_inst.cpu_core.ex_rs1_data[20] ;
 wire \soc_inst.cpu_core.ex_rs1_data[21] ;
 wire \soc_inst.cpu_core.ex_rs1_data[22] ;
 wire \soc_inst.cpu_core.ex_rs1_data[23] ;
 wire \soc_inst.cpu_core.ex_rs1_data[24] ;
 wire \soc_inst.cpu_core.ex_rs1_data[25] ;
 wire \soc_inst.cpu_core.ex_rs1_data[26] ;
 wire \soc_inst.cpu_core.ex_rs1_data[27] ;
 wire \soc_inst.cpu_core.ex_rs1_data[28] ;
 wire \soc_inst.cpu_core.ex_rs1_data[29] ;
 wire \soc_inst.cpu_core.ex_rs1_data[2] ;
 wire \soc_inst.cpu_core.ex_rs1_data[30] ;
 wire \soc_inst.cpu_core.ex_rs1_data[31] ;
 wire \soc_inst.cpu_core.ex_rs1_data[3] ;
 wire \soc_inst.cpu_core.ex_rs1_data[4] ;
 wire \soc_inst.cpu_core.ex_rs1_data[5] ;
 wire \soc_inst.cpu_core.ex_rs1_data[6] ;
 wire \soc_inst.cpu_core.ex_rs1_data[7] ;
 wire \soc_inst.cpu_core.ex_rs1_data[8] ;
 wire \soc_inst.cpu_core.ex_rs1_data[9] ;
 wire \soc_inst.cpu_core.ex_rs2_data[0] ;
 wire \soc_inst.cpu_core.ex_rs2_data[10] ;
 wire \soc_inst.cpu_core.ex_rs2_data[11] ;
 wire \soc_inst.cpu_core.ex_rs2_data[12] ;
 wire \soc_inst.cpu_core.ex_rs2_data[13] ;
 wire \soc_inst.cpu_core.ex_rs2_data[14] ;
 wire \soc_inst.cpu_core.ex_rs2_data[15] ;
 wire \soc_inst.cpu_core.ex_rs2_data[16] ;
 wire \soc_inst.cpu_core.ex_rs2_data[17] ;
 wire \soc_inst.cpu_core.ex_rs2_data[18] ;
 wire \soc_inst.cpu_core.ex_rs2_data[19] ;
 wire \soc_inst.cpu_core.ex_rs2_data[1] ;
 wire \soc_inst.cpu_core.ex_rs2_data[20] ;
 wire \soc_inst.cpu_core.ex_rs2_data[21] ;
 wire \soc_inst.cpu_core.ex_rs2_data[22] ;
 wire \soc_inst.cpu_core.ex_rs2_data[23] ;
 wire \soc_inst.cpu_core.ex_rs2_data[24] ;
 wire \soc_inst.cpu_core.ex_rs2_data[25] ;
 wire \soc_inst.cpu_core.ex_rs2_data[26] ;
 wire \soc_inst.cpu_core.ex_rs2_data[27] ;
 wire \soc_inst.cpu_core.ex_rs2_data[28] ;
 wire \soc_inst.cpu_core.ex_rs2_data[29] ;
 wire \soc_inst.cpu_core.ex_rs2_data[2] ;
 wire \soc_inst.cpu_core.ex_rs2_data[30] ;
 wire \soc_inst.cpu_core.ex_rs2_data[31] ;
 wire \soc_inst.cpu_core.ex_rs2_data[3] ;
 wire \soc_inst.cpu_core.ex_rs2_data[4] ;
 wire \soc_inst.cpu_core.ex_rs2_data[5] ;
 wire \soc_inst.cpu_core.ex_rs2_data[6] ;
 wire \soc_inst.cpu_core.ex_rs2_data[7] ;
 wire \soc_inst.cpu_core.ex_rs2_data[8] ;
 wire \soc_inst.cpu_core.ex_rs2_data[9] ;
 wire \soc_inst.cpu_core.i_mem_ready ;
 wire \soc_inst.cpu_core.id_funct3[0] ;
 wire \soc_inst.cpu_core.id_funct3[1] ;
 wire \soc_inst.cpu_core.id_funct3[2] ;
 wire \soc_inst.cpu_core.id_imm12[0] ;
 wire \soc_inst.cpu_core.id_imm12[10] ;
 wire \soc_inst.cpu_core.id_imm12[11] ;
 wire \soc_inst.cpu_core.id_imm12[1] ;
 wire \soc_inst.cpu_core.id_imm12[2] ;
 wire \soc_inst.cpu_core.id_imm12[3] ;
 wire \soc_inst.cpu_core.id_imm12[4] ;
 wire \soc_inst.cpu_core.id_imm12[5] ;
 wire \soc_inst.cpu_core.id_imm12[6] ;
 wire \soc_inst.cpu_core.id_imm12[7] ;
 wire \soc_inst.cpu_core.id_imm12[8] ;
 wire \soc_inst.cpu_core.id_imm12[9] ;
 wire \soc_inst.cpu_core.id_imm[0] ;
 wire \soc_inst.cpu_core.id_imm[10] ;
 wire \soc_inst.cpu_core.id_imm[11] ;
 wire \soc_inst.cpu_core.id_imm[12] ;
 wire \soc_inst.cpu_core.id_imm[13] ;
 wire \soc_inst.cpu_core.id_imm[14] ;
 wire \soc_inst.cpu_core.id_imm[15] ;
 wire \soc_inst.cpu_core.id_imm[16] ;
 wire \soc_inst.cpu_core.id_imm[17] ;
 wire \soc_inst.cpu_core.id_imm[18] ;
 wire \soc_inst.cpu_core.id_imm[19] ;
 wire \soc_inst.cpu_core.id_imm[1] ;
 wire \soc_inst.cpu_core.id_imm[20] ;
 wire \soc_inst.cpu_core.id_imm[21] ;
 wire \soc_inst.cpu_core.id_imm[22] ;
 wire \soc_inst.cpu_core.id_imm[23] ;
 wire \soc_inst.cpu_core.id_imm[24] ;
 wire \soc_inst.cpu_core.id_imm[25] ;
 wire \soc_inst.cpu_core.id_imm[26] ;
 wire \soc_inst.cpu_core.id_imm[27] ;
 wire \soc_inst.cpu_core.id_imm[28] ;
 wire \soc_inst.cpu_core.id_imm[29] ;
 wire \soc_inst.cpu_core.id_imm[2] ;
 wire \soc_inst.cpu_core.id_imm[30] ;
 wire \soc_inst.cpu_core.id_imm[31] ;
 wire \soc_inst.cpu_core.id_imm[3] ;
 wire \soc_inst.cpu_core.id_imm[4] ;
 wire \soc_inst.cpu_core.id_imm[5] ;
 wire \soc_inst.cpu_core.id_imm[6] ;
 wire \soc_inst.cpu_core.id_imm[7] ;
 wire \soc_inst.cpu_core.id_imm[8] ;
 wire \soc_inst.cpu_core.id_imm[9] ;
 wire \soc_inst.cpu_core.id_instr[10] ;
 wire \soc_inst.cpu_core.id_instr[11] ;
 wire \soc_inst.cpu_core.id_instr[15] ;
 wire \soc_inst.cpu_core.id_instr[16] ;
 wire \soc_inst.cpu_core.id_instr[17] ;
 wire \soc_inst.cpu_core.id_instr[18] ;
 wire \soc_inst.cpu_core.id_instr[19] ;
 wire \soc_inst.cpu_core.id_instr[2] ;
 wire \soc_inst.cpu_core.id_instr[3] ;
 wire \soc_inst.cpu_core.id_instr[5] ;
 wire \soc_inst.cpu_core.id_instr[6] ;
 wire \soc_inst.cpu_core.id_instr[7] ;
 wire \soc_inst.cpu_core.id_instr[8] ;
 wire \soc_inst.cpu_core.id_instr[9] ;
 wire \soc_inst.cpu_core.id_int_is_interrupt ;
 wire \soc_inst.cpu_core.id_is_compressed ;
 wire \soc_inst.cpu_core.id_pc[0] ;
 wire \soc_inst.cpu_core.id_pc[10] ;
 wire \soc_inst.cpu_core.id_pc[11] ;
 wire \soc_inst.cpu_core.id_pc[12] ;
 wire \soc_inst.cpu_core.id_pc[13] ;
 wire \soc_inst.cpu_core.id_pc[14] ;
 wire \soc_inst.cpu_core.id_pc[15] ;
 wire \soc_inst.cpu_core.id_pc[16] ;
 wire \soc_inst.cpu_core.id_pc[17] ;
 wire \soc_inst.cpu_core.id_pc[18] ;
 wire \soc_inst.cpu_core.id_pc[19] ;
 wire \soc_inst.cpu_core.id_pc[1] ;
 wire \soc_inst.cpu_core.id_pc[20] ;
 wire \soc_inst.cpu_core.id_pc[21] ;
 wire \soc_inst.cpu_core.id_pc[22] ;
 wire \soc_inst.cpu_core.id_pc[23] ;
 wire \soc_inst.cpu_core.id_pc[2] ;
 wire \soc_inst.cpu_core.id_pc[3] ;
 wire \soc_inst.cpu_core.id_pc[4] ;
 wire \soc_inst.cpu_core.id_pc[5] ;
 wire \soc_inst.cpu_core.id_pc[6] ;
 wire \soc_inst.cpu_core.id_pc[7] ;
 wire \soc_inst.cpu_core.id_pc[8] ;
 wire \soc_inst.cpu_core.id_pc[9] ;
 wire \soc_inst.cpu_core.id_rs1_data[0] ;
 wire \soc_inst.cpu_core.id_rs1_data[10] ;
 wire \soc_inst.cpu_core.id_rs1_data[11] ;
 wire \soc_inst.cpu_core.id_rs1_data[12] ;
 wire \soc_inst.cpu_core.id_rs1_data[13] ;
 wire \soc_inst.cpu_core.id_rs1_data[14] ;
 wire \soc_inst.cpu_core.id_rs1_data[15] ;
 wire \soc_inst.cpu_core.id_rs1_data[16] ;
 wire \soc_inst.cpu_core.id_rs1_data[17] ;
 wire \soc_inst.cpu_core.id_rs1_data[18] ;
 wire \soc_inst.cpu_core.id_rs1_data[19] ;
 wire \soc_inst.cpu_core.id_rs1_data[1] ;
 wire \soc_inst.cpu_core.id_rs1_data[20] ;
 wire \soc_inst.cpu_core.id_rs1_data[21] ;
 wire \soc_inst.cpu_core.id_rs1_data[22] ;
 wire \soc_inst.cpu_core.id_rs1_data[23] ;
 wire \soc_inst.cpu_core.id_rs1_data[24] ;
 wire \soc_inst.cpu_core.id_rs1_data[25] ;
 wire \soc_inst.cpu_core.id_rs1_data[26] ;
 wire \soc_inst.cpu_core.id_rs1_data[27] ;
 wire \soc_inst.cpu_core.id_rs1_data[28] ;
 wire \soc_inst.cpu_core.id_rs1_data[29] ;
 wire \soc_inst.cpu_core.id_rs1_data[2] ;
 wire \soc_inst.cpu_core.id_rs1_data[30] ;
 wire \soc_inst.cpu_core.id_rs1_data[31] ;
 wire \soc_inst.cpu_core.id_rs1_data[3] ;
 wire \soc_inst.cpu_core.id_rs1_data[4] ;
 wire \soc_inst.cpu_core.id_rs1_data[5] ;
 wire \soc_inst.cpu_core.id_rs1_data[6] ;
 wire \soc_inst.cpu_core.id_rs1_data[7] ;
 wire \soc_inst.cpu_core.id_rs1_data[8] ;
 wire \soc_inst.cpu_core.id_rs1_data[9] ;
 wire \soc_inst.cpu_core.id_rs2_data[0] ;
 wire \soc_inst.cpu_core.id_rs2_data[10] ;
 wire \soc_inst.cpu_core.id_rs2_data[11] ;
 wire \soc_inst.cpu_core.id_rs2_data[12] ;
 wire \soc_inst.cpu_core.id_rs2_data[13] ;
 wire \soc_inst.cpu_core.id_rs2_data[14] ;
 wire \soc_inst.cpu_core.id_rs2_data[15] ;
 wire \soc_inst.cpu_core.id_rs2_data[16] ;
 wire \soc_inst.cpu_core.id_rs2_data[17] ;
 wire \soc_inst.cpu_core.id_rs2_data[18] ;
 wire \soc_inst.cpu_core.id_rs2_data[19] ;
 wire \soc_inst.cpu_core.id_rs2_data[1] ;
 wire \soc_inst.cpu_core.id_rs2_data[20] ;
 wire \soc_inst.cpu_core.id_rs2_data[21] ;
 wire \soc_inst.cpu_core.id_rs2_data[22] ;
 wire \soc_inst.cpu_core.id_rs2_data[23] ;
 wire \soc_inst.cpu_core.id_rs2_data[24] ;
 wire \soc_inst.cpu_core.id_rs2_data[25] ;
 wire \soc_inst.cpu_core.id_rs2_data[26] ;
 wire \soc_inst.cpu_core.id_rs2_data[27] ;
 wire \soc_inst.cpu_core.id_rs2_data[28] ;
 wire \soc_inst.cpu_core.id_rs2_data[29] ;
 wire \soc_inst.cpu_core.id_rs2_data[2] ;
 wire \soc_inst.cpu_core.id_rs2_data[30] ;
 wire \soc_inst.cpu_core.id_rs2_data[31] ;
 wire \soc_inst.cpu_core.id_rs2_data[3] ;
 wire \soc_inst.cpu_core.id_rs2_data[4] ;
 wire \soc_inst.cpu_core.id_rs2_data[5] ;
 wire \soc_inst.cpu_core.id_rs2_data[6] ;
 wire \soc_inst.cpu_core.id_rs2_data[7] ;
 wire \soc_inst.cpu_core.id_rs2_data[8] ;
 wire \soc_inst.cpu_core.id_rs2_data[9] ;
 wire \soc_inst.cpu_core.if_funct3[0] ;
 wire \soc_inst.cpu_core.if_funct3[1] ;
 wire \soc_inst.cpu_core.if_funct3[2] ;
 wire \soc_inst.cpu_core.if_funct7[0] ;
 wire \soc_inst.cpu_core.if_funct7[1] ;
 wire \soc_inst.cpu_core.if_funct7[2] ;
 wire \soc_inst.cpu_core.if_funct7[3] ;
 wire \soc_inst.cpu_core.if_funct7[4] ;
 wire \soc_inst.cpu_core.if_funct7[5] ;
 wire \soc_inst.cpu_core.if_funct7[6] ;
 wire \soc_inst.cpu_core.if_imm12[0] ;
 wire \soc_inst.cpu_core.if_imm12[1] ;
 wire \soc_inst.cpu_core.if_imm12[2] ;
 wire \soc_inst.cpu_core.if_imm12[3] ;
 wire \soc_inst.cpu_core.if_imm12[4] ;
 wire \soc_inst.cpu_core.if_instr[10] ;
 wire \soc_inst.cpu_core.if_instr[11] ;
 wire \soc_inst.cpu_core.if_instr[15] ;
 wire \soc_inst.cpu_core.if_instr[16] ;
 wire \soc_inst.cpu_core.if_instr[17] ;
 wire \soc_inst.cpu_core.if_instr[18] ;
 wire \soc_inst.cpu_core.if_instr[19] ;
 wire \soc_inst.cpu_core.if_instr[2] ;
 wire \soc_inst.cpu_core.if_instr[3] ;
 wire \soc_inst.cpu_core.if_instr[5] ;
 wire \soc_inst.cpu_core.if_instr[6] ;
 wire \soc_inst.cpu_core.if_instr[7] ;
 wire \soc_inst.cpu_core.if_instr[8] ;
 wire \soc_inst.cpu_core.if_instr[9] ;
 wire \soc_inst.cpu_core.if_is_compressed ;
 wire \soc_inst.cpu_core.if_pc[0] ;
 wire \soc_inst.cpu_core.if_pc[10] ;
 wire \soc_inst.cpu_core.if_pc[11] ;
 wire \soc_inst.cpu_core.if_pc[12] ;
 wire \soc_inst.cpu_core.if_pc[13] ;
 wire \soc_inst.cpu_core.if_pc[14] ;
 wire \soc_inst.cpu_core.if_pc[15] ;
 wire \soc_inst.cpu_core.if_pc[16] ;
 wire \soc_inst.cpu_core.if_pc[17] ;
 wire \soc_inst.cpu_core.if_pc[18] ;
 wire \soc_inst.cpu_core.if_pc[19] ;
 wire \soc_inst.cpu_core.if_pc[1] ;
 wire \soc_inst.cpu_core.if_pc[20] ;
 wire \soc_inst.cpu_core.if_pc[21] ;
 wire \soc_inst.cpu_core.if_pc[22] ;
 wire \soc_inst.cpu_core.if_pc[23] ;
 wire \soc_inst.cpu_core.if_pc[2] ;
 wire \soc_inst.cpu_core.if_pc[3] ;
 wire \soc_inst.cpu_core.if_pc[4] ;
 wire \soc_inst.cpu_core.if_pc[5] ;
 wire \soc_inst.cpu_core.if_pc[6] ;
 wire \soc_inst.cpu_core.if_pc[7] ;
 wire \soc_inst.cpu_core.if_pc[8] ;
 wire \soc_inst.cpu_core.if_pc[9] ;
 wire \soc_inst.cpu_core.mem_instr[15] ;
 wire \soc_inst.cpu_core.mem_instr[16] ;
 wire \soc_inst.cpu_core.mem_instr[17] ;
 wire \soc_inst.cpu_core.mem_instr[18] ;
 wire \soc_inst.cpu_core.mem_instr[19] ;
 wire \soc_inst.cpu_core.mem_instr[2] ;
 wire \soc_inst.cpu_core.mem_instr[3] ;
 wire \soc_inst.cpu_core.mem_instr[5] ;
 wire \soc_inst.cpu_core.mem_instr[6] ;
 wire \soc_inst.cpu_core.mem_reg_we ;
 wire \soc_inst.cpu_core.mem_rs1_data[0] ;
 wire \soc_inst.cpu_core.mem_rs1_data[10] ;
 wire \soc_inst.cpu_core.mem_rs1_data[11] ;
 wire \soc_inst.cpu_core.mem_rs1_data[12] ;
 wire \soc_inst.cpu_core.mem_rs1_data[13] ;
 wire \soc_inst.cpu_core.mem_rs1_data[14] ;
 wire \soc_inst.cpu_core.mem_rs1_data[15] ;
 wire \soc_inst.cpu_core.mem_rs1_data[16] ;
 wire \soc_inst.cpu_core.mem_rs1_data[17] ;
 wire \soc_inst.cpu_core.mem_rs1_data[18] ;
 wire \soc_inst.cpu_core.mem_rs1_data[19] ;
 wire \soc_inst.cpu_core.mem_rs1_data[1] ;
 wire \soc_inst.cpu_core.mem_rs1_data[20] ;
 wire \soc_inst.cpu_core.mem_rs1_data[21] ;
 wire \soc_inst.cpu_core.mem_rs1_data[22] ;
 wire \soc_inst.cpu_core.mem_rs1_data[23] ;
 wire \soc_inst.cpu_core.mem_rs1_data[24] ;
 wire \soc_inst.cpu_core.mem_rs1_data[25] ;
 wire \soc_inst.cpu_core.mem_rs1_data[26] ;
 wire \soc_inst.cpu_core.mem_rs1_data[27] ;
 wire \soc_inst.cpu_core.mem_rs1_data[28] ;
 wire \soc_inst.cpu_core.mem_rs1_data[29] ;
 wire \soc_inst.cpu_core.mem_rs1_data[2] ;
 wire \soc_inst.cpu_core.mem_rs1_data[30] ;
 wire \soc_inst.cpu_core.mem_rs1_data[31] ;
 wire \soc_inst.cpu_core.mem_rs1_data[3] ;
 wire \soc_inst.cpu_core.mem_rs1_data[4] ;
 wire \soc_inst.cpu_core.mem_rs1_data[5] ;
 wire \soc_inst.cpu_core.mem_rs1_data[6] ;
 wire \soc_inst.cpu_core.mem_rs1_data[7] ;
 wire \soc_inst.cpu_core.mem_rs1_data[8] ;
 wire \soc_inst.cpu_core.mem_rs1_data[9] ;
 wire \soc_inst.cpu_core.mem_stall ;
 wire \soc_inst.cpu_core.register_file.registers[10][0] ;
 wire \soc_inst.cpu_core.register_file.registers[10][10] ;
 wire \soc_inst.cpu_core.register_file.registers[10][11] ;
 wire \soc_inst.cpu_core.register_file.registers[10][12] ;
 wire \soc_inst.cpu_core.register_file.registers[10][13] ;
 wire \soc_inst.cpu_core.register_file.registers[10][14] ;
 wire \soc_inst.cpu_core.register_file.registers[10][15] ;
 wire \soc_inst.cpu_core.register_file.registers[10][16] ;
 wire \soc_inst.cpu_core.register_file.registers[10][17] ;
 wire \soc_inst.cpu_core.register_file.registers[10][18] ;
 wire \soc_inst.cpu_core.register_file.registers[10][19] ;
 wire \soc_inst.cpu_core.register_file.registers[10][1] ;
 wire \soc_inst.cpu_core.register_file.registers[10][20] ;
 wire \soc_inst.cpu_core.register_file.registers[10][21] ;
 wire \soc_inst.cpu_core.register_file.registers[10][22] ;
 wire \soc_inst.cpu_core.register_file.registers[10][23] ;
 wire \soc_inst.cpu_core.register_file.registers[10][24] ;
 wire \soc_inst.cpu_core.register_file.registers[10][25] ;
 wire \soc_inst.cpu_core.register_file.registers[10][26] ;
 wire \soc_inst.cpu_core.register_file.registers[10][27] ;
 wire \soc_inst.cpu_core.register_file.registers[10][28] ;
 wire \soc_inst.cpu_core.register_file.registers[10][29] ;
 wire \soc_inst.cpu_core.register_file.registers[10][2] ;
 wire \soc_inst.cpu_core.register_file.registers[10][30] ;
 wire \soc_inst.cpu_core.register_file.registers[10][31] ;
 wire \soc_inst.cpu_core.register_file.registers[10][3] ;
 wire \soc_inst.cpu_core.register_file.registers[10][4] ;
 wire \soc_inst.cpu_core.register_file.registers[10][5] ;
 wire \soc_inst.cpu_core.register_file.registers[10][6] ;
 wire \soc_inst.cpu_core.register_file.registers[10][7] ;
 wire \soc_inst.cpu_core.register_file.registers[10][8] ;
 wire \soc_inst.cpu_core.register_file.registers[10][9] ;
 wire \soc_inst.cpu_core.register_file.registers[11][0] ;
 wire \soc_inst.cpu_core.register_file.registers[11][10] ;
 wire \soc_inst.cpu_core.register_file.registers[11][11] ;
 wire \soc_inst.cpu_core.register_file.registers[11][12] ;
 wire \soc_inst.cpu_core.register_file.registers[11][13] ;
 wire \soc_inst.cpu_core.register_file.registers[11][14] ;
 wire \soc_inst.cpu_core.register_file.registers[11][15] ;
 wire \soc_inst.cpu_core.register_file.registers[11][16] ;
 wire \soc_inst.cpu_core.register_file.registers[11][17] ;
 wire \soc_inst.cpu_core.register_file.registers[11][18] ;
 wire \soc_inst.cpu_core.register_file.registers[11][19] ;
 wire \soc_inst.cpu_core.register_file.registers[11][1] ;
 wire \soc_inst.cpu_core.register_file.registers[11][20] ;
 wire \soc_inst.cpu_core.register_file.registers[11][21] ;
 wire \soc_inst.cpu_core.register_file.registers[11][22] ;
 wire \soc_inst.cpu_core.register_file.registers[11][23] ;
 wire \soc_inst.cpu_core.register_file.registers[11][24] ;
 wire \soc_inst.cpu_core.register_file.registers[11][25] ;
 wire \soc_inst.cpu_core.register_file.registers[11][26] ;
 wire \soc_inst.cpu_core.register_file.registers[11][27] ;
 wire \soc_inst.cpu_core.register_file.registers[11][28] ;
 wire \soc_inst.cpu_core.register_file.registers[11][29] ;
 wire \soc_inst.cpu_core.register_file.registers[11][2] ;
 wire \soc_inst.cpu_core.register_file.registers[11][30] ;
 wire \soc_inst.cpu_core.register_file.registers[11][31] ;
 wire \soc_inst.cpu_core.register_file.registers[11][3] ;
 wire \soc_inst.cpu_core.register_file.registers[11][4] ;
 wire \soc_inst.cpu_core.register_file.registers[11][5] ;
 wire \soc_inst.cpu_core.register_file.registers[11][6] ;
 wire \soc_inst.cpu_core.register_file.registers[11][7] ;
 wire \soc_inst.cpu_core.register_file.registers[11][8] ;
 wire \soc_inst.cpu_core.register_file.registers[11][9] ;
 wire \soc_inst.cpu_core.register_file.registers[12][0] ;
 wire \soc_inst.cpu_core.register_file.registers[12][10] ;
 wire \soc_inst.cpu_core.register_file.registers[12][11] ;
 wire \soc_inst.cpu_core.register_file.registers[12][12] ;
 wire \soc_inst.cpu_core.register_file.registers[12][13] ;
 wire \soc_inst.cpu_core.register_file.registers[12][14] ;
 wire \soc_inst.cpu_core.register_file.registers[12][15] ;
 wire \soc_inst.cpu_core.register_file.registers[12][16] ;
 wire \soc_inst.cpu_core.register_file.registers[12][17] ;
 wire \soc_inst.cpu_core.register_file.registers[12][18] ;
 wire \soc_inst.cpu_core.register_file.registers[12][19] ;
 wire \soc_inst.cpu_core.register_file.registers[12][1] ;
 wire \soc_inst.cpu_core.register_file.registers[12][20] ;
 wire \soc_inst.cpu_core.register_file.registers[12][21] ;
 wire \soc_inst.cpu_core.register_file.registers[12][22] ;
 wire \soc_inst.cpu_core.register_file.registers[12][23] ;
 wire \soc_inst.cpu_core.register_file.registers[12][24] ;
 wire \soc_inst.cpu_core.register_file.registers[12][25] ;
 wire \soc_inst.cpu_core.register_file.registers[12][26] ;
 wire \soc_inst.cpu_core.register_file.registers[12][27] ;
 wire \soc_inst.cpu_core.register_file.registers[12][28] ;
 wire \soc_inst.cpu_core.register_file.registers[12][29] ;
 wire \soc_inst.cpu_core.register_file.registers[12][2] ;
 wire \soc_inst.cpu_core.register_file.registers[12][30] ;
 wire \soc_inst.cpu_core.register_file.registers[12][31] ;
 wire \soc_inst.cpu_core.register_file.registers[12][3] ;
 wire \soc_inst.cpu_core.register_file.registers[12][4] ;
 wire \soc_inst.cpu_core.register_file.registers[12][5] ;
 wire \soc_inst.cpu_core.register_file.registers[12][6] ;
 wire \soc_inst.cpu_core.register_file.registers[12][7] ;
 wire \soc_inst.cpu_core.register_file.registers[12][8] ;
 wire \soc_inst.cpu_core.register_file.registers[12][9] ;
 wire \soc_inst.cpu_core.register_file.registers[13][0] ;
 wire \soc_inst.cpu_core.register_file.registers[13][10] ;
 wire \soc_inst.cpu_core.register_file.registers[13][11] ;
 wire \soc_inst.cpu_core.register_file.registers[13][12] ;
 wire \soc_inst.cpu_core.register_file.registers[13][13] ;
 wire \soc_inst.cpu_core.register_file.registers[13][14] ;
 wire \soc_inst.cpu_core.register_file.registers[13][15] ;
 wire \soc_inst.cpu_core.register_file.registers[13][16] ;
 wire \soc_inst.cpu_core.register_file.registers[13][17] ;
 wire \soc_inst.cpu_core.register_file.registers[13][18] ;
 wire \soc_inst.cpu_core.register_file.registers[13][19] ;
 wire \soc_inst.cpu_core.register_file.registers[13][1] ;
 wire \soc_inst.cpu_core.register_file.registers[13][20] ;
 wire \soc_inst.cpu_core.register_file.registers[13][21] ;
 wire \soc_inst.cpu_core.register_file.registers[13][22] ;
 wire \soc_inst.cpu_core.register_file.registers[13][23] ;
 wire \soc_inst.cpu_core.register_file.registers[13][24] ;
 wire \soc_inst.cpu_core.register_file.registers[13][25] ;
 wire \soc_inst.cpu_core.register_file.registers[13][26] ;
 wire \soc_inst.cpu_core.register_file.registers[13][27] ;
 wire \soc_inst.cpu_core.register_file.registers[13][28] ;
 wire \soc_inst.cpu_core.register_file.registers[13][29] ;
 wire \soc_inst.cpu_core.register_file.registers[13][2] ;
 wire \soc_inst.cpu_core.register_file.registers[13][30] ;
 wire \soc_inst.cpu_core.register_file.registers[13][31] ;
 wire \soc_inst.cpu_core.register_file.registers[13][3] ;
 wire \soc_inst.cpu_core.register_file.registers[13][4] ;
 wire \soc_inst.cpu_core.register_file.registers[13][5] ;
 wire \soc_inst.cpu_core.register_file.registers[13][6] ;
 wire \soc_inst.cpu_core.register_file.registers[13][7] ;
 wire \soc_inst.cpu_core.register_file.registers[13][8] ;
 wire \soc_inst.cpu_core.register_file.registers[13][9] ;
 wire \soc_inst.cpu_core.register_file.registers[14][0] ;
 wire \soc_inst.cpu_core.register_file.registers[14][10] ;
 wire \soc_inst.cpu_core.register_file.registers[14][11] ;
 wire \soc_inst.cpu_core.register_file.registers[14][12] ;
 wire \soc_inst.cpu_core.register_file.registers[14][13] ;
 wire \soc_inst.cpu_core.register_file.registers[14][14] ;
 wire \soc_inst.cpu_core.register_file.registers[14][15] ;
 wire \soc_inst.cpu_core.register_file.registers[14][16] ;
 wire \soc_inst.cpu_core.register_file.registers[14][17] ;
 wire \soc_inst.cpu_core.register_file.registers[14][18] ;
 wire \soc_inst.cpu_core.register_file.registers[14][19] ;
 wire \soc_inst.cpu_core.register_file.registers[14][1] ;
 wire \soc_inst.cpu_core.register_file.registers[14][20] ;
 wire \soc_inst.cpu_core.register_file.registers[14][21] ;
 wire \soc_inst.cpu_core.register_file.registers[14][22] ;
 wire \soc_inst.cpu_core.register_file.registers[14][23] ;
 wire \soc_inst.cpu_core.register_file.registers[14][24] ;
 wire \soc_inst.cpu_core.register_file.registers[14][25] ;
 wire \soc_inst.cpu_core.register_file.registers[14][26] ;
 wire \soc_inst.cpu_core.register_file.registers[14][27] ;
 wire \soc_inst.cpu_core.register_file.registers[14][28] ;
 wire \soc_inst.cpu_core.register_file.registers[14][29] ;
 wire \soc_inst.cpu_core.register_file.registers[14][2] ;
 wire \soc_inst.cpu_core.register_file.registers[14][30] ;
 wire \soc_inst.cpu_core.register_file.registers[14][31] ;
 wire \soc_inst.cpu_core.register_file.registers[14][3] ;
 wire \soc_inst.cpu_core.register_file.registers[14][4] ;
 wire \soc_inst.cpu_core.register_file.registers[14][5] ;
 wire \soc_inst.cpu_core.register_file.registers[14][6] ;
 wire \soc_inst.cpu_core.register_file.registers[14][7] ;
 wire \soc_inst.cpu_core.register_file.registers[14][8] ;
 wire \soc_inst.cpu_core.register_file.registers[14][9] ;
 wire \soc_inst.cpu_core.register_file.registers[15][0] ;
 wire \soc_inst.cpu_core.register_file.registers[15][10] ;
 wire \soc_inst.cpu_core.register_file.registers[15][11] ;
 wire \soc_inst.cpu_core.register_file.registers[15][12] ;
 wire \soc_inst.cpu_core.register_file.registers[15][13] ;
 wire \soc_inst.cpu_core.register_file.registers[15][14] ;
 wire \soc_inst.cpu_core.register_file.registers[15][15] ;
 wire \soc_inst.cpu_core.register_file.registers[15][16] ;
 wire \soc_inst.cpu_core.register_file.registers[15][17] ;
 wire \soc_inst.cpu_core.register_file.registers[15][18] ;
 wire \soc_inst.cpu_core.register_file.registers[15][19] ;
 wire \soc_inst.cpu_core.register_file.registers[15][1] ;
 wire \soc_inst.cpu_core.register_file.registers[15][20] ;
 wire \soc_inst.cpu_core.register_file.registers[15][21] ;
 wire \soc_inst.cpu_core.register_file.registers[15][22] ;
 wire \soc_inst.cpu_core.register_file.registers[15][23] ;
 wire \soc_inst.cpu_core.register_file.registers[15][24] ;
 wire \soc_inst.cpu_core.register_file.registers[15][25] ;
 wire \soc_inst.cpu_core.register_file.registers[15][26] ;
 wire \soc_inst.cpu_core.register_file.registers[15][27] ;
 wire \soc_inst.cpu_core.register_file.registers[15][28] ;
 wire \soc_inst.cpu_core.register_file.registers[15][29] ;
 wire \soc_inst.cpu_core.register_file.registers[15][2] ;
 wire \soc_inst.cpu_core.register_file.registers[15][30] ;
 wire \soc_inst.cpu_core.register_file.registers[15][31] ;
 wire \soc_inst.cpu_core.register_file.registers[15][3] ;
 wire \soc_inst.cpu_core.register_file.registers[15][4] ;
 wire \soc_inst.cpu_core.register_file.registers[15][5] ;
 wire \soc_inst.cpu_core.register_file.registers[15][6] ;
 wire \soc_inst.cpu_core.register_file.registers[15][7] ;
 wire \soc_inst.cpu_core.register_file.registers[15][8] ;
 wire \soc_inst.cpu_core.register_file.registers[15][9] ;
 wire \soc_inst.cpu_core.register_file.registers[1][0] ;
 wire \soc_inst.cpu_core.register_file.registers[1][10] ;
 wire \soc_inst.cpu_core.register_file.registers[1][11] ;
 wire \soc_inst.cpu_core.register_file.registers[1][12] ;
 wire \soc_inst.cpu_core.register_file.registers[1][13] ;
 wire \soc_inst.cpu_core.register_file.registers[1][14] ;
 wire \soc_inst.cpu_core.register_file.registers[1][15] ;
 wire \soc_inst.cpu_core.register_file.registers[1][16] ;
 wire \soc_inst.cpu_core.register_file.registers[1][17] ;
 wire \soc_inst.cpu_core.register_file.registers[1][18] ;
 wire \soc_inst.cpu_core.register_file.registers[1][19] ;
 wire \soc_inst.cpu_core.register_file.registers[1][1] ;
 wire \soc_inst.cpu_core.register_file.registers[1][20] ;
 wire \soc_inst.cpu_core.register_file.registers[1][21] ;
 wire \soc_inst.cpu_core.register_file.registers[1][22] ;
 wire \soc_inst.cpu_core.register_file.registers[1][23] ;
 wire \soc_inst.cpu_core.register_file.registers[1][24] ;
 wire \soc_inst.cpu_core.register_file.registers[1][25] ;
 wire \soc_inst.cpu_core.register_file.registers[1][26] ;
 wire \soc_inst.cpu_core.register_file.registers[1][27] ;
 wire \soc_inst.cpu_core.register_file.registers[1][28] ;
 wire \soc_inst.cpu_core.register_file.registers[1][29] ;
 wire \soc_inst.cpu_core.register_file.registers[1][2] ;
 wire \soc_inst.cpu_core.register_file.registers[1][30] ;
 wire \soc_inst.cpu_core.register_file.registers[1][31] ;
 wire \soc_inst.cpu_core.register_file.registers[1][3] ;
 wire \soc_inst.cpu_core.register_file.registers[1][4] ;
 wire \soc_inst.cpu_core.register_file.registers[1][5] ;
 wire \soc_inst.cpu_core.register_file.registers[1][6] ;
 wire \soc_inst.cpu_core.register_file.registers[1][7] ;
 wire \soc_inst.cpu_core.register_file.registers[1][8] ;
 wire \soc_inst.cpu_core.register_file.registers[1][9] ;
 wire \soc_inst.cpu_core.register_file.registers[2][0] ;
 wire \soc_inst.cpu_core.register_file.registers[2][10] ;
 wire \soc_inst.cpu_core.register_file.registers[2][11] ;
 wire \soc_inst.cpu_core.register_file.registers[2][12] ;
 wire \soc_inst.cpu_core.register_file.registers[2][13] ;
 wire \soc_inst.cpu_core.register_file.registers[2][14] ;
 wire \soc_inst.cpu_core.register_file.registers[2][15] ;
 wire \soc_inst.cpu_core.register_file.registers[2][16] ;
 wire \soc_inst.cpu_core.register_file.registers[2][17] ;
 wire \soc_inst.cpu_core.register_file.registers[2][18] ;
 wire \soc_inst.cpu_core.register_file.registers[2][19] ;
 wire \soc_inst.cpu_core.register_file.registers[2][1] ;
 wire \soc_inst.cpu_core.register_file.registers[2][20] ;
 wire \soc_inst.cpu_core.register_file.registers[2][21] ;
 wire \soc_inst.cpu_core.register_file.registers[2][22] ;
 wire \soc_inst.cpu_core.register_file.registers[2][23] ;
 wire \soc_inst.cpu_core.register_file.registers[2][24] ;
 wire \soc_inst.cpu_core.register_file.registers[2][25] ;
 wire \soc_inst.cpu_core.register_file.registers[2][26] ;
 wire \soc_inst.cpu_core.register_file.registers[2][27] ;
 wire \soc_inst.cpu_core.register_file.registers[2][28] ;
 wire \soc_inst.cpu_core.register_file.registers[2][29] ;
 wire \soc_inst.cpu_core.register_file.registers[2][2] ;
 wire \soc_inst.cpu_core.register_file.registers[2][30] ;
 wire \soc_inst.cpu_core.register_file.registers[2][31] ;
 wire \soc_inst.cpu_core.register_file.registers[2][3] ;
 wire \soc_inst.cpu_core.register_file.registers[2][4] ;
 wire \soc_inst.cpu_core.register_file.registers[2][5] ;
 wire \soc_inst.cpu_core.register_file.registers[2][6] ;
 wire \soc_inst.cpu_core.register_file.registers[2][7] ;
 wire \soc_inst.cpu_core.register_file.registers[2][8] ;
 wire \soc_inst.cpu_core.register_file.registers[2][9] ;
 wire \soc_inst.cpu_core.register_file.registers[3][0] ;
 wire \soc_inst.cpu_core.register_file.registers[3][10] ;
 wire \soc_inst.cpu_core.register_file.registers[3][11] ;
 wire \soc_inst.cpu_core.register_file.registers[3][12] ;
 wire \soc_inst.cpu_core.register_file.registers[3][13] ;
 wire \soc_inst.cpu_core.register_file.registers[3][14] ;
 wire \soc_inst.cpu_core.register_file.registers[3][15] ;
 wire \soc_inst.cpu_core.register_file.registers[3][16] ;
 wire \soc_inst.cpu_core.register_file.registers[3][17] ;
 wire \soc_inst.cpu_core.register_file.registers[3][18] ;
 wire \soc_inst.cpu_core.register_file.registers[3][19] ;
 wire \soc_inst.cpu_core.register_file.registers[3][1] ;
 wire \soc_inst.cpu_core.register_file.registers[3][20] ;
 wire \soc_inst.cpu_core.register_file.registers[3][21] ;
 wire \soc_inst.cpu_core.register_file.registers[3][22] ;
 wire \soc_inst.cpu_core.register_file.registers[3][23] ;
 wire \soc_inst.cpu_core.register_file.registers[3][24] ;
 wire \soc_inst.cpu_core.register_file.registers[3][25] ;
 wire \soc_inst.cpu_core.register_file.registers[3][26] ;
 wire \soc_inst.cpu_core.register_file.registers[3][27] ;
 wire \soc_inst.cpu_core.register_file.registers[3][28] ;
 wire \soc_inst.cpu_core.register_file.registers[3][29] ;
 wire \soc_inst.cpu_core.register_file.registers[3][2] ;
 wire \soc_inst.cpu_core.register_file.registers[3][30] ;
 wire \soc_inst.cpu_core.register_file.registers[3][31] ;
 wire \soc_inst.cpu_core.register_file.registers[3][3] ;
 wire \soc_inst.cpu_core.register_file.registers[3][4] ;
 wire \soc_inst.cpu_core.register_file.registers[3][5] ;
 wire \soc_inst.cpu_core.register_file.registers[3][6] ;
 wire \soc_inst.cpu_core.register_file.registers[3][7] ;
 wire \soc_inst.cpu_core.register_file.registers[3][8] ;
 wire \soc_inst.cpu_core.register_file.registers[3][9] ;
 wire \soc_inst.cpu_core.register_file.registers[4][0] ;
 wire \soc_inst.cpu_core.register_file.registers[4][10] ;
 wire \soc_inst.cpu_core.register_file.registers[4][11] ;
 wire \soc_inst.cpu_core.register_file.registers[4][12] ;
 wire \soc_inst.cpu_core.register_file.registers[4][13] ;
 wire \soc_inst.cpu_core.register_file.registers[4][14] ;
 wire \soc_inst.cpu_core.register_file.registers[4][15] ;
 wire \soc_inst.cpu_core.register_file.registers[4][16] ;
 wire \soc_inst.cpu_core.register_file.registers[4][17] ;
 wire \soc_inst.cpu_core.register_file.registers[4][18] ;
 wire \soc_inst.cpu_core.register_file.registers[4][19] ;
 wire \soc_inst.cpu_core.register_file.registers[4][1] ;
 wire \soc_inst.cpu_core.register_file.registers[4][20] ;
 wire \soc_inst.cpu_core.register_file.registers[4][21] ;
 wire \soc_inst.cpu_core.register_file.registers[4][22] ;
 wire \soc_inst.cpu_core.register_file.registers[4][23] ;
 wire \soc_inst.cpu_core.register_file.registers[4][24] ;
 wire \soc_inst.cpu_core.register_file.registers[4][25] ;
 wire \soc_inst.cpu_core.register_file.registers[4][26] ;
 wire \soc_inst.cpu_core.register_file.registers[4][27] ;
 wire \soc_inst.cpu_core.register_file.registers[4][28] ;
 wire \soc_inst.cpu_core.register_file.registers[4][29] ;
 wire \soc_inst.cpu_core.register_file.registers[4][2] ;
 wire \soc_inst.cpu_core.register_file.registers[4][30] ;
 wire \soc_inst.cpu_core.register_file.registers[4][31] ;
 wire \soc_inst.cpu_core.register_file.registers[4][3] ;
 wire \soc_inst.cpu_core.register_file.registers[4][4] ;
 wire \soc_inst.cpu_core.register_file.registers[4][5] ;
 wire \soc_inst.cpu_core.register_file.registers[4][6] ;
 wire \soc_inst.cpu_core.register_file.registers[4][7] ;
 wire \soc_inst.cpu_core.register_file.registers[4][8] ;
 wire \soc_inst.cpu_core.register_file.registers[4][9] ;
 wire \soc_inst.cpu_core.register_file.registers[5][0] ;
 wire \soc_inst.cpu_core.register_file.registers[5][10] ;
 wire \soc_inst.cpu_core.register_file.registers[5][11] ;
 wire \soc_inst.cpu_core.register_file.registers[5][12] ;
 wire \soc_inst.cpu_core.register_file.registers[5][13] ;
 wire \soc_inst.cpu_core.register_file.registers[5][14] ;
 wire \soc_inst.cpu_core.register_file.registers[5][15] ;
 wire \soc_inst.cpu_core.register_file.registers[5][16] ;
 wire \soc_inst.cpu_core.register_file.registers[5][17] ;
 wire \soc_inst.cpu_core.register_file.registers[5][18] ;
 wire \soc_inst.cpu_core.register_file.registers[5][19] ;
 wire \soc_inst.cpu_core.register_file.registers[5][1] ;
 wire \soc_inst.cpu_core.register_file.registers[5][20] ;
 wire \soc_inst.cpu_core.register_file.registers[5][21] ;
 wire \soc_inst.cpu_core.register_file.registers[5][22] ;
 wire \soc_inst.cpu_core.register_file.registers[5][23] ;
 wire \soc_inst.cpu_core.register_file.registers[5][24] ;
 wire \soc_inst.cpu_core.register_file.registers[5][25] ;
 wire \soc_inst.cpu_core.register_file.registers[5][26] ;
 wire \soc_inst.cpu_core.register_file.registers[5][27] ;
 wire \soc_inst.cpu_core.register_file.registers[5][28] ;
 wire \soc_inst.cpu_core.register_file.registers[5][29] ;
 wire \soc_inst.cpu_core.register_file.registers[5][2] ;
 wire \soc_inst.cpu_core.register_file.registers[5][30] ;
 wire \soc_inst.cpu_core.register_file.registers[5][31] ;
 wire \soc_inst.cpu_core.register_file.registers[5][3] ;
 wire \soc_inst.cpu_core.register_file.registers[5][4] ;
 wire \soc_inst.cpu_core.register_file.registers[5][5] ;
 wire \soc_inst.cpu_core.register_file.registers[5][6] ;
 wire \soc_inst.cpu_core.register_file.registers[5][7] ;
 wire \soc_inst.cpu_core.register_file.registers[5][8] ;
 wire \soc_inst.cpu_core.register_file.registers[5][9] ;
 wire \soc_inst.cpu_core.register_file.registers[6][0] ;
 wire \soc_inst.cpu_core.register_file.registers[6][10] ;
 wire \soc_inst.cpu_core.register_file.registers[6][11] ;
 wire \soc_inst.cpu_core.register_file.registers[6][12] ;
 wire \soc_inst.cpu_core.register_file.registers[6][13] ;
 wire \soc_inst.cpu_core.register_file.registers[6][14] ;
 wire \soc_inst.cpu_core.register_file.registers[6][15] ;
 wire \soc_inst.cpu_core.register_file.registers[6][16] ;
 wire \soc_inst.cpu_core.register_file.registers[6][17] ;
 wire \soc_inst.cpu_core.register_file.registers[6][18] ;
 wire \soc_inst.cpu_core.register_file.registers[6][19] ;
 wire \soc_inst.cpu_core.register_file.registers[6][1] ;
 wire \soc_inst.cpu_core.register_file.registers[6][20] ;
 wire \soc_inst.cpu_core.register_file.registers[6][21] ;
 wire \soc_inst.cpu_core.register_file.registers[6][22] ;
 wire \soc_inst.cpu_core.register_file.registers[6][23] ;
 wire \soc_inst.cpu_core.register_file.registers[6][24] ;
 wire \soc_inst.cpu_core.register_file.registers[6][25] ;
 wire \soc_inst.cpu_core.register_file.registers[6][26] ;
 wire \soc_inst.cpu_core.register_file.registers[6][27] ;
 wire \soc_inst.cpu_core.register_file.registers[6][28] ;
 wire \soc_inst.cpu_core.register_file.registers[6][29] ;
 wire \soc_inst.cpu_core.register_file.registers[6][2] ;
 wire \soc_inst.cpu_core.register_file.registers[6][30] ;
 wire \soc_inst.cpu_core.register_file.registers[6][31] ;
 wire \soc_inst.cpu_core.register_file.registers[6][3] ;
 wire \soc_inst.cpu_core.register_file.registers[6][4] ;
 wire \soc_inst.cpu_core.register_file.registers[6][5] ;
 wire \soc_inst.cpu_core.register_file.registers[6][6] ;
 wire \soc_inst.cpu_core.register_file.registers[6][7] ;
 wire \soc_inst.cpu_core.register_file.registers[6][8] ;
 wire \soc_inst.cpu_core.register_file.registers[6][9] ;
 wire \soc_inst.cpu_core.register_file.registers[7][0] ;
 wire \soc_inst.cpu_core.register_file.registers[7][10] ;
 wire \soc_inst.cpu_core.register_file.registers[7][11] ;
 wire \soc_inst.cpu_core.register_file.registers[7][12] ;
 wire \soc_inst.cpu_core.register_file.registers[7][13] ;
 wire \soc_inst.cpu_core.register_file.registers[7][14] ;
 wire \soc_inst.cpu_core.register_file.registers[7][15] ;
 wire \soc_inst.cpu_core.register_file.registers[7][16] ;
 wire \soc_inst.cpu_core.register_file.registers[7][17] ;
 wire \soc_inst.cpu_core.register_file.registers[7][18] ;
 wire \soc_inst.cpu_core.register_file.registers[7][19] ;
 wire \soc_inst.cpu_core.register_file.registers[7][1] ;
 wire \soc_inst.cpu_core.register_file.registers[7][20] ;
 wire \soc_inst.cpu_core.register_file.registers[7][21] ;
 wire \soc_inst.cpu_core.register_file.registers[7][22] ;
 wire \soc_inst.cpu_core.register_file.registers[7][23] ;
 wire \soc_inst.cpu_core.register_file.registers[7][24] ;
 wire \soc_inst.cpu_core.register_file.registers[7][25] ;
 wire \soc_inst.cpu_core.register_file.registers[7][26] ;
 wire \soc_inst.cpu_core.register_file.registers[7][27] ;
 wire \soc_inst.cpu_core.register_file.registers[7][28] ;
 wire \soc_inst.cpu_core.register_file.registers[7][29] ;
 wire \soc_inst.cpu_core.register_file.registers[7][2] ;
 wire \soc_inst.cpu_core.register_file.registers[7][30] ;
 wire \soc_inst.cpu_core.register_file.registers[7][31] ;
 wire \soc_inst.cpu_core.register_file.registers[7][3] ;
 wire \soc_inst.cpu_core.register_file.registers[7][4] ;
 wire \soc_inst.cpu_core.register_file.registers[7][5] ;
 wire \soc_inst.cpu_core.register_file.registers[7][6] ;
 wire \soc_inst.cpu_core.register_file.registers[7][7] ;
 wire \soc_inst.cpu_core.register_file.registers[7][8] ;
 wire \soc_inst.cpu_core.register_file.registers[7][9] ;
 wire \soc_inst.cpu_core.register_file.registers[8][0] ;
 wire \soc_inst.cpu_core.register_file.registers[8][10] ;
 wire \soc_inst.cpu_core.register_file.registers[8][11] ;
 wire \soc_inst.cpu_core.register_file.registers[8][12] ;
 wire \soc_inst.cpu_core.register_file.registers[8][13] ;
 wire \soc_inst.cpu_core.register_file.registers[8][14] ;
 wire \soc_inst.cpu_core.register_file.registers[8][15] ;
 wire \soc_inst.cpu_core.register_file.registers[8][16] ;
 wire \soc_inst.cpu_core.register_file.registers[8][17] ;
 wire \soc_inst.cpu_core.register_file.registers[8][18] ;
 wire \soc_inst.cpu_core.register_file.registers[8][19] ;
 wire \soc_inst.cpu_core.register_file.registers[8][1] ;
 wire \soc_inst.cpu_core.register_file.registers[8][20] ;
 wire \soc_inst.cpu_core.register_file.registers[8][21] ;
 wire \soc_inst.cpu_core.register_file.registers[8][22] ;
 wire \soc_inst.cpu_core.register_file.registers[8][23] ;
 wire \soc_inst.cpu_core.register_file.registers[8][24] ;
 wire \soc_inst.cpu_core.register_file.registers[8][25] ;
 wire \soc_inst.cpu_core.register_file.registers[8][26] ;
 wire \soc_inst.cpu_core.register_file.registers[8][27] ;
 wire \soc_inst.cpu_core.register_file.registers[8][28] ;
 wire \soc_inst.cpu_core.register_file.registers[8][29] ;
 wire \soc_inst.cpu_core.register_file.registers[8][2] ;
 wire \soc_inst.cpu_core.register_file.registers[8][30] ;
 wire \soc_inst.cpu_core.register_file.registers[8][31] ;
 wire \soc_inst.cpu_core.register_file.registers[8][3] ;
 wire \soc_inst.cpu_core.register_file.registers[8][4] ;
 wire \soc_inst.cpu_core.register_file.registers[8][5] ;
 wire \soc_inst.cpu_core.register_file.registers[8][6] ;
 wire \soc_inst.cpu_core.register_file.registers[8][7] ;
 wire \soc_inst.cpu_core.register_file.registers[8][8] ;
 wire \soc_inst.cpu_core.register_file.registers[8][9] ;
 wire \soc_inst.cpu_core.register_file.registers[9][0] ;
 wire \soc_inst.cpu_core.register_file.registers[9][10] ;
 wire \soc_inst.cpu_core.register_file.registers[9][11] ;
 wire \soc_inst.cpu_core.register_file.registers[9][12] ;
 wire \soc_inst.cpu_core.register_file.registers[9][13] ;
 wire \soc_inst.cpu_core.register_file.registers[9][14] ;
 wire \soc_inst.cpu_core.register_file.registers[9][15] ;
 wire \soc_inst.cpu_core.register_file.registers[9][16] ;
 wire \soc_inst.cpu_core.register_file.registers[9][17] ;
 wire \soc_inst.cpu_core.register_file.registers[9][18] ;
 wire \soc_inst.cpu_core.register_file.registers[9][19] ;
 wire \soc_inst.cpu_core.register_file.registers[9][1] ;
 wire \soc_inst.cpu_core.register_file.registers[9][20] ;
 wire \soc_inst.cpu_core.register_file.registers[9][21] ;
 wire \soc_inst.cpu_core.register_file.registers[9][22] ;
 wire \soc_inst.cpu_core.register_file.registers[9][23] ;
 wire \soc_inst.cpu_core.register_file.registers[9][24] ;
 wire \soc_inst.cpu_core.register_file.registers[9][25] ;
 wire \soc_inst.cpu_core.register_file.registers[9][26] ;
 wire \soc_inst.cpu_core.register_file.registers[9][27] ;
 wire \soc_inst.cpu_core.register_file.registers[9][28] ;
 wire \soc_inst.cpu_core.register_file.registers[9][29] ;
 wire \soc_inst.cpu_core.register_file.registers[9][2] ;
 wire \soc_inst.cpu_core.register_file.registers[9][30] ;
 wire \soc_inst.cpu_core.register_file.registers[9][31] ;
 wire \soc_inst.cpu_core.register_file.registers[9][3] ;
 wire \soc_inst.cpu_core.register_file.registers[9][4] ;
 wire \soc_inst.cpu_core.register_file.registers[9][5] ;
 wire \soc_inst.cpu_core.register_file.registers[9][6] ;
 wire \soc_inst.cpu_core.register_file.registers[9][7] ;
 wire \soc_inst.cpu_core.register_file.registers[9][8] ;
 wire \soc_inst.cpu_core.register_file.registers[9][9] ;
 wire \soc_inst.flash_cs_n ;
 wire \soc_inst.gpio_inst.gpio_out[0] ;
 wire \soc_inst.gpio_inst.gpio_out[1] ;
 wire \soc_inst.gpio_inst.gpio_out[2] ;
 wire \soc_inst.gpio_inst.gpio_out[3] ;
 wire \soc_inst.gpio_inst.gpio_out[4] ;
 wire \soc_inst.gpio_inst.gpio_out[5] ;
 wire \soc_inst.gpio_inst.gpio_sync1[0] ;
 wire \soc_inst.gpio_inst.gpio_sync1[1] ;
 wire \soc_inst.gpio_inst.gpio_sync1[2] ;
 wire \soc_inst.gpio_inst.gpio_sync1[3] ;
 wire \soc_inst.gpio_inst.gpio_sync1[4] ;
 wire \soc_inst.gpio_inst.gpio_sync1[5] ;
 wire \soc_inst.gpio_inst.gpio_sync1[6] ;
 wire \soc_inst.gpio_inst.gpio_sync2[0] ;
 wire \soc_inst.gpio_inst.gpio_sync2[1] ;
 wire \soc_inst.gpio_inst.gpio_sync2[2] ;
 wire \soc_inst.gpio_inst.gpio_sync2[3] ;
 wire \soc_inst.gpio_inst.gpio_sync2[4] ;
 wire \soc_inst.gpio_inst.gpio_sync2[5] ;
 wire \soc_inst.gpio_inst.gpio_sync2[6] ;
 wire \soc_inst.gpio_inst.int_en_reg[0] ;
 wire \soc_inst.gpio_inst.int_en_reg[1] ;
 wire \soc_inst.gpio_inst.int_en_reg[2] ;
 wire \soc_inst.gpio_inst.int_en_reg[3] ;
 wire \soc_inst.gpio_inst.int_en_reg[4] ;
 wire \soc_inst.gpio_inst.int_en_reg[5] ;
 wire \soc_inst.gpio_inst.int_en_reg[6] ;
 wire \soc_inst.gpio_inst.int_pend_reg[0] ;
 wire \soc_inst.gpio_inst.int_pend_reg[1] ;
 wire \soc_inst.gpio_inst.int_pend_reg[2] ;
 wire \soc_inst.gpio_inst.int_pend_reg[3] ;
 wire \soc_inst.gpio_inst.int_pend_reg[4] ;
 wire \soc_inst.gpio_inst.int_pend_reg[5] ;
 wire \soc_inst.gpio_inst.int_pend_reg[6] ;
 wire \soc_inst.i2c_ena ;
 wire \soc_inst.i2c_inst.ack_enable ;
 wire \soc_inst.i2c_inst.ack_received ;
 wire \soc_inst.i2c_inst.arb_lost ;
 wire \soc_inst.i2c_inst.bit_cnt[0] ;
 wire \soc_inst.i2c_inst.bit_cnt[1] ;
 wire \soc_inst.i2c_inst.bit_cnt[2] ;
 wire \soc_inst.i2c_inst.bit_cnt[3] ;
 wire \soc_inst.i2c_inst.clk_cnt[0] ;
 wire \soc_inst.i2c_inst.clk_cnt[1] ;
 wire \soc_inst.i2c_inst.clk_cnt[2] ;
 wire \soc_inst.i2c_inst.clk_cnt[3] ;
 wire \soc_inst.i2c_inst.clk_cnt[4] ;
 wire \soc_inst.i2c_inst.clk_cnt[5] ;
 wire \soc_inst.i2c_inst.clk_cnt[6] ;
 wire \soc_inst.i2c_inst.clk_cnt[7] ;
 wire \soc_inst.i2c_inst.ctrl_reg[2] ;
 wire \soc_inst.i2c_inst.ctrl_reg[4] ;
 wire \soc_inst.i2c_inst.data_reg[0] ;
 wire \soc_inst.i2c_inst.data_reg[1] ;
 wire \soc_inst.i2c_inst.data_reg[2] ;
 wire \soc_inst.i2c_inst.data_reg[3] ;
 wire \soc_inst.i2c_inst.data_reg[4] ;
 wire \soc_inst.i2c_inst.data_reg[5] ;
 wire \soc_inst.i2c_inst.data_reg[6] ;
 wire \soc_inst.i2c_inst.data_reg[7] ;
 wire \soc_inst.i2c_inst.prescale_reg[5] ;
 wire \soc_inst.i2c_inst.prescale_reg[6] ;
 wire \soc_inst.i2c_inst.restart_pending ;
 wire \soc_inst.i2c_inst.shift_reg[0] ;
 wire \soc_inst.i2c_inst.shift_reg[1] ;
 wire \soc_inst.i2c_inst.shift_reg[2] ;
 wire \soc_inst.i2c_inst.shift_reg[3] ;
 wire \soc_inst.i2c_inst.shift_reg[4] ;
 wire \soc_inst.i2c_inst.shift_reg[5] ;
 wire \soc_inst.i2c_inst.shift_reg[6] ;
 wire \soc_inst.i2c_inst.shift_reg[7] ;
 wire \soc_inst.i2c_inst.start_pending ;
 wire \soc_inst.i2c_inst.state[0] ;
 wire \soc_inst.i2c_inst.state[1] ;
 wire \soc_inst.i2c_inst.state[2] ;
 wire \soc_inst.i2c_inst.state[3] ;
 wire \soc_inst.i2c_inst.status_reg[0] ;
 wire \soc_inst.i2c_inst.status_reg[1] ;
 wire \soc_inst.i2c_inst.status_reg[2] ;
 wire \soc_inst.i2c_inst.status_reg[3] ;
 wire \soc_inst.i2c_inst.stop_pending ;
 wire \soc_inst.i2c_inst.transfer_done ;
 wire \soc_inst.mem_ctrl.access_state[1] ;
 wire \soc_inst.mem_ctrl.access_state[2] ;
 wire \soc_inst.mem_ctrl.access_state[3] ;
 wire \soc_inst.mem_ctrl.access_state[4] ;
 wire \soc_inst.mem_ctrl.instr_ready_reg ;
 wire \soc_inst.mem_ctrl.next_instr_addr[0] ;
 wire \soc_inst.mem_ctrl.next_instr_data[0] ;
 wire \soc_inst.mem_ctrl.next_instr_data[10] ;
 wire \soc_inst.mem_ctrl.next_instr_data[11] ;
 wire \soc_inst.mem_ctrl.next_instr_data[12] ;
 wire \soc_inst.mem_ctrl.next_instr_data[13] ;
 wire \soc_inst.mem_ctrl.next_instr_data[14] ;
 wire \soc_inst.mem_ctrl.next_instr_data[15] ;
 wire \soc_inst.mem_ctrl.next_instr_data[16] ;
 wire \soc_inst.mem_ctrl.next_instr_data[17] ;
 wire \soc_inst.mem_ctrl.next_instr_data[18] ;
 wire \soc_inst.mem_ctrl.next_instr_data[19] ;
 wire \soc_inst.mem_ctrl.next_instr_data[1] ;
 wire \soc_inst.mem_ctrl.next_instr_data[20] ;
 wire \soc_inst.mem_ctrl.next_instr_data[21] ;
 wire \soc_inst.mem_ctrl.next_instr_data[22] ;
 wire \soc_inst.mem_ctrl.next_instr_data[23] ;
 wire \soc_inst.mem_ctrl.next_instr_data[24] ;
 wire \soc_inst.mem_ctrl.next_instr_data[25] ;
 wire \soc_inst.mem_ctrl.next_instr_data[26] ;
 wire \soc_inst.mem_ctrl.next_instr_data[27] ;
 wire \soc_inst.mem_ctrl.next_instr_data[28] ;
 wire \soc_inst.mem_ctrl.next_instr_data[29] ;
 wire \soc_inst.mem_ctrl.next_instr_data[2] ;
 wire \soc_inst.mem_ctrl.next_instr_data[30] ;
 wire \soc_inst.mem_ctrl.next_instr_data[31] ;
 wire \soc_inst.mem_ctrl.next_instr_data[3] ;
 wire \soc_inst.mem_ctrl.next_instr_data[4] ;
 wire \soc_inst.mem_ctrl.next_instr_data[5] ;
 wire \soc_inst.mem_ctrl.next_instr_data[6] ;
 wire \soc_inst.mem_ctrl.next_instr_data[7] ;
 wire \soc_inst.mem_ctrl.next_instr_data[8] ;
 wire \soc_inst.mem_ctrl.next_instr_data[9] ;
 wire \soc_inst.mem_ctrl.next_instr_ready_reg ;
 wire \soc_inst.mem_ctrl.ram_cs_n ;
 wire \soc_inst.mem_ctrl.spi_addr[10] ;
 wire \soc_inst.mem_ctrl.spi_addr[11] ;
 wire \soc_inst.mem_ctrl.spi_addr[12] ;
 wire \soc_inst.mem_ctrl.spi_addr[13] ;
 wire \soc_inst.mem_ctrl.spi_addr[14] ;
 wire \soc_inst.mem_ctrl.spi_addr[15] ;
 wire \soc_inst.mem_ctrl.spi_addr[16] ;
 wire \soc_inst.mem_ctrl.spi_addr[17] ;
 wire \soc_inst.mem_ctrl.spi_addr[18] ;
 wire \soc_inst.mem_ctrl.spi_addr[19] ;
 wire \soc_inst.mem_ctrl.spi_addr[1] ;
 wire \soc_inst.mem_ctrl.spi_addr[20] ;
 wire \soc_inst.mem_ctrl.spi_addr[21] ;
 wire \soc_inst.mem_ctrl.spi_addr[22] ;
 wire \soc_inst.mem_ctrl.spi_addr[23] ;
 wire \soc_inst.mem_ctrl.spi_addr[2] ;
 wire \soc_inst.mem_ctrl.spi_addr[3] ;
 wire \soc_inst.mem_ctrl.spi_addr[4] ;
 wire \soc_inst.mem_ctrl.spi_addr[5] ;
 wire \soc_inst.mem_ctrl.spi_addr[6] ;
 wire \soc_inst.mem_ctrl.spi_addr[7] ;
 wire \soc_inst.mem_ctrl.spi_addr[8] ;
 wire \soc_inst.mem_ctrl.spi_addr[9] ;
 wire \soc_inst.mem_ctrl.spi_data_in[0] ;
 wire \soc_inst.mem_ctrl.spi_data_in[10] ;
 wire \soc_inst.mem_ctrl.spi_data_in[11] ;
 wire \soc_inst.mem_ctrl.spi_data_in[12] ;
 wire \soc_inst.mem_ctrl.spi_data_in[13] ;
 wire \soc_inst.mem_ctrl.spi_data_in[14] ;
 wire \soc_inst.mem_ctrl.spi_data_in[15] ;
 wire \soc_inst.mem_ctrl.spi_data_in[16] ;
 wire \soc_inst.mem_ctrl.spi_data_in[17] ;
 wire \soc_inst.mem_ctrl.spi_data_in[18] ;
 wire \soc_inst.mem_ctrl.spi_data_in[19] ;
 wire \soc_inst.mem_ctrl.spi_data_in[1] ;
 wire \soc_inst.mem_ctrl.spi_data_in[20] ;
 wire \soc_inst.mem_ctrl.spi_data_in[21] ;
 wire \soc_inst.mem_ctrl.spi_data_in[22] ;
 wire \soc_inst.mem_ctrl.spi_data_in[23] ;
 wire \soc_inst.mem_ctrl.spi_data_in[24] ;
 wire \soc_inst.mem_ctrl.spi_data_in[25] ;
 wire \soc_inst.mem_ctrl.spi_data_in[26] ;
 wire \soc_inst.mem_ctrl.spi_data_in[27] ;
 wire \soc_inst.mem_ctrl.spi_data_in[28] ;
 wire \soc_inst.mem_ctrl.spi_data_in[29] ;
 wire \soc_inst.mem_ctrl.spi_data_in[2] ;
 wire \soc_inst.mem_ctrl.spi_data_in[30] ;
 wire \soc_inst.mem_ctrl.spi_data_in[31] ;
 wire \soc_inst.mem_ctrl.spi_data_in[3] ;
 wire \soc_inst.mem_ctrl.spi_data_in[4] ;
 wire \soc_inst.mem_ctrl.spi_data_in[5] ;
 wire \soc_inst.mem_ctrl.spi_data_in[6] ;
 wire \soc_inst.mem_ctrl.spi_data_in[7] ;
 wire \soc_inst.mem_ctrl.spi_data_in[8] ;
 wire \soc_inst.mem_ctrl.spi_data_in[9] ;
 wire \soc_inst.mem_ctrl.spi_data_len[3] ;
 wire \soc_inst.mem_ctrl.spi_data_len[4] ;
 wire \soc_inst.mem_ctrl.spi_data_len[5] ;
 wire \soc_inst.mem_ctrl.spi_data_out[0] ;
 wire \soc_inst.mem_ctrl.spi_data_out[10] ;
 wire \soc_inst.mem_ctrl.spi_data_out[11] ;
 wire \soc_inst.mem_ctrl.spi_data_out[12] ;
 wire \soc_inst.mem_ctrl.spi_data_out[13] ;
 wire \soc_inst.mem_ctrl.spi_data_out[14] ;
 wire \soc_inst.mem_ctrl.spi_data_out[15] ;
 wire \soc_inst.mem_ctrl.spi_data_out[16] ;
 wire \soc_inst.mem_ctrl.spi_data_out[17] ;
 wire \soc_inst.mem_ctrl.spi_data_out[18] ;
 wire \soc_inst.mem_ctrl.spi_data_out[19] ;
 wire \soc_inst.mem_ctrl.spi_data_out[1] ;
 wire \soc_inst.mem_ctrl.spi_data_out[20] ;
 wire \soc_inst.mem_ctrl.spi_data_out[21] ;
 wire \soc_inst.mem_ctrl.spi_data_out[22] ;
 wire \soc_inst.mem_ctrl.spi_data_out[23] ;
 wire \soc_inst.mem_ctrl.spi_data_out[24] ;
 wire \soc_inst.mem_ctrl.spi_data_out[25] ;
 wire \soc_inst.mem_ctrl.spi_data_out[26] ;
 wire \soc_inst.mem_ctrl.spi_data_out[27] ;
 wire \soc_inst.mem_ctrl.spi_data_out[28] ;
 wire \soc_inst.mem_ctrl.spi_data_out[29] ;
 wire \soc_inst.mem_ctrl.spi_data_out[2] ;
 wire \soc_inst.mem_ctrl.spi_data_out[30] ;
 wire \soc_inst.mem_ctrl.spi_data_out[31] ;
 wire \soc_inst.mem_ctrl.spi_data_out[3] ;
 wire \soc_inst.mem_ctrl.spi_data_out[4] ;
 wire \soc_inst.mem_ctrl.spi_data_out[5] ;
 wire \soc_inst.mem_ctrl.spi_data_out[6] ;
 wire \soc_inst.mem_ctrl.spi_data_out[7] ;
 wire \soc_inst.mem_ctrl.spi_data_out[8] ;
 wire \soc_inst.mem_ctrl.spi_data_out[9] ;
 wire \soc_inst.mem_ctrl.spi_done ;
 wire \soc_inst.mem_ctrl.spi_is_instr ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.flash_in_cont_mode ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.initialized ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.is_write_op ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.ram_in_quad_mode ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[12] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[23] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[28] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[30] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[31] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[18] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[25] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.start ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.stop ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.write_enable ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.write_mosi ;
 wire \soc_inst.mem_ctrl.spi_read_enable ;
 wire \soc_inst.pwm_ena[0] ;
 wire \soc_inst.pwm_ena[1] ;
 wire \soc_inst.pwm_inst.channel_counter[0][0] ;
 wire \soc_inst.pwm_inst.channel_counter[0][10] ;
 wire \soc_inst.pwm_inst.channel_counter[0][11] ;
 wire \soc_inst.pwm_inst.channel_counter[0][12] ;
 wire \soc_inst.pwm_inst.channel_counter[0][13] ;
 wire \soc_inst.pwm_inst.channel_counter[0][14] ;
 wire \soc_inst.pwm_inst.channel_counter[0][15] ;
 wire \soc_inst.pwm_inst.channel_counter[0][1] ;
 wire \soc_inst.pwm_inst.channel_counter[0][2] ;
 wire \soc_inst.pwm_inst.channel_counter[0][3] ;
 wire \soc_inst.pwm_inst.channel_counter[0][4] ;
 wire \soc_inst.pwm_inst.channel_counter[0][5] ;
 wire \soc_inst.pwm_inst.channel_counter[0][6] ;
 wire \soc_inst.pwm_inst.channel_counter[0][7] ;
 wire \soc_inst.pwm_inst.channel_counter[0][8] ;
 wire \soc_inst.pwm_inst.channel_counter[0][9] ;
 wire \soc_inst.pwm_inst.channel_counter[1][0] ;
 wire \soc_inst.pwm_inst.channel_counter[1][10] ;
 wire \soc_inst.pwm_inst.channel_counter[1][11] ;
 wire \soc_inst.pwm_inst.channel_counter[1][12] ;
 wire \soc_inst.pwm_inst.channel_counter[1][13] ;
 wire \soc_inst.pwm_inst.channel_counter[1][14] ;
 wire \soc_inst.pwm_inst.channel_counter[1][15] ;
 wire \soc_inst.pwm_inst.channel_counter[1][1] ;
 wire \soc_inst.pwm_inst.channel_counter[1][2] ;
 wire \soc_inst.pwm_inst.channel_counter[1][3] ;
 wire \soc_inst.pwm_inst.channel_counter[1][4] ;
 wire \soc_inst.pwm_inst.channel_counter[1][5] ;
 wire \soc_inst.pwm_inst.channel_counter[1][6] ;
 wire \soc_inst.pwm_inst.channel_counter[1][7] ;
 wire \soc_inst.pwm_inst.channel_counter[1][8] ;
 wire \soc_inst.pwm_inst.channel_counter[1][9] ;
 wire \soc_inst.pwm_inst.channel_duty[0][0] ;
 wire \soc_inst.pwm_inst.channel_duty[0][10] ;
 wire \soc_inst.pwm_inst.channel_duty[0][11] ;
 wire \soc_inst.pwm_inst.channel_duty[0][12] ;
 wire \soc_inst.pwm_inst.channel_duty[0][13] ;
 wire \soc_inst.pwm_inst.channel_duty[0][14] ;
 wire \soc_inst.pwm_inst.channel_duty[0][15] ;
 wire \soc_inst.pwm_inst.channel_duty[0][1] ;
 wire \soc_inst.pwm_inst.channel_duty[0][2] ;
 wire \soc_inst.pwm_inst.channel_duty[0][3] ;
 wire \soc_inst.pwm_inst.channel_duty[0][4] ;
 wire \soc_inst.pwm_inst.channel_duty[0][5] ;
 wire \soc_inst.pwm_inst.channel_duty[0][6] ;
 wire \soc_inst.pwm_inst.channel_duty[0][7] ;
 wire \soc_inst.pwm_inst.channel_duty[0][8] ;
 wire \soc_inst.pwm_inst.channel_duty[0][9] ;
 wire \soc_inst.pwm_inst.channel_duty[1][0] ;
 wire \soc_inst.pwm_inst.channel_duty[1][10] ;
 wire \soc_inst.pwm_inst.channel_duty[1][11] ;
 wire \soc_inst.pwm_inst.channel_duty[1][12] ;
 wire \soc_inst.pwm_inst.channel_duty[1][13] ;
 wire \soc_inst.pwm_inst.channel_duty[1][14] ;
 wire \soc_inst.pwm_inst.channel_duty[1][15] ;
 wire \soc_inst.pwm_inst.channel_duty[1][1] ;
 wire \soc_inst.pwm_inst.channel_duty[1][2] ;
 wire \soc_inst.pwm_inst.channel_duty[1][3] ;
 wire \soc_inst.pwm_inst.channel_duty[1][4] ;
 wire \soc_inst.pwm_inst.channel_duty[1][5] ;
 wire \soc_inst.pwm_inst.channel_duty[1][6] ;
 wire \soc_inst.pwm_inst.channel_duty[1][7] ;
 wire \soc_inst.pwm_inst.channel_duty[1][8] ;
 wire \soc_inst.pwm_inst.channel_duty[1][9] ;
 wire \soc_inst.spi_ena ;
 wire \soc_inst.spi_inst.bit_counter[0] ;
 wire \soc_inst.spi_inst.bit_counter[1] ;
 wire \soc_inst.spi_inst.bit_counter[2] ;
 wire \soc_inst.spi_inst.bit_counter[3] ;
 wire \soc_inst.spi_inst.bit_counter[4] ;
 wire \soc_inst.spi_inst.bit_counter[5] ;
 wire \soc_inst.spi_inst.busy ;
 wire \soc_inst.spi_inst.clk_counter[0] ;
 wire \soc_inst.spi_inst.clk_counter[1] ;
 wire \soc_inst.spi_inst.clk_counter[2] ;
 wire \soc_inst.spi_inst.clk_counter[3] ;
 wire \soc_inst.spi_inst.clk_counter[4] ;
 wire \soc_inst.spi_inst.clk_counter[5] ;
 wire \soc_inst.spi_inst.clk_counter[6] ;
 wire \soc_inst.spi_inst.clk_counter[7] ;
 wire \soc_inst.spi_inst.clock_divider[5] ;
 wire \soc_inst.spi_inst.clock_divider[6] ;
 wire \soc_inst.spi_inst.clock_divider[7] ;
 wire \soc_inst.spi_inst.cpha ;
 wire \soc_inst.spi_inst.cpol ;
 wire \soc_inst.spi_inst.done ;
 wire \soc_inst.spi_inst.len_sel[0] ;
 wire \soc_inst.spi_inst.len_sel[1] ;
 wire \soc_inst.spi_inst.next_state[0] ;
 wire \soc_inst.spi_inst.next_state[1] ;
 wire \soc_inst.spi_inst.rx_shift_reg[0] ;
 wire \soc_inst.spi_inst.rx_shift_reg[10] ;
 wire \soc_inst.spi_inst.rx_shift_reg[11] ;
 wire \soc_inst.spi_inst.rx_shift_reg[12] ;
 wire \soc_inst.spi_inst.rx_shift_reg[13] ;
 wire \soc_inst.spi_inst.rx_shift_reg[14] ;
 wire \soc_inst.spi_inst.rx_shift_reg[15] ;
 wire \soc_inst.spi_inst.rx_shift_reg[16] ;
 wire \soc_inst.spi_inst.rx_shift_reg[17] ;
 wire \soc_inst.spi_inst.rx_shift_reg[18] ;
 wire \soc_inst.spi_inst.rx_shift_reg[19] ;
 wire \soc_inst.spi_inst.rx_shift_reg[1] ;
 wire \soc_inst.spi_inst.rx_shift_reg[20] ;
 wire \soc_inst.spi_inst.rx_shift_reg[21] ;
 wire \soc_inst.spi_inst.rx_shift_reg[22] ;
 wire \soc_inst.spi_inst.rx_shift_reg[23] ;
 wire \soc_inst.spi_inst.rx_shift_reg[24] ;
 wire \soc_inst.spi_inst.rx_shift_reg[25] ;
 wire \soc_inst.spi_inst.rx_shift_reg[26] ;
 wire \soc_inst.spi_inst.rx_shift_reg[27] ;
 wire \soc_inst.spi_inst.rx_shift_reg[28] ;
 wire \soc_inst.spi_inst.rx_shift_reg[29] ;
 wire \soc_inst.spi_inst.rx_shift_reg[2] ;
 wire \soc_inst.spi_inst.rx_shift_reg[30] ;
 wire \soc_inst.spi_inst.rx_shift_reg[31] ;
 wire \soc_inst.spi_inst.rx_shift_reg[3] ;
 wire \soc_inst.spi_inst.rx_shift_reg[4] ;
 wire \soc_inst.spi_inst.rx_shift_reg[5] ;
 wire \soc_inst.spi_inst.rx_shift_reg[6] ;
 wire \soc_inst.spi_inst.rx_shift_reg[7] ;
 wire \soc_inst.spi_inst.rx_shift_reg[8] ;
 wire \soc_inst.spi_inst.rx_shift_reg[9] ;
 wire \soc_inst.spi_inst.spi_clk_en ;
 wire \soc_inst.spi_inst.spi_mosi ;
 wire \soc_inst.spi_inst.spi_sclk ;
 wire \soc_inst.spi_inst.start_pending ;
 wire \soc_inst.spi_inst.state[0] ;
 wire \soc_inst.spi_inst.state[1] ;
 wire \soc_inst.spi_inst.tx_shift_reg[0] ;
 wire \soc_inst.spi_inst.tx_shift_reg[10] ;
 wire \soc_inst.spi_inst.tx_shift_reg[11] ;
 wire \soc_inst.spi_inst.tx_shift_reg[12] ;
 wire \soc_inst.spi_inst.tx_shift_reg[13] ;
 wire \soc_inst.spi_inst.tx_shift_reg[14] ;
 wire \soc_inst.spi_inst.tx_shift_reg[15] ;
 wire \soc_inst.spi_inst.tx_shift_reg[16] ;
 wire \soc_inst.spi_inst.tx_shift_reg[17] ;
 wire \soc_inst.spi_inst.tx_shift_reg[18] ;
 wire \soc_inst.spi_inst.tx_shift_reg[19] ;
 wire \soc_inst.spi_inst.tx_shift_reg[1] ;
 wire \soc_inst.spi_inst.tx_shift_reg[20] ;
 wire \soc_inst.spi_inst.tx_shift_reg[21] ;
 wire \soc_inst.spi_inst.tx_shift_reg[22] ;
 wire \soc_inst.spi_inst.tx_shift_reg[23] ;
 wire \soc_inst.spi_inst.tx_shift_reg[24] ;
 wire \soc_inst.spi_inst.tx_shift_reg[25] ;
 wire \soc_inst.spi_inst.tx_shift_reg[26] ;
 wire \soc_inst.spi_inst.tx_shift_reg[27] ;
 wire \soc_inst.spi_inst.tx_shift_reg[28] ;
 wire \soc_inst.spi_inst.tx_shift_reg[29] ;
 wire \soc_inst.spi_inst.tx_shift_reg[2] ;
 wire \soc_inst.spi_inst.tx_shift_reg[30] ;
 wire \soc_inst.spi_inst.tx_shift_reg[31] ;
 wire \soc_inst.spi_inst.tx_shift_reg[3] ;
 wire \soc_inst.spi_inst.tx_shift_reg[4] ;
 wire \soc_inst.spi_inst.tx_shift_reg[5] ;
 wire \soc_inst.spi_inst.tx_shift_reg[6] ;
 wire \soc_inst.spi_inst.tx_shift_reg[7] ;
 wire \soc_inst.spi_inst.tx_shift_reg[8] ;
 wire \soc_inst.spi_inst.tx_shift_reg[9] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_sample ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg_0 ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_rx_break_reg ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ;
 wire net77;
 wire net78;
 wire clknet_leaf_0_clk;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0_0_clk;
 wire clknet_6_1_0_clk;
 wire clknet_6_2_0_clk;
 wire clknet_6_3_0_clk;
 wire clknet_6_4_0_clk;
 wire clknet_6_5_0_clk;
 wire clknet_6_6_0_clk;
 wire clknet_6_7_0_clk;
 wire clknet_6_8_0_clk;
 wire clknet_6_9_0_clk;
 wire clknet_6_10_0_clk;
 wire clknet_6_11_0_clk;
 wire clknet_6_12_0_clk;
 wire clknet_6_13_0_clk;
 wire clknet_6_14_0_clk;
 wire clknet_6_15_0_clk;
 wire clknet_6_16_0_clk;
 wire clknet_6_17_0_clk;
 wire clknet_6_18_0_clk;
 wire clknet_6_19_0_clk;
 wire clknet_6_20_0_clk;
 wire clknet_6_21_0_clk;
 wire clknet_6_22_0_clk;
 wire clknet_6_23_0_clk;
 wire clknet_6_24_0_clk;
 wire clknet_6_25_0_clk;
 wire clknet_6_26_0_clk;
 wire clknet_6_27_0_clk;
 wire clknet_6_28_0_clk;
 wire clknet_6_29_0_clk;
 wire clknet_6_30_0_clk;
 wire clknet_6_31_0_clk;
 wire clknet_6_32_0_clk;
 wire clknet_6_33_0_clk;
 wire clknet_6_34_0_clk;
 wire clknet_6_35_0_clk;
 wire clknet_6_36_0_clk;
 wire clknet_6_37_0_clk;
 wire clknet_6_38_0_clk;
 wire clknet_6_39_0_clk;
 wire clknet_6_40_0_clk;
 wire clknet_6_41_0_clk;
 wire clknet_6_42_0_clk;
 wire clknet_6_43_0_clk;
 wire clknet_6_44_0_clk;
 wire clknet_6_45_0_clk;
 wire clknet_6_46_0_clk;
 wire clknet_6_47_0_clk;
 wire clknet_6_48_0_clk;
 wire clknet_6_49_0_clk;
 wire clknet_6_50_0_clk;
 wire clknet_6_51_0_clk;
 wire clknet_6_52_0_clk;
 wire clknet_6_53_0_clk;
 wire clknet_6_54_0_clk;
 wire clknet_6_55_0_clk;
 wire clknet_6_56_0_clk;
 wire clknet_6_57_0_clk;
 wire clknet_6_58_0_clk;
 wire clknet_6_59_0_clk;
 wire clknet_6_60_0_clk;
 wire clknet_6_61_0_clk;
 wire clknet_6_62_0_clk;
 wire clknet_6_63_0_clk;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire [0:0] _10277_;
 wire [0:0] _10278_;
 wire [0:0] _10279_;
 wire [0:0] \soc_inst.gpio_bidir_oe ;
 wire [0:0] \soc_inst.gpio_bidir_out ;
 wire [0:0] \soc_inst.pwm_inst.channel_idx ;
 wire [0:0] \soc_inst.uart_tx ;

 sg13g2_inv_1 _10280_ (.Y(_05373_),
    .A(net1698));
 sg13g2_inv_2 _10281_ (.Y(_05374_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ));
 sg13g2_inv_1 _10282_ (.Y(_05375_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ));
 sg13g2_inv_2 _10283_ (.Y(_05376_),
    .A(net2577));
 sg13g2_inv_1 _10284_ (.Y(_05377_),
    .A(net2597));
 sg13g2_inv_1 _10285_ (.Y(_05378_),
    .A(net1276));
 sg13g2_inv_1 _10286_ (.Y(_05379_),
    .A(net1299));
 sg13g2_inv_1 _10287_ (.Y(_05380_),
    .A(net1991));
 sg13g2_inv_2 _10288_ (.Y(_05381_),
    .A(net597));
 sg13g2_inv_1 _10289_ (.Y(_05382_),
    .A(net655));
 sg13g2_inv_1 _10290_ (.Y(_05383_),
    .A(net1019));
 sg13g2_inv_1 _10291_ (.Y(_05384_),
    .A(net620));
 sg13g2_inv_1 _10292_ (.Y(_05385_),
    .A(net605));
 sg13g2_inv_1 _10293_ (.Y(_05386_),
    .A(net4762));
 sg13g2_inv_1 _10294_ (.Y(_05387_),
    .A(net4758));
 sg13g2_inv_1 _10295_ (.Y(_05388_),
    .A(_00329_));
 sg13g2_inv_2 _10296_ (.Y(_05389_),
    .A(_00328_));
 sg13g2_inv_1 _10297_ (.Y(_05390_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ));
 sg13g2_inv_1 _10298_ (.Y(_05391_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ));
 sg13g2_inv_1 _10299_ (.Y(_05392_),
    .A(net2892));
 sg13g2_inv_1 _10300_ (.Y(_05393_),
    .A(net517));
 sg13g2_inv_1 _10301_ (.Y(_05394_),
    .A(_00324_));
 sg13g2_inv_1 _10302_ (.Y(_05395_),
    .A(_00323_));
 sg13g2_inv_1 _10303_ (.Y(_05396_),
    .A(_00297_));
 sg13g2_inv_1 _10304_ (.Y(_05397_),
    .A(net2074));
 sg13g2_inv_1 _10305_ (.Y(_05398_),
    .A(net2382));
 sg13g2_inv_1 _10306_ (.Y(_05399_),
    .A(_00287_));
 sg13g2_inv_1 _10307_ (.Y(_05400_),
    .A(_00280_));
 sg13g2_inv_1 _10308_ (.Y(_05401_),
    .A(_00279_));
 sg13g2_inv_1 _10309_ (.Y(_05402_),
    .A(_00278_));
 sg13g2_inv_2 _10310_ (.Y(_05403_),
    .A(net603));
 sg13g2_inv_1 _10311_ (.Y(_05404_),
    .A(_00258_));
 sg13g2_inv_1 _10312_ (.Y(_05405_),
    .A(net158));
 sg13g2_inv_1 _10313_ (.Y(_05406_),
    .A(_00220_));
 sg13g2_inv_1 _10314_ (.Y(_05407_),
    .A(_00219_));
 sg13g2_inv_1 _10315_ (.Y(_05408_),
    .A(_00218_));
 sg13g2_inv_1 _10316_ (.Y(_05409_),
    .A(_00217_));
 sg13g2_inv_1 _10317_ (.Y(_00169_),
    .A(net556));
 sg13g2_inv_1 _10318_ (.Y(_05410_),
    .A(net2738));
 sg13g2_inv_1 _10319_ (.Y(_05411_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ));
 sg13g2_inv_2 _10320_ (.Y(_05412_),
    .A(net2776));
 sg13g2_inv_2 _10321_ (.Y(_05413_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ));
 sg13g2_inv_2 _10322_ (.Y(_05414_),
    .A(net2554));
 sg13g2_inv_2 _10323_ (.Y(_05415_),
    .A(net4872));
 sg13g2_inv_2 _10324_ (.Y(_05416_),
    .A(net4866));
 sg13g2_inv_8 _10325_ (.Y(_05417_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ));
 sg13g2_inv_1 _10326_ (.Y(_05418_),
    .A(net2583));
 sg13g2_inv_1 _10327_ (.Y(_05419_),
    .A(net2371));
 sg13g2_inv_2 _10328_ (.Y(_05420_),
    .A(net1807));
 sg13g2_inv_2 _10329_ (.Y(_05421_),
    .A(net2195));
 sg13g2_inv_1 _10330_ (.Y(_05422_),
    .A(net2935));
 sg13g2_inv_2 _10331_ (.Y(_05423_),
    .A(net4787));
 sg13g2_inv_4 _10332_ (.A(net2951),
    .Y(_05424_));
 sg13g2_inv_4 _10333_ (.A(net2489),
    .Y(_05425_));
 sg13g2_inv_1 _10334_ (.Y(_05426_),
    .A(net2515));
 sg13g2_inv_1 _10335_ (.Y(_05427_),
    .A(net2725));
 sg13g2_inv_1 _10336_ (.Y(_05428_),
    .A(net2672));
 sg13g2_inv_1 _10337_ (.Y(_05429_),
    .A(net2791));
 sg13g2_inv_1 _10338_ (.Y(_05430_),
    .A(net2548));
 sg13g2_inv_1 _10339_ (.Y(_05431_),
    .A(net2730));
 sg13g2_inv_1 _10340_ (.Y(_05432_),
    .A(net2433));
 sg13g2_inv_2 _10341_ (.Y(_05433_),
    .A(\soc_inst.core_mem_addr[27] ));
 sg13g2_inv_2 _10342_ (.Y(_05434_),
    .A(net1878));
 sg13g2_inv_1 _10343_ (.Y(_05435_),
    .A(net2173));
 sg13g2_inv_2 _10344_ (.Y(_05436_),
    .A(net2533));
 sg13g2_inv_2 _10345_ (.Y(_05437_),
    .A(\soc_inst.core_instr_addr[2] ));
 sg13g2_inv_2 _10346_ (.Y(_05438_),
    .A(\soc_inst.core_instr_addr[3] ));
 sg13g2_inv_1 _10347_ (.Y(_05439_),
    .A(\soc_inst.mem_ctrl.spi_addr[4] ));
 sg13g2_inv_2 _10348_ (.Y(_05440_),
    .A(\soc_inst.core_instr_addr[4] ));
 sg13g2_inv_2 _10349_ (.Y(_05441_),
    .A(\soc_inst.mem_ctrl.spi_addr[5] ));
 sg13g2_inv_1 _10350_ (.Y(_05442_),
    .A(net2629));
 sg13g2_inv_1 _10351_ (.Y(_05443_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ));
 sg13g2_inv_2 _10352_ (.Y(_05444_),
    .A(net2782));
 sg13g2_inv_2 _10353_ (.Y(_05445_),
    .A(net2737));
 sg13g2_inv_4 _10354_ (.A(net2707),
    .Y(_05446_));
 sg13g2_inv_1 _10355_ (.Y(_05447_),
    .A(\soc_inst.mem_ctrl.spi_addr[9] ));
 sg13g2_inv_4 _10356_ (.A(net2781),
    .Y(_05448_));
 sg13g2_inv_1 _10357_ (.Y(_05449_),
    .A(\soc_inst.mem_ctrl.spi_addr[10] ));
 sg13g2_inv_2 _10358_ (.Y(_05450_),
    .A(\soc_inst.core_instr_addr[10] ));
 sg13g2_inv_1 _10359_ (.Y(_05451_),
    .A(\soc_inst.mem_ctrl.spi_addr[11] ));
 sg13g2_inv_2 _10360_ (.Y(_05452_),
    .A(net2789));
 sg13g2_inv_2 _10361_ (.Y(_05453_),
    .A(net2931));
 sg13g2_inv_1 _10362_ (.Y(_05454_),
    .A(net2607));
 sg13g2_inv_2 _10363_ (.Y(_05455_),
    .A(\soc_inst.core_instr_addr[14] ));
 sg13g2_inv_2 _10364_ (.Y(_05456_),
    .A(net2832));
 sg13g2_inv_4 _10365_ (.A(net2853),
    .Y(_05457_));
 sg13g2_inv_4 _10366_ (.A(net2770),
    .Y(_05458_));
 sg13g2_inv_2 _10367_ (.Y(_05459_),
    .A(net2883));
 sg13g2_inv_2 _10368_ (.Y(_05460_),
    .A(net2855));
 sg13g2_inv_2 _10369_ (.Y(_05461_),
    .A(net2901));
 sg13g2_inv_2 _10370_ (.Y(_05462_),
    .A(net2909));
 sg13g2_inv_2 _10371_ (.Y(_05463_),
    .A(net1777));
 sg13g2_inv_4 _10372_ (.A(net2854),
    .Y(_05464_));
 sg13g2_inv_2 _10373_ (.Y(_05465_),
    .A(net2831));
 sg13g2_inv_1 _10374_ (.Y(_05466_),
    .A(net4779));
 sg13g2_inv_1 _10375_ (.Y(_05467_),
    .A(net4772));
 sg13g2_inv_1 _10376_ (.Y(_05468_),
    .A(\soc_inst.spi_inst.state[1] ));
 sg13g2_inv_2 _10377_ (.Y(_05469_),
    .A(net2566));
 sg13g2_inv_1 _10378_ (.Y(_05470_),
    .A(\soc_inst.mem_ctrl.spi_done ));
 sg13g2_inv_2 _10379_ (.Y(_05471_),
    .A(net2662));
 sg13g2_inv_1 _10380_ (.Y(_05472_),
    .A(net13));
 sg13g2_inv_1 _10381_ (.Y(_05473_),
    .A(net5128));
 sg13g2_inv_4 _10382_ (.A(net5054),
    .Y(_05474_));
 sg13g2_inv_2 _10383_ (.Y(_05475_),
    .A(net2014));
 sg13g2_inv_1 _10384_ (.Y(_05476_),
    .A(net1687));
 sg13g2_inv_1 _10385_ (.Y(_05477_),
    .A(net2804));
 sg13g2_inv_1 _10386_ (.Y(_05478_),
    .A(net2845));
 sg13g2_inv_1 _10387_ (.Y(_05479_),
    .A(net2786));
 sg13g2_inv_4 _10388_ (.A(net4884),
    .Y(_05480_));
 sg13g2_inv_2 _10389_ (.Y(_05481_),
    .A(\soc_inst.cpu_core.mem_reg_we ));
 sg13g2_inv_1 _10390_ (.Y(_05482_),
    .A(net2827));
 sg13g2_inv_1 _10391_ (.Y(_05483_),
    .A(net2760));
 sg13g2_inv_4 _10392_ (.A(net4799),
    .Y(_05484_));
 sg13g2_inv_4 _10393_ (.A(net4796),
    .Y(_05485_));
 sg13g2_inv_1 _10394_ (.Y(_05486_),
    .A(net2017));
 sg13g2_inv_4 _10395_ (.A(\soc_inst.pwm_inst.channel_idx [0]),
    .Y(_05487_));
 sg13g2_inv_1 _10396_ (.Y(_05488_),
    .A(net1902));
 sg13g2_inv_1 _10397_ (.Y(_05489_),
    .A(net1798));
 sg13g2_inv_1 _10398_ (.Y(_05490_),
    .A(net4782));
 sg13g2_inv_2 _10399_ (.Y(_05491_),
    .A(net2899));
 sg13g2_inv_2 _10400_ (.Y(_05492_),
    .A(net2868));
 sg13g2_inv_1 _10401_ (.Y(_05493_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ));
 sg13g2_inv_1 _10402_ (.Y(_05494_),
    .A(net5059));
 sg13g2_inv_4 _10403_ (.A(net2159),
    .Y(_05495_));
 sg13g2_inv_1 _10404_ (.Y(_05496_),
    .A(net496));
 sg13g2_inv_1 _10405_ (.Y(_05497_),
    .A(net2944));
 sg13g2_inv_1 _10406_ (.Y(_05498_),
    .A(net474));
 sg13g2_inv_1 _10407_ (.Y(_05499_),
    .A(net582));
 sg13g2_inv_1 _10408_ (.Y(_05500_),
    .A(net1034));
 sg13g2_inv_8 _10409_ (.Y(_05501_),
    .A(net5080));
 sg13g2_inv_1 _10410_ (.Y(_05502_),
    .A(\soc_inst.spi_inst.clock_divider[7] ));
 sg13g2_inv_1 _10411_ (.Y(_05503_),
    .A(net1120));
 sg13g2_inv_1 _10412_ (.Y(_05504_),
    .A(net397));
 sg13g2_inv_1 _10413_ (.Y(_05505_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ));
 sg13g2_inv_2 _10414_ (.Y(_05506_),
    .A(net2578));
 sg13g2_inv_1 _10415_ (.Y(_05507_),
    .A(\soc_inst.cpu_core.csr_file.mtime[3] ));
 sg13g2_inv_1 _10416_ (.Y(_05508_),
    .A(\soc_inst.cpu_core.csr_file.mtime[2] ));
 sg13g2_inv_1 _10417_ (.Y(_05509_),
    .A(\soc_inst.cpu_core.csr_file.mtime[7] ));
 sg13g2_inv_1 _10418_ (.Y(_05510_),
    .A(\soc_inst.cpu_core.csr_file.mtime[10] ));
 sg13g2_inv_1 _10419_ (.Y(_05511_),
    .A(\soc_inst.cpu_core.csr_file.mtime[9] ));
 sg13g2_inv_2 _10420_ (.Y(_05512_),
    .A(net2692));
 sg13g2_inv_1 _10421_ (.Y(_05513_),
    .A(net1772));
 sg13g2_inv_1 _10422_ (.Y(_05514_),
    .A(net1932));
 sg13g2_inv_1 _10423_ (.Y(_05515_),
    .A(net2587));
 sg13g2_inv_1 _10424_ (.Y(_05516_),
    .A(net2769));
 sg13g2_inv_1 _10425_ (.Y(_05517_),
    .A(\soc_inst.cpu_core.id_instr[2] ));
 sg13g2_inv_2 _10426_ (.Y(_05518_),
    .A(net2864));
 sg13g2_inv_1 _10427_ (.Y(_05519_),
    .A(net2135));
 sg13g2_inv_1 _10428_ (.Y(_05520_),
    .A(net2200));
 sg13g2_inv_1 _10429_ (.Y(_05521_),
    .A(net2034));
 sg13g2_inv_2 _10430_ (.Y(_05522_),
    .A(net978));
 sg13g2_inv_1 _10431_ (.Y(_05523_),
    .A(net2402));
 sg13g2_inv_1 _10432_ (.Y(_05524_),
    .A(net2287));
 sg13g2_inv_1 _10433_ (.Y(_05525_),
    .A(net2315));
 sg13g2_inv_1 _10434_ (.Y(_05526_),
    .A(net2229));
 sg13g2_inv_1 _10435_ (.Y(_05527_),
    .A(net2030));
 sg13g2_inv_1 _10436_ (.Y(_05528_),
    .A(net2285));
 sg13g2_inv_1 _10437_ (.Y(_05529_),
    .A(net2032));
 sg13g2_inv_1 _10438_ (.Y(_05530_),
    .A(net1898));
 sg13g2_inv_1 _10439_ (.Y(_05531_),
    .A(net1988));
 sg13g2_inv_1 _10440_ (.Y(_05532_),
    .A(net1816));
 sg13g2_inv_1 _10441_ (.Y(_05533_),
    .A(net1975));
 sg13g2_inv_1 _10442_ (.Y(_05534_),
    .A(net1946));
 sg13g2_inv_1 _10443_ (.Y(_05535_),
    .A(net1721));
 sg13g2_inv_1 _10444_ (.Y(_05536_),
    .A(net2368));
 sg13g2_inv_1 _10445_ (.Y(_05537_),
    .A(net2343));
 sg13g2_inv_1 _10446_ (.Y(_05538_),
    .A(net2026));
 sg13g2_inv_1 _10447_ (.Y(_05539_),
    .A(net1871));
 sg13g2_inv_1 _10448_ (.Y(_05540_),
    .A(net1741));
 sg13g2_inv_1 _10449_ (.Y(_05541_),
    .A(net2006));
 sg13g2_inv_1 _10450_ (.Y(_05542_),
    .A(net2164));
 sg13g2_inv_1 _10451_ (.Y(_05543_),
    .A(net616));
 sg13g2_inv_1 _10452_ (.Y(_05544_),
    .A(\soc_inst.spi_inst.rx_shift_reg[8] ));
 sg13g2_inv_1 _10453_ (.Y(_05545_),
    .A(\soc_inst.spi_inst.rx_shift_reg[24] ));
 sg13g2_inv_1 _10454_ (.Y(_05546_),
    .A(\soc_inst.spi_inst.rx_shift_reg[26] ));
 sg13g2_inv_1 _10455_ (.Y(_05547_),
    .A(\soc_inst.spi_inst.rx_shift_reg[27] ));
 sg13g2_inv_1 _10456_ (.Y(_05548_),
    .A(\soc_inst.spi_inst.rx_shift_reg[28] ));
 sg13g2_inv_1 _10457_ (.Y(_05549_),
    .A(\soc_inst.spi_inst.rx_shift_reg[29] ));
 sg13g2_inv_1 _10458_ (.Y(_05550_),
    .A(\soc_inst.spi_inst.rx_shift_reg[30] ));
 sg13g2_inv_1 _10459_ (.Y(_05551_),
    .A(net323));
 sg13g2_inv_1 _10460_ (.Y(_05552_),
    .A(net559));
 sg13g2_inv_1 _10461_ (.Y(_05553_),
    .A(net325));
 sg13g2_inv_1 _10462_ (.Y(_05554_),
    .A(net301));
 sg13g2_inv_1 _10463_ (.Y(_05555_),
    .A(net442));
 sg13g2_inv_1 _10464_ (.Y(_05556_),
    .A(net385));
 sg13g2_inv_1 _10465_ (.Y(_05557_),
    .A(net393));
 sg13g2_inv_1 _10466_ (.Y(_05558_),
    .A(net420));
 sg13g2_inv_1 _10467_ (.Y(_05559_),
    .A(net329));
 sg13g2_inv_1 _10468_ (.Y(_05560_),
    .A(net307));
 sg13g2_inv_1 _10469_ (.Y(_05561_),
    .A(net341));
 sg13g2_inv_1 _10470_ (.Y(_05562_),
    .A(net379));
 sg13g2_inv_1 _10471_ (.Y(_05563_),
    .A(net482));
 sg13g2_inv_1 _10472_ (.Y(_05564_),
    .A(net339));
 sg13g2_inv_1 _10473_ (.Y(_05565_),
    .A(net348));
 sg13g2_inv_1 _10474_ (.Y(_05566_),
    .A(net366));
 sg13g2_inv_1 _10475_ (.Y(_05567_),
    .A(\soc_inst.spi_inst.bit_counter[3] ));
 sg13g2_inv_1 _10476_ (.Y(_05568_),
    .A(net1122));
 sg13g2_inv_1 _10477_ (.Y(_05569_),
    .A(\soc_inst.pwm_inst.channel_counter[1][12] ));
 sg13g2_inv_1 _10478_ (.Y(_05570_),
    .A(\soc_inst.pwm_inst.channel_counter[1][11] ));
 sg13g2_inv_1 _10479_ (.Y(_05571_),
    .A(\soc_inst.pwm_inst.channel_counter[1][8] ));
 sg13g2_inv_1 _10480_ (.Y(_05572_),
    .A(\soc_inst.pwm_inst.channel_counter[1][3] ));
 sg13g2_inv_1 _10481_ (.Y(_05573_),
    .A(net910));
 sg13g2_inv_1 _10482_ (.Y(_05574_),
    .A(\soc_inst.pwm_inst.channel_counter[1][1] ));
 sg13g2_inv_1 _10483_ (.Y(_05575_),
    .A(net148));
 sg13g2_inv_1 _10484_ (.Y(_05576_),
    .A(\soc_inst.pwm_inst.channel_counter[0][10] ));
 sg13g2_inv_1 _10485_ (.Y(_05577_),
    .A(net5127));
 sg13g2_inv_1 _10486_ (.Y(_05578_),
    .A(\soc_inst.pwm_inst.channel_counter[0][8] ));
 sg13g2_inv_1 _10487_ (.Y(_05579_),
    .A(\soc_inst.pwm_inst.channel_counter[0][6] ));
 sg13g2_inv_1 _10488_ (.Y(_05580_),
    .A(\soc_inst.pwm_inst.channel_counter[0][5] ));
 sg13g2_inv_1 _10489_ (.Y(_05581_),
    .A(\soc_inst.pwm_inst.channel_counter[0][1] ));
 sg13g2_inv_1 _10490_ (.Y(_05582_),
    .A(\soc_inst.pwm_inst.channel_counter[0][0] ));
 sg13g2_inv_4 _10491_ (.A(net2072),
    .Y(_05583_));
 sg13g2_inv_4 _10492_ (.A(net2097),
    .Y(_05584_));
 sg13g2_inv_2 _10493_ (.Y(_05585_),
    .A(\soc_inst.mem_ctrl.spi_data_out[1] ));
 sg13g2_inv_2 _10494_ (.Y(_05586_),
    .A(\soc_inst.mem_ctrl.spi_data_out[3] ));
 sg13g2_inv_2 _10495_ (.Y(_05587_),
    .A(\soc_inst.mem_ctrl.spi_data_out[5] ));
 sg13g2_inv_1 _10496_ (.Y(_05588_),
    .A(\soc_inst.gpio_inst.gpio_out[0] ));
 sg13g2_inv_1 _10497_ (.Y(_05589_),
    .A(\soc_inst.pwm_inst.channel_duty[0][1] ));
 sg13g2_inv_1 _10498_ (.Y(_05590_),
    .A(\soc_inst.pwm_inst.channel_duty[1][1] ));
 sg13g2_inv_1 _10499_ (.Y(_05591_),
    .A(\soc_inst.spi_inst.done ));
 sg13g2_inv_1 _10500_ (.Y(_05592_),
    .A(\soc_inst.pwm_inst.channel_duty[0][2] ));
 sg13g2_inv_1 _10501_ (.Y(_05593_),
    .A(\soc_inst.pwm_inst.channel_duty[1][2] ));
 sg13g2_inv_1 _10502_ (.Y(_05594_),
    .A(\soc_inst.gpio_inst.gpio_out[3] ));
 sg13g2_inv_1 _10503_ (.Y(_05595_),
    .A(\soc_inst.pwm_inst.channel_duty[1][4] ));
 sg13g2_inv_2 _10504_ (.Y(_05596_),
    .A(\soc_inst.gpio_inst.gpio_out[4] ));
 sg13g2_inv_1 _10505_ (.Y(_05597_),
    .A(\soc_inst.pwm_inst.channel_duty[1][5] ));
 sg13g2_inv_2 _10506_ (.Y(_05598_),
    .A(\soc_inst.gpio_inst.gpio_out[5] ));
 sg13g2_inv_1 _10507_ (.Y(_05599_),
    .A(\soc_inst.pwm_inst.channel_duty[0][6] ));
 sg13g2_inv_1 _10508_ (.Y(_05600_),
    .A(\soc_inst.pwm_inst.channel_duty[1][6] ));
 sg13g2_inv_1 _10509_ (.Y(_05601_),
    .A(\soc_inst.pwm_inst.channel_duty[0][7] ));
 sg13g2_inv_1 _10510_ (.Y(_05602_),
    .A(\soc_inst.pwm_inst.channel_duty[1][7] ));
 sg13g2_inv_1 _10511_ (.Y(_05603_),
    .A(\soc_inst.spi_inst.rx_shift_reg[31] ));
 sg13g2_inv_1 _10512_ (.Y(_05604_),
    .A(\soc_inst.pwm_inst.channel_duty[0][8] ));
 sg13g2_inv_1 _10513_ (.Y(_05605_),
    .A(\soc_inst.pwm_inst.channel_duty[0][9] ));
 sg13g2_inv_1 _10514_ (.Y(_05606_),
    .A(\soc_inst.pwm_inst.channel_duty[1][10] ));
 sg13g2_inv_1 _10515_ (.Y(_05607_),
    .A(\soc_inst.pwm_inst.channel_duty[0][11] ));
 sg13g2_inv_1 _10516_ (.Y(_05608_),
    .A(\soc_inst.pwm_inst.channel_duty[1][11] ));
 sg13g2_inv_1 _10517_ (.Y(_05609_),
    .A(\soc_inst.pwm_inst.channel_duty[0][12] ));
 sg13g2_inv_1 _10518_ (.Y(_05610_),
    .A(\soc_inst.pwm_inst.channel_duty[0][13] ));
 sg13g2_inv_1 _10519_ (.Y(_05611_),
    .A(net1623));
 sg13g2_inv_1 _10520_ (.Y(_05612_),
    .A(net2843));
 sg13g2_inv_1 _10521_ (.Y(_05613_),
    .A(net752));
 sg13g2_inv_1 _10522_ (.Y(_05614_),
    .A(net2721));
 sg13g2_inv_1 _10523_ (.Y(_05615_),
    .A(net2902));
 sg13g2_inv_1 _10524_ (.Y(_05616_),
    .A(net1435));
 sg13g2_inv_1 _10525_ (.Y(_05617_),
    .A(net837));
 sg13g2_inv_1 _10526_ (.Y(_05618_),
    .A(net2683));
 sg13g2_inv_1 _10527_ (.Y(_05619_),
    .A(net1016));
 sg13g2_inv_1 _10528_ (.Y(_05620_),
    .A(net999));
 sg13g2_inv_1 _10529_ (.Y(_05621_),
    .A(net1208));
 sg13g2_inv_1 _10530_ (.Y(_05622_),
    .A(net949));
 sg13g2_inv_1 _10531_ (.Y(_05623_),
    .A(net2484));
 sg13g2_inv_1 _10532_ (.Y(_05624_),
    .A(net2559));
 sg13g2_inv_2 _10533_ (.Y(_05625_),
    .A(net1072));
 sg13g2_inv_1 _10534_ (.Y(_05626_),
    .A(net789));
 sg13g2_inv_1 _10535_ (.Y(_05627_),
    .A(net1914));
 sg13g2_inv_1 _10536_ (.Y(_05628_),
    .A(net538));
 sg13g2_inv_1 _10537_ (.Y(_05629_),
    .A(net832));
 sg13g2_inv_1 _10538_ (.Y(_05630_),
    .A(net930));
 sg13g2_inv_1 _10539_ (.Y(_05631_),
    .A(net2061));
 sg13g2_inv_2 _10540_ (.Y(_05632_),
    .A(net618));
 sg13g2_inv_1 _10541_ (.Y(_05633_),
    .A(net2115));
 sg13g2_inv_2 _10542_ (.Y(_05634_),
    .A(net733));
 sg13g2_inv_1 _10543_ (.Y(_05635_),
    .A(net1104));
 sg13g2_inv_1 _10544_ (.Y(_05636_),
    .A(net1197));
 sg13g2_inv_1 _10545_ (.Y(_05637_),
    .A(net1307));
 sg13g2_inv_2 _10546_ (.Y(_05638_),
    .A(net631));
 sg13g2_inv_1 _10547_ (.Y(_05639_),
    .A(net1634));
 sg13g2_inv_1 _10548_ (.Y(_05640_),
    .A(net1578));
 sg13g2_inv_1 _10549_ (.Y(_05641_),
    .A(net1713));
 sg13g2_inv_1 _10550_ (.Y(_05642_),
    .A(net1886));
 sg13g2_inv_1 _10551_ (.Y(_05643_),
    .A(net925));
 sg13g2_inv_1 _10552_ (.Y(_05644_),
    .A(net1408));
 sg13g2_inv_1 _10553_ (.Y(_05645_),
    .A(net1949));
 sg13g2_inv_1 _10554_ (.Y(_05646_),
    .A(net1199));
 sg13g2_inv_1 _10555_ (.Y(_05647_),
    .A(net472));
 sg13g2_inv_2 _10556_ (.Y(_05648_),
    .A(net5082));
 sg13g2_inv_4 _10557_ (.A(net5095),
    .Y(_05649_));
 sg13g2_inv_2 _10558_ (.Y(_05650_),
    .A(net5091));
 sg13g2_inv_2 _10559_ (.Y(_05651_),
    .A(\soc_inst.cpu_core.id_rs2_data[0] ));
 sg13g2_inv_2 _10560_ (.Y(_05652_),
    .A(\soc_inst.cpu_core.id_rs1_data[7] ));
 sg13g2_inv_2 _10561_ (.Y(_05653_),
    .A(\soc_inst.cpu_core.id_rs1_data[6] ));
 sg13g2_inv_2 _10562_ (.Y(_05654_),
    .A(\soc_inst.cpu_core.id_rs1_data[5] ));
 sg13g2_inv_2 _10563_ (.Y(_05655_),
    .A(\soc_inst.cpu_core.id_rs2_data[5] ));
 sg13g2_inv_2 _10564_ (.Y(_05656_),
    .A(\soc_inst.cpu_core.id_rs1_data[4] ));
 sg13g2_inv_2 _10565_ (.Y(_05657_),
    .A(\soc_inst.cpu_core.id_rs2_data[4] ));
 sg13g2_inv_2 _10566_ (.Y(_05658_),
    .A(\soc_inst.cpu_core.id_rs1_data[15] ));
 sg13g2_inv_4 _10567_ (.A(\soc_inst.cpu_core.id_rs2_data[15] ),
    .Y(_05659_));
 sg13g2_inv_1 _10568_ (.Y(_05660_),
    .A(\soc_inst.cpu_core.id_rs1_data[14] ));
 sg13g2_inv_4 _10569_ (.A(\soc_inst.cpu_core.id_rs2_data[10] ),
    .Y(_05661_));
 sg13g2_inv_4 _10570_ (.A(\soc_inst.cpu_core.id_rs2_data[8] ),
    .Y(_05662_));
 sg13g2_inv_2 _10571_ (.Y(_05663_),
    .A(\soc_inst.cpu_core.id_rs1_data[30] ));
 sg13g2_inv_4 _10572_ (.A(\soc_inst.cpu_core.id_rs2_data[28] ),
    .Y(_05664_));
 sg13g2_inv_4 _10573_ (.A(\soc_inst.cpu_core.id_rs2_data[27] ),
    .Y(_05665_));
 sg13g2_inv_2 _10574_ (.Y(_05666_),
    .A(\soc_inst.cpu_core.id_rs1_data[26] ));
 sg13g2_inv_4 _10575_ (.A(\soc_inst.cpu_core.id_rs2_data[24] ),
    .Y(_05667_));
 sg13g2_inv_2 _10576_ (.Y(_05668_),
    .A(\soc_inst.cpu_core.id_rs1_data[23] ));
 sg13g2_inv_2 _10577_ (.Y(_05669_),
    .A(\soc_inst.cpu_core.id_rs2_data[23] ));
 sg13g2_inv_1 _10578_ (.Y(_05670_),
    .A(\soc_inst.cpu_core.id_rs1_data[22] ));
 sg13g2_inv_4 _10579_ (.A(net2235),
    .Y(_05671_));
 sg13g2_inv_2 _10580_ (.Y(_05672_),
    .A(\soc_inst.cpu_core.id_rs1_data[21] ));
 sg13g2_inv_2 _10581_ (.Y(_05673_),
    .A(net1648));
 sg13g2_inv_1 _10582_ (.Y(_05674_),
    .A(\soc_inst.cpu_core.id_rs1_data[19] ));
 sg13g2_inv_8 _10583_ (.Y(_05675_),
    .A(\soc_inst.cpu_core.id_rs2_data[19] ));
 sg13g2_inv_2 _10584_ (.Y(_05676_),
    .A(\soc_inst.cpu_core.id_rs1_data[18] ));
 sg13g2_inv_1 _10585_ (.Y(_05677_),
    .A(\soc_inst.cpu_core.id_pc[0] ));
 sg13g2_inv_1 _10586_ (.Y(_05678_),
    .A(\soc_inst.cpu_core.id_pc[1] ));
 sg13g2_inv_1 _10587_ (.Y(_05679_),
    .A(\soc_inst.cpu_core.id_pc[2] ));
 sg13g2_inv_1 _10588_ (.Y(_05680_),
    .A(\soc_inst.cpu_core.id_pc[3] ));
 sg13g2_inv_2 _10589_ (.Y(_05681_),
    .A(net2582));
 sg13g2_inv_2 _10590_ (.Y(_05682_),
    .A(\soc_inst.cpu_core.id_pc[5] ));
 sg13g2_inv_2 _10591_ (.Y(_05683_),
    .A(\soc_inst.cpu_core.id_pc[6] ));
 sg13g2_inv_1 _10592_ (.Y(_05684_),
    .A(\soc_inst.cpu_core.id_pc[7] ));
 sg13g2_inv_1 _10593_ (.Y(_05685_),
    .A(\soc_inst.cpu_core.id_pc[8] ));
 sg13g2_inv_1 _10594_ (.Y(_05686_),
    .A(\soc_inst.cpu_core.id_pc[9] ));
 sg13g2_inv_2 _10595_ (.Y(_05687_),
    .A(\soc_inst.cpu_core.id_pc[10] ));
 sg13g2_inv_1 _10596_ (.Y(_05688_),
    .A(\soc_inst.cpu_core.id_imm[10] ));
 sg13g2_inv_2 _10597_ (.Y(_05689_),
    .A(\soc_inst.cpu_core.id_pc[11] ));
 sg13g2_inv_1 _10598_ (.Y(_05690_),
    .A(\soc_inst.cpu_core.id_imm[11] ));
 sg13g2_inv_2 _10599_ (.Y(_05691_),
    .A(\soc_inst.cpu_core.id_pc[12] ));
 sg13g2_inv_1 _10600_ (.Y(_05692_),
    .A(\soc_inst.cpu_core.id_pc[13] ));
 sg13g2_inv_4 _10601_ (.A(\soc_inst.cpu_core.id_pc[14] ),
    .Y(_05693_));
 sg13g2_inv_2 _10602_ (.Y(_05694_),
    .A(\soc_inst.cpu_core.id_pc[15] ));
 sg13g2_inv_1 _10603_ (.Y(_05695_),
    .A(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_inv_1 _10604_ (.Y(_05696_),
    .A(\soc_inst.cpu_core.id_pc[16] ));
 sg13g2_inv_2 _10605_ (.Y(_05697_),
    .A(\soc_inst.cpu_core.id_pc[17] ));
 sg13g2_inv_2 _10606_ (.Y(_05698_),
    .A(\soc_inst.cpu_core.id_pc[18] ));
 sg13g2_inv_2 _10607_ (.Y(_05699_),
    .A(net2985));
 sg13g2_inv_2 _10608_ (.Y(_05700_),
    .A(\soc_inst.cpu_core.id_pc[20] ));
 sg13g2_inv_1 _10609_ (.Y(_05701_),
    .A(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_inv_2 _10610_ (.Y(_05702_),
    .A(\soc_inst.cpu_core.id_pc[21] ));
 sg13g2_inv_1 _10611_ (.Y(_05703_),
    .A(\soc_inst.cpu_core.id_pc[22] ));
 sg13g2_inv_4 _10612_ (.A(\soc_inst.cpu_core.id_pc[23] ),
    .Y(_05704_));
 sg13g2_inv_1 _10613_ (.Y(_05705_),
    .A(\soc_inst.cpu_core.id_imm[23] ));
 sg13g2_inv_1 _10614_ (.Y(_05706_),
    .A(\soc_inst.cpu_core.id_imm[30] ));
 sg13g2_inv_2 _10615_ (.Y(_05707_),
    .A(net1888));
 sg13g2_inv_1 _10616_ (.Y(_05708_),
    .A(net2384));
 sg13g2_inv_2 _10617_ (.Y(_05709_),
    .A(net630));
 sg13g2_inv_1 _10618_ (.Y(_05710_),
    .A(net1037));
 sg13g2_inv_1 _10619_ (.Y(_05711_),
    .A(net2516));
 sg13g2_inv_1 _10620_ (.Y(_05712_),
    .A(net2746));
 sg13g2_inv_1 _10621_ (.Y(_05713_),
    .A(net2520));
 sg13g2_inv_1 _10622_ (.Y(_05714_),
    .A(net2062));
 sg13g2_inv_1 _10623_ (.Y(_05715_),
    .A(net2225));
 sg13g2_inv_2 _10624_ (.Y(_05716_),
    .A(net2350));
 sg13g2_inv_1 _10625_ (.Y(_05717_),
    .A(net2768));
 sg13g2_inv_1 _10626_ (.Y(_05718_),
    .A(net1069));
 sg13g2_inv_1 _10627_ (.Y(_05719_),
    .A(net675));
 sg13g2_inv_1 _10628_ (.Y(_05720_),
    .A(net526));
 sg13g2_inv_1 _10629_ (.Y(_05721_),
    .A(\soc_inst.cpu_core.if_instr[5] ));
 sg13g2_inv_1 _10630_ (.Y(_05722_),
    .A(net905));
 sg13g2_inv_1 _10631_ (.Y(_05723_),
    .A(net512));
 sg13g2_inv_1 _10632_ (.Y(_05724_),
    .A(net548));
 sg13g2_inv_1 _10633_ (.Y(_05725_),
    .A(net1986));
 sg13g2_inv_1 _10634_ (.Y(_05726_),
    .A(\soc_inst.cpu_core.register_file.registers[1][14] ));
 sg13g2_inv_1 _10635_ (.Y(_05727_),
    .A(\soc_inst.cpu_core.register_file.registers[1][15] ));
 sg13g2_inv_1 _10636_ (.Y(_05728_),
    .A(\soc_inst.cpu_core.register_file.registers[1][17] ));
 sg13g2_inv_1 _10637_ (.Y(_05729_),
    .A(net561));
 sg13g2_inv_1 _10638_ (.Y(_05730_),
    .A(\soc_inst.cpu_core.register_file.registers[1][24] ));
 sg13g2_inv_1 _10639_ (.Y(_05731_),
    .A(net1268));
 sg13g2_inv_1 _10640_ (.Y(_05732_),
    .A(net454));
 sg13g2_inv_1 _10641_ (.Y(_05733_),
    .A(net528));
 sg13g2_inv_1 _10642_ (.Y(_05734_),
    .A(net1296));
 sg13g2_inv_1 _10643_ (.Y(_05735_),
    .A(net2185));
 sg13g2_inv_1 _10644_ (.Y(_05736_),
    .A(net1070));
 sg13g2_inv_1 _10645_ (.Y(_05737_),
    .A(net2245));
 sg13g2_inv_1 _10646_ (.Y(_05738_),
    .A(net1350));
 sg13g2_inv_1 _10647_ (.Y(_05739_),
    .A(net1748));
 sg13g2_inv_1 _10648_ (.Y(_05740_),
    .A(net1737));
 sg13g2_inv_1 _10649_ (.Y(_05741_),
    .A(net943));
 sg13g2_inv_1 _10650_ (.Y(_05742_),
    .A(net1206));
 sg13g2_inv_1 _10651_ (.Y(_05743_),
    .A(net859));
 sg13g2_inv_1 _10652_ (.Y(_05744_),
    .A(net2051));
 sg13g2_inv_1 _10653_ (.Y(_05745_),
    .A(net918));
 sg13g2_inv_1 _10654_ (.Y(_05746_),
    .A(net1195));
 sg13g2_inv_1 _10655_ (.Y(_05747_),
    .A(net887));
 sg13g2_inv_1 _10656_ (.Y(_05748_),
    .A(net1166));
 sg13g2_inv_1 _10657_ (.Y(_05749_),
    .A(net1161));
 sg13g2_inv_1 _10658_ (.Y(_05750_),
    .A(net1957));
 sg13g2_inv_1 _10659_ (.Y(_05751_),
    .A(net1658));
 sg13g2_inv_1 _10660_ (.Y(_05752_),
    .A(net1246));
 sg13g2_inv_1 _10661_ (.Y(_05753_),
    .A(net1419));
 sg13g2_inv_1 _10662_ (.Y(_05754_),
    .A(net1509));
 sg13g2_inv_1 _10663_ (.Y(_05755_),
    .A(net1569));
 sg13g2_inv_1 _10664_ (.Y(_05756_),
    .A(net1646));
 sg13g2_inv_1 _10665_ (.Y(_05757_),
    .A(net1439));
 sg13g2_inv_1 _10666_ (.Y(_05758_),
    .A(net2751));
 sg13g2_inv_1 _10667_ (.Y(_05759_),
    .A(net2777));
 sg13g2_inv_1 _10668_ (.Y(_05760_),
    .A(net2743));
 sg13g2_inv_1 _10669_ (.Y(_05761_),
    .A(net2923));
 sg13g2_inv_1 _10670_ (.Y(_05762_),
    .A(net2908));
 sg13g2_inv_4 _10671_ (.A(net2105),
    .Y(_05763_));
 sg13g2_inv_1 _10672_ (.Y(_05764_),
    .A(net2867));
 sg13g2_inv_1 _10673_ (.Y(_05765_),
    .A(net2817));
 sg13g2_inv_1 _10674_ (.Y(_05766_),
    .A(net2802));
 sg13g2_inv_1 _10675_ (.Y(_05767_),
    .A(net2426));
 sg13g2_inv_1 _10676_ (.Y(_05768_),
    .A(net2773));
 sg13g2_inv_1 _10677_ (.Y(_05769_),
    .A(net2833));
 sg13g2_inv_1 _10678_ (.Y(_05770_),
    .A(net2649));
 sg13g2_inv_1 _10679_ (.Y(_05771_),
    .A(net2815));
 sg13g2_inv_1 _10680_ (.Y(_05772_),
    .A(net2673));
 sg13g2_inv_1 _10681_ (.Y(_05773_),
    .A(net1784));
 sg13g2_inv_2 _10682_ (.Y(_05774_),
    .A(net1157));
 sg13g2_inv_2 _10683_ (.Y(_05775_),
    .A(net742));
 sg13g2_inv_1 _10684_ (.Y(_05776_),
    .A(net1391));
 sg13g2_inv_1 _10685_ (.Y(_05777_),
    .A(net1876));
 sg13g2_inv_2 _10686_ (.Y(_05778_),
    .A(net424));
 sg13g2_inv_2 _10687_ (.Y(_05779_),
    .A(net1228));
 sg13g2_inv_1 _10688_ (.Y(_05780_),
    .A(net1821));
 sg13g2_inv_2 _10689_ (.Y(_05781_),
    .A(net448));
 sg13g2_inv_1 _10690_ (.Y(_05782_),
    .A(net1459));
 sg13g2_inv_1 _10691_ (.Y(_05783_),
    .A(net1530));
 sg13g2_inv_1 _10692_ (.Y(_05784_),
    .A(\soc_inst.spi_inst.spi_mosi ));
 sg13g2_inv_1 _10693_ (.Y(_05785_),
    .A(net2283));
 sg13g2_inv_1 _10694_ (.Y(_05786_),
    .A(net1694));
 sg13g2_inv_1 _10695_ (.Y(_05787_),
    .A(net2911));
 sg13g2_inv_1 _10696_ (.Y(_05788_),
    .A(net2429));
 sg13g2_inv_1 _10697_ (.Y(_05789_),
    .A(net1602));
 sg13g2_inv_1 _10698_ (.Y(_05790_),
    .A(net2718));
 sg13g2_inv_1 _10699_ (.Y(_05791_),
    .A(net2028));
 sg13g2_inv_1 _10700_ (.Y(_05792_),
    .A(net1858));
 sg13g2_inv_1 _10701_ (.Y(_05793_),
    .A(net2470));
 sg13g2_inv_1 _10702_ (.Y(_05794_),
    .A(net1130));
 sg13g2_inv_1 _10703_ (.Y(_05795_),
    .A(net2389));
 sg13g2_inv_2 _10704_ (.Y(_05796_),
    .A(net2826));
 sg13g2_inv_1 _10705_ (.Y(_05797_),
    .A(net2591));
 sg13g2_inv_1 _10706_ (.Y(_05798_),
    .A(net2688));
 sg13g2_inv_1 _10707_ (.Y(_05799_),
    .A(net2627));
 sg13g2_inv_1 _10708_ (.Y(_05800_),
    .A(net4860));
 sg13g2_inv_1 _10709_ (.Y(_05801_),
    .A(net2617));
 sg13g2_inv_1 _10710_ (.Y(_05802_),
    .A(net4861));
 sg13g2_inv_1 _10711_ (.Y(_05803_),
    .A(net2480));
 sg13g2_inv_1 _10712_ (.Y(_05804_),
    .A(net4862));
 sg13g2_inv_2 _10713_ (.Y(_05805_),
    .A(net1317));
 sg13g2_inv_4 _10714_ (.A(net2711),
    .Y(_05806_));
 sg13g2_inv_1 _10715_ (.Y(_05807_),
    .A(net1897));
 sg13g2_inv_1 _10716_ (.Y(_05808_),
    .A(net2601));
 sg13g2_inv_2 _10717_ (.Y(_05809_),
    .A(net2144));
 sg13g2_inv_4 _10718_ (.A(net2792),
    .Y(_05810_));
 sg13g2_inv_2 _10719_ (.Y(_05811_),
    .A(net854));
 sg13g2_inv_4 _10720_ (.A(net2465),
    .Y(_05812_));
 sg13g2_inv_1 _10721_ (.Y(_05813_),
    .A(net2621));
 sg13g2_inv_1 _10722_ (.Y(_05814_),
    .A(net4863));
 sg13g2_inv_1 _10723_ (.Y(_05815_),
    .A(net1895));
 sg13g2_inv_2 _10724_ (.Y(_05816_),
    .A(net2895));
 sg13g2_inv_1 _10725_ (.Y(_05817_),
    .A(net1415));
 sg13g2_inv_1 _10726_ (.Y(_05818_),
    .A(net2519));
 sg13g2_inv_1 _10727_ (.Y(_05819_),
    .A(net1960));
 sg13g2_inv_2 _10728_ (.Y(_05820_),
    .A(net2719));
 sg13g2_inv_1 _10729_ (.Y(_05821_),
    .A(net1495));
 sg13g2_inv_2 _10730_ (.Y(_05822_),
    .A(net2417));
 sg13g2_inv_1 _10731_ (.Y(_05823_),
    .A(net2474));
 sg13g2_inv_2 _10732_ (.Y(_05824_),
    .A(net2380));
 sg13g2_inv_1 _10733_ (.Y(_05825_),
    .A(net1411));
 sg13g2_inv_1 _10734_ (.Y(_05826_),
    .A(net1688));
 sg13g2_inv_1 _10735_ (.Y(_05827_),
    .A(net1386));
 sg13g2_inv_2 _10736_ (.Y(_05828_),
    .A(net1922));
 sg13g2_inv_1 _10737_ (.Y(_05829_),
    .A(net1159));
 sg13g2_inv_2 _10738_ (.Y(_05830_),
    .A(net2333));
 sg13g2_inv_1 _10739_ (.Y(_05831_),
    .A(net4806));
 sg13g2_inv_4 _10740_ (.A(net2518),
    .Y(_05832_));
 sg13g2_inv_1 _10741_ (.Y(_05833_),
    .A(net4815));
 sg13g2_inv_1 _10742_ (.Y(_05834_),
    .A(net2455));
 sg13g2_inv_1 _10743_ (.Y(_05835_),
    .A(net4817));
 sg13g2_inv_1 _10744_ (.Y(_05836_),
    .A(net998));
 sg13g2_inv_1 _10745_ (.Y(_05837_),
    .A(net4838));
 sg13g2_inv_1 _10746_ (.Y(_05838_),
    .A(net2396));
 sg13g2_inv_4 _10747_ (.A(net4850),
    .Y(_05839_));
 sg13g2_inv_1 _10748_ (.Y(_05840_),
    .A(net2345));
 sg13g2_inv_1 _10749_ (.Y(_05841_),
    .A(net696));
 sg13g2_inv_1 _10750_ (.Y(_05842_),
    .A(net861));
 sg13g2_inv_1 _10751_ (.Y(_05843_),
    .A(net589));
 sg13g2_inv_1 _10752_ (.Y(_05844_),
    .A(net806));
 sg13g2_inv_1 _10753_ (.Y(_05845_),
    .A(net1395));
 sg13g2_inv_1 _10754_ (.Y(_05846_),
    .A(net1031));
 sg13g2_inv_1 _10755_ (.Y(_05847_),
    .A(net914));
 sg13g2_inv_1 _10756_ (.Y(_05848_),
    .A(net704));
 sg13g2_inv_1 _10757_ (.Y(_05849_),
    .A(net628));
 sg13g2_inv_1 _10758_ (.Y(_05850_),
    .A(net700));
 sg13g2_inv_1 _10759_ (.Y(_05851_),
    .A(net852));
 sg13g2_inv_1 _10760_ (.Y(_05852_),
    .A(net692));
 sg13g2_inv_1 _10761_ (.Y(_05853_),
    .A(net406));
 sg13g2_inv_1 _10762_ (.Y(_05854_),
    .A(net955));
 sg13g2_inv_1 _10763_ (.Y(_05855_),
    .A(net414));
 sg13g2_inv_1 _10764_ (.Y(_05856_),
    .A(net595));
 sg13g2_inv_1 _10765_ (.Y(_05857_),
    .A(net612));
 sg13g2_inv_1 _10766_ (.Y(_05858_),
    .A(net436));
 sg13g2_inv_1 _10767_ (.Y(_05859_),
    .A(net377));
 sg13g2_inv_1 _10768_ (.Y(_05860_),
    .A(net740));
 sg13g2_inv_1 _10769_ (.Y(_05861_),
    .A(net346));
 sg13g2_inv_1 _10770_ (.Y(_05862_),
    .A(net1678));
 sg13g2_inv_4 _10771_ (.A(net2599),
    .Y(_05863_));
 sg13g2_inv_1 _10772_ (.Y(_05864_),
    .A(net2404));
 sg13g2_inv_1 _10773_ (.Y(_05865_),
    .A(net5073));
 sg13g2_inv_1 _10774_ (.Y(_05866_),
    .A(net2808));
 sg13g2_nor2_1 _10775_ (.A(net599),
    .B(\soc_inst.core_mem_re ),
    .Y(_05867_));
 sg13g2_nor2_1 _10776_ (.A(\soc_inst.core_mem_we ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .Y(_05868_));
 sg13g2_and2_1 _10777_ (.A(_05867_),
    .B(_05868_),
    .X(_05869_));
 sg13g2_nand2_2 _10778_ (.Y(_05870_),
    .A(_05867_),
    .B(_05868_));
 sg13g2_and2_1 _10779_ (.A(net5074),
    .B(_05870_),
    .X(_05871_));
 sg13g2_nand2_2 _10780_ (.Y(_05872_),
    .A(net5074),
    .B(_05870_));
 sg13g2_nor4_2 _10781_ (.A(\soc_inst.core_mem_addr[21] ),
    .B(\soc_inst.core_mem_addr[20] ),
    .C(\soc_inst.core_mem_addr[23] ),
    .Y(_05873_),
    .D(\soc_inst.core_mem_addr[22] ));
 sg13g2_nor4_2 _10782_ (.A(\soc_inst.core_mem_addr[17] ),
    .B(\soc_inst.core_mem_addr[16] ),
    .C(\soc_inst.core_mem_addr[19] ),
    .Y(_05874_),
    .D(\soc_inst.core_mem_addr[18] ));
 sg13g2_nand2_2 _10783_ (.Y(_05875_),
    .A(_05873_),
    .B(_05874_));
 sg13g2_nand3_1 _10784_ (.B(_05873_),
    .C(_05874_),
    .A(\soc_inst.core_mem_addr[13] ),
    .Y(_05876_));
 sg13g2_nand4_1 _10785_ (.B(_05421_),
    .C(_05424_),
    .A(_05420_),
    .Y(_05877_),
    .D(\soc_inst.core_mem_addr[30] ));
 sg13g2_nor3_2 _10786_ (.A(\soc_inst.core_mem_addr[29] ),
    .B(\soc_inst.core_mem_addr[28] ),
    .C(\soc_inst.core_mem_addr[31] ),
    .Y(_05878_));
 sg13g2_nor4_2 _10787_ (.A(\soc_inst.core_mem_addr[25] ),
    .B(\soc_inst.core_mem_addr[24] ),
    .C(\soc_inst.core_mem_addr[27] ),
    .Y(_05879_),
    .D(\soc_inst.core_mem_addr[26] ));
 sg13g2_nand2_1 _10788_ (.Y(_05880_),
    .A(_05878_),
    .B(_05879_));
 sg13g2_nor4_2 _10789_ (.A(\soc_inst.core_mem_addr[8] ),
    .B(\soc_inst.core_mem_addr[9] ),
    .C(_05877_),
    .Y(_05881_),
    .D(_05880_));
 sg13g2_and2_1 _10790_ (.A(_05425_),
    .B(_05881_),
    .X(_05882_));
 sg13g2_nor2b_1 _10791_ (.A(_05876_),
    .B_N(_05882_),
    .Y(_05883_));
 sg13g2_nor2_1 _10792_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(_05875_),
    .Y(_05884_));
 sg13g2_and2_1 _10793_ (.A(_05881_),
    .B(_05884_),
    .X(_05885_));
 sg13g2_o21ai_1 _10794_ (.B1(_05870_),
    .Y(_05886_),
    .A1(_05883_),
    .A2(_05885_));
 sg13g2_nand2_2 _10795_ (.Y(_05887_),
    .A(\soc_inst.core_mem_addr[12] ),
    .B(_05884_));
 sg13g2_nor3_1 _10796_ (.A(\soc_inst.core_mem_addr[8] ),
    .B(\soc_inst.core_mem_addr[9] ),
    .C(\soc_inst.core_mem_addr[11] ),
    .Y(_05888_));
 sg13g2_nor2_1 _10797_ (.A(\soc_inst.core_mem_addr[10] ),
    .B(_05434_),
    .Y(_05889_));
 sg13g2_nand4_1 _10798_ (.B(_05879_),
    .C(_05888_),
    .A(_05878_),
    .Y(_05890_),
    .D(_05889_));
 sg13g2_nor3_1 _10799_ (.A(\soc_inst.core_mem_addr[15] ),
    .B(\soc_inst.core_mem_addr[14] ),
    .C(_05890_),
    .Y(_05891_));
 sg13g2_nor3_2 _10800_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(net4787),
    .C(_05875_),
    .Y(_05892_));
 sg13g2_and2_1 _10801_ (.A(\soc_inst.core_mem_addr[30] ),
    .B(_05879_),
    .X(_05893_));
 sg13g2_nand4_1 _10802_ (.B(_05878_),
    .C(_05888_),
    .A(_05421_),
    .Y(_05894_),
    .D(_05893_));
 sg13g2_nand3b_1 _10803_ (.B(_05425_),
    .C(_05424_),
    .Y(_05895_),
    .A_N(_05894_));
 sg13g2_nor2_2 _10804_ (.A(_05876_),
    .B(_05895_),
    .Y(_05896_));
 sg13g2_nor2_2 _10805_ (.A(_05887_),
    .B(_05895_),
    .Y(_05897_));
 sg13g2_nor3_1 _10806_ (.A(\soc_inst.core_mem_addr[15] ),
    .B(_05425_),
    .C(_05894_),
    .Y(_05898_));
 sg13g2_nor2b_2 _10807_ (.A(_05887_),
    .B_N(_05898_),
    .Y(_05899_));
 sg13g2_nor3_1 _10808_ (.A(\soc_inst.core_mem_addr[15] ),
    .B(_05887_),
    .C(_05894_),
    .Y(_05900_));
 sg13g2_nor4_2 _10809_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(net4787),
    .C(_05875_),
    .Y(_05901_),
    .D(_05895_));
 sg13g2_and2_1 _10810_ (.A(_05892_),
    .B(_05898_),
    .X(_05902_));
 sg13g2_nor4_1 _10811_ (.A(_05896_),
    .B(_05900_),
    .C(_05901_),
    .D(_05902_),
    .Y(_05903_));
 sg13g2_nor2_2 _10812_ (.A(_05869_),
    .B(_05903_),
    .Y(_05904_));
 sg13g2_or2_1 _10813_ (.X(_05905_),
    .B(_05903_),
    .A(_05869_));
 sg13g2_nor2_2 _10814_ (.A(_05871_),
    .B(net4015),
    .Y(_05906_));
 sg13g2_nand2_1 _10815_ (.Y(_05907_),
    .A(_05872_),
    .B(net4066));
 sg13g2_nor3_1 _10816_ (.A(net5074),
    .B(_05469_),
    .C(_05470_),
    .Y(_05908_));
 sg13g2_o21ai_1 _10817_ (.B1(_05906_),
    .Y(_05909_),
    .A1(net2748),
    .A2(_05908_));
 sg13g2_xor2_1 _10818_ (.B(\soc_inst.core_instr_addr[7] ),
    .A(\soc_inst.mem_ctrl.spi_addr[7] ),
    .X(_05910_));
 sg13g2_xor2_1 _10819_ (.B(\soc_inst.core_instr_addr[1] ),
    .A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .X(_05911_));
 sg13g2_xor2_1 _10820_ (.B(\soc_inst.core_instr_addr[16] ),
    .A(\soc_inst.mem_ctrl.spi_addr[16] ),
    .X(_05912_));
 sg13g2_xnor2_1 _10821_ (.Y(_05913_),
    .A(\soc_inst.mem_ctrl.spi_addr[14] ),
    .B(\soc_inst.core_instr_addr[14] ));
 sg13g2_xor2_1 _10822_ (.B(\soc_inst.core_instr_addr[15] ),
    .A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .X(_05914_));
 sg13g2_xor2_1 _10823_ (.B(\soc_inst.core_instr_addr[20] ),
    .A(\soc_inst.mem_ctrl.spi_addr[20] ),
    .X(_05915_));
 sg13g2_xnor2_1 _10824_ (.Y(_05916_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .B(\soc_inst.core_instr_addr[6] ));
 sg13g2_xor2_1 _10825_ (.B(\soc_inst.core_instr_addr[2] ),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .X(_05917_));
 sg13g2_xor2_1 _10826_ (.B(\soc_inst.core_instr_addr[13] ),
    .A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .X(_05918_));
 sg13g2_xor2_1 _10827_ (.B(\soc_inst.core_instr_addr[5] ),
    .A(\soc_inst.mem_ctrl.spi_addr[5] ),
    .X(_05919_));
 sg13g2_xnor2_1 _10828_ (.Y(_05920_),
    .A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .B(\soc_inst.core_instr_addr[3] ));
 sg13g2_xor2_1 _10829_ (.B(\soc_inst.core_instr_addr[8] ),
    .A(\soc_inst.mem_ctrl.spi_addr[8] ),
    .X(_05921_));
 sg13g2_xor2_1 _10830_ (.B(\soc_inst.core_instr_addr[10] ),
    .A(\soc_inst.mem_ctrl.spi_addr[10] ),
    .X(_05922_));
 sg13g2_xor2_1 _10831_ (.B(\soc_inst.core_instr_addr[23] ),
    .A(\soc_inst.mem_ctrl.spi_addr[23] ),
    .X(_05923_));
 sg13g2_a21oi_1 _10832_ (.A1(_05463_),
    .A2(\soc_inst.core_instr_addr[22] ),
    .Y(_05924_),
    .B1(_05923_));
 sg13g2_xor2_1 _10833_ (.B(\soc_inst.core_instr_addr[4] ),
    .A(\soc_inst.mem_ctrl.spi_addr[4] ),
    .X(_05925_));
 sg13g2_xor2_1 _10834_ (.B(\soc_inst.core_instr_addr[0] ),
    .A(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .X(_05926_));
 sg13g2_xor2_1 _10835_ (.B(\soc_inst.core_instr_addr[17] ),
    .A(\soc_inst.mem_ctrl.spi_addr[17] ),
    .X(_05927_));
 sg13g2_xor2_1 _10836_ (.B(\soc_inst.core_instr_addr[11] ),
    .A(\soc_inst.mem_ctrl.spi_addr[11] ),
    .X(_05928_));
 sg13g2_inv_1 _10837_ (.Y(_05929_),
    .A(_05928_));
 sg13g2_xnor2_1 _10838_ (.Y(_05930_),
    .A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .B(\soc_inst.core_instr_addr[21] ));
 sg13g2_xor2_1 _10839_ (.B(\soc_inst.core_instr_addr[12] ),
    .A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .X(_05931_));
 sg13g2_xnor2_1 _10840_ (.Y(_05932_),
    .A(\soc_inst.mem_ctrl.spi_addr[19] ),
    .B(\soc_inst.core_instr_addr[19] ));
 sg13g2_nand2_1 _10841_ (.Y(_05933_),
    .A(\soc_inst.mem_ctrl.spi_addr[22] ),
    .B(_05464_));
 sg13g2_xor2_1 _10842_ (.B(\soc_inst.core_instr_addr[18] ),
    .A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .X(_05934_));
 sg13g2_xor2_1 _10843_ (.B(\soc_inst.core_instr_addr[9] ),
    .A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .X(_05935_));
 sg13g2_inv_1 _10844_ (.Y(_05936_),
    .A(_05935_));
 sg13g2_nor2_1 _10845_ (.A(_05921_),
    .B(_05925_),
    .Y(_05937_));
 sg13g2_nor4_1 _10846_ (.A(_05911_),
    .B(_05915_),
    .C(_05926_),
    .D(_05927_),
    .Y(_05938_));
 sg13g2_nor4_1 _10847_ (.A(_05912_),
    .B(_05917_),
    .C(_05922_),
    .D(_05934_),
    .Y(_05939_));
 sg13g2_nand4_1 _10848_ (.B(_05937_),
    .C(_05938_),
    .A(_05913_),
    .Y(_05940_),
    .D(_05939_));
 sg13g2_nand4_1 _10849_ (.B(_05930_),
    .C(_05932_),
    .A(_05929_),
    .Y(_05941_),
    .D(_05936_));
 sg13g2_nor4_1 _10850_ (.A(_05914_),
    .B(_05918_),
    .C(_05919_),
    .D(_05931_),
    .Y(_05942_));
 sg13g2_nand2_1 _10851_ (.Y(_05943_),
    .A(_05916_),
    .B(_05933_));
 sg13g2_nor2_1 _10852_ (.A(_05910_),
    .B(_05943_),
    .Y(_05944_));
 sg13g2_nand4_1 _10853_ (.B(_05924_),
    .C(_05942_),
    .A(_05920_),
    .Y(_05945_),
    .D(_05944_));
 sg13g2_nor3_2 _10854_ (.A(_05940_),
    .B(_05941_),
    .C(_05945_),
    .Y(_05946_));
 sg13g2_nand2_2 _10855_ (.Y(_05947_),
    .A(net641),
    .B(_05946_));
 sg13g2_nor2_1 _10856_ (.A(_05870_),
    .B(_05947_),
    .Y(_05948_));
 sg13g2_nand2_1 _10857_ (.Y(_05949_),
    .A(_05866_),
    .B(_05948_));
 sg13g2_o21ai_1 _10858_ (.B1(_05949_),
    .Y(_05950_),
    .A1(net2808),
    .A2(net4066));
 sg13g2_nor2b_1 _10859_ (.A(_05950_),
    .B_N(_05909_),
    .Y(_00332_));
 sg13g2_nor2_1 _10860_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .B(net2203),
    .Y(_05951_));
 sg13g2_nor3_1 _10861_ (.A(net5061),
    .B(net5123),
    .C(net2204),
    .Y(_00331_));
 sg13g2_and2_1 _10862_ (.A(net330),
    .B(net2211),
    .X(_05952_));
 sg13g2_a221oi_1 _10863_ (.B2(net1969),
    .C1(_05952_),
    .B1(net357),
    .A1(net513),
    .Y(_05953_),
    .A2(net2178));
 sg13g2_a22oi_1 _10864_ (.Y(_05954_),
    .B1(net562),
    .B2(net2169),
    .A2(net2101),
    .A1(net483));
 sg13g2_a22oi_1 _10865_ (.Y(_05955_),
    .B1(net380),
    .B2(net2409),
    .A2(net2150),
    .A1(net467));
 sg13g2_nand3_1 _10866_ (.B(_05954_),
    .C(_05955_),
    .A(_05953_),
    .Y(_00069_));
 sg13g2_and2_1 _10867_ (.A(\soc_inst.core_instr_data[0] ),
    .B(net5113),
    .X(_05956_));
 sg13g2_a21o_2 _10868_ (.A2(\soc_inst.core_instr_data[1] ),
    .A1(\soc_inst.core_instr_data[0] ),
    .B1(\soc_inst.mem_ctrl.spi_addr[1] ),
    .X(_05957_));
 sg13g2_nand2_1 _10869_ (.Y(_05958_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .B(_05957_));
 sg13g2_nand3_1 _10870_ (.B(\soc_inst.mem_ctrl.spi_addr[3] ),
    .C(_05957_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .Y(_05959_));
 sg13g2_nand4_1 _10871_ (.B(\soc_inst.mem_ctrl.spi_addr[3] ),
    .C(\soc_inst.mem_ctrl.spi_addr[4] ),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .Y(_05960_),
    .D(_05957_));
 sg13g2_nor2_2 _10872_ (.A(_05441_),
    .B(_05960_),
    .Y(_05961_));
 sg13g2_nand2_1 _10873_ (.Y(_05962_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .B(_05961_));
 sg13g2_nand3_1 _10874_ (.B(\soc_inst.mem_ctrl.spi_addr[7] ),
    .C(_05961_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .Y(_05963_));
 sg13g2_nand4_1 _10875_ (.B(\soc_inst.mem_ctrl.spi_addr[7] ),
    .C(\soc_inst.mem_ctrl.spi_addr[8] ),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .Y(_05964_),
    .D(_05961_));
 sg13g2_nor2_1 _10876_ (.A(_05447_),
    .B(_05964_),
    .Y(_05965_));
 sg13g2_nor4_2 _10877_ (.A(_05447_),
    .B(_05449_),
    .C(_05451_),
    .Y(_05966_),
    .D(_05964_));
 sg13g2_nand2_1 _10878_ (.Y(_05967_),
    .A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .B(_05966_));
 sg13g2_nand3_1 _10879_ (.B(\soc_inst.mem_ctrl.spi_addr[13] ),
    .C(_05966_),
    .A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .Y(_05968_));
 sg13g2_and4_1 _10880_ (.A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .B(\soc_inst.mem_ctrl.spi_addr[13] ),
    .C(\soc_inst.mem_ctrl.spi_addr[14] ),
    .D(_05966_),
    .X(_05969_));
 sg13g2_and2_1 _10881_ (.A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .B(_05969_),
    .X(_05970_));
 sg13g2_nand2_1 _10882_ (.Y(_05971_),
    .A(\soc_inst.mem_ctrl.spi_addr[16] ),
    .B(_05970_));
 sg13g2_and3_2 _10883_ (.X(_05972_),
    .A(\soc_inst.mem_ctrl.spi_addr[16] ),
    .B(\soc_inst.mem_ctrl.spi_addr[17] ),
    .C(_05970_));
 sg13g2_nand2_1 _10884_ (.Y(_05973_),
    .A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .B(_05972_));
 sg13g2_nand3_1 _10885_ (.B(\soc_inst.mem_ctrl.spi_addr[19] ),
    .C(_05972_),
    .A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .Y(_05974_));
 sg13g2_and4_1 _10886_ (.A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .B(\soc_inst.mem_ctrl.spi_addr[19] ),
    .C(\soc_inst.mem_ctrl.spi_addr[20] ),
    .D(_05972_),
    .X(_05975_));
 sg13g2_nand2_1 _10887_ (.Y(_05976_),
    .A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .B(_05975_));
 sg13g2_o21ai_1 _10888_ (.B1(_05933_),
    .Y(_05977_),
    .A1(_05923_),
    .A2(_05976_));
 sg13g2_o21ai_1 _10889_ (.B1(_05977_),
    .Y(_05978_),
    .A1(_05924_),
    .A2(_05976_));
 sg13g2_or2_1 _10890_ (.X(_05979_),
    .B(_05977_),
    .A(_05924_));
 sg13g2_xor2_1 _10891_ (.B(_05974_),
    .A(_05915_),
    .X(_05980_));
 sg13g2_xnor2_1 _10892_ (.Y(_05981_),
    .A(_05932_),
    .B(_05973_));
 sg13g2_xnor2_1 _10893_ (.Y(_05982_),
    .A(_05934_),
    .B(_05972_));
 sg13g2_xnor2_1 _10894_ (.Y(_05983_),
    .A(_05927_),
    .B(_05971_));
 sg13g2_xor2_1 _10895_ (.B(_05970_),
    .A(_05912_),
    .X(_05984_));
 sg13g2_xor2_1 _10896_ (.B(_05969_),
    .A(_05914_),
    .X(_05985_));
 sg13g2_xnor2_1 _10897_ (.Y(_05986_),
    .A(_05913_),
    .B(_05968_));
 sg13g2_xor2_1 _10898_ (.B(_05967_),
    .A(_05918_),
    .X(_05987_));
 sg13g2_xor2_1 _10899_ (.B(_05966_),
    .A(_05931_),
    .X(_05988_));
 sg13g2_a21oi_1 _10900_ (.A1(\soc_inst.mem_ctrl.spi_addr[10] ),
    .A2(_05965_),
    .Y(_05989_),
    .B1(_05929_));
 sg13g2_o21ai_1 _10901_ (.B1(_05910_),
    .Y(_05990_),
    .A1(\soc_inst.core_instr_addr[7] ),
    .A2(_05921_));
 sg13g2_nor2b_1 _10902_ (.A(_05962_),
    .B_N(_05990_),
    .Y(_05991_));
 sg13g2_xor2_1 _10903_ (.B(_05958_),
    .A(_05920_),
    .X(_05992_));
 sg13g2_nor2_1 _10904_ (.A(_05911_),
    .B(_05956_),
    .Y(_05993_));
 sg13g2_xnor2_1 _10905_ (.Y(_05994_),
    .A(_05917_),
    .B(_05957_));
 sg13g2_xnor2_1 _10906_ (.Y(_05995_),
    .A(_05919_),
    .B(_05960_));
 sg13g2_or2_1 _10907_ (.X(_05996_),
    .B(_05975_),
    .A(_05930_));
 sg13g2_o21ai_1 _10908_ (.B1(_05922_),
    .Y(_05997_),
    .A1(\soc_inst.core_instr_addr[10] ),
    .A2(_05928_));
 sg13g2_mux2_1 _10909_ (.A0(_05922_),
    .A1(_05997_),
    .S(_05965_),
    .X(_05998_));
 sg13g2_xnor2_1 _10910_ (.Y(_05999_),
    .A(_05936_),
    .B(_05964_));
 sg13g2_o21ai_1 _10911_ (.B1(_05994_),
    .Y(_06000_),
    .A1(_05925_),
    .A2(_05959_));
 sg13g2_a221oi_1 _10912_ (.B2(_05921_),
    .C1(_06000_),
    .B1(_05963_),
    .A1(_05916_),
    .Y(_06001_),
    .A2(_05961_));
 sg13g2_a21o_1 _10913_ (.A2(_05956_),
    .A1(_05911_),
    .B1(_05926_),
    .X(_06002_));
 sg13g2_nor4_1 _10914_ (.A(_05991_),
    .B(_05992_),
    .C(_05995_),
    .D(_06002_),
    .Y(_06003_));
 sg13g2_a21oi_1 _10915_ (.A1(_05925_),
    .A2(_05959_),
    .Y(_06004_),
    .B1(_05993_));
 sg13g2_o21ai_1 _10916_ (.B1(_06004_),
    .Y(_06005_),
    .A1(_05916_),
    .A2(_05961_));
 sg13g2_a21oi_1 _10917_ (.A1(_05910_),
    .A2(_05962_),
    .Y(_06006_),
    .B1(_06005_));
 sg13g2_nand4_1 _10918_ (.B(_06001_),
    .C(_06003_),
    .A(_05999_),
    .Y(_06007_),
    .D(_06006_));
 sg13g2_nor4_1 _10919_ (.A(_05988_),
    .B(_05989_),
    .C(_05998_),
    .D(_06007_),
    .Y(_06008_));
 sg13g2_nand3_1 _10920_ (.B(_05987_),
    .C(_06008_),
    .A(_05986_),
    .Y(_06009_));
 sg13g2_nor4_1 _10921_ (.A(_05983_),
    .B(_05984_),
    .C(_05985_),
    .D(_06009_),
    .Y(_06010_));
 sg13g2_nand4_1 _10922_ (.B(_05981_),
    .C(_05982_),
    .A(_05980_),
    .Y(_06011_),
    .D(_06010_));
 sg13g2_a21oi_1 _10923_ (.A1(_05930_),
    .A2(_05975_),
    .Y(_06012_),
    .B1(_06011_));
 sg13g2_and4_1 _10924_ (.A(_05978_),
    .B(_05979_),
    .C(_05996_),
    .D(_06012_),
    .X(_06013_));
 sg13g2_nor3_1 _10925_ (.A(_05467_),
    .B(_05946_),
    .C(_06013_),
    .Y(_06014_));
 sg13g2_nor3_1 _10926_ (.A(_05466_),
    .B(_05946_),
    .C(_06013_),
    .Y(_06015_));
 sg13g2_nor3_1 _10927_ (.A(_05871_),
    .B(_06014_),
    .C(_06015_),
    .Y(_06016_));
 sg13g2_nor2_1 _10928_ (.A(net4015),
    .B(_06016_),
    .Y(_00089_));
 sg13g2_a21o_1 _10929_ (.A2(net4015),
    .A1(net2748),
    .B1(_00089_),
    .X(_00009_));
 sg13g2_or3_1 _10930_ (.A(net2808),
    .B(_05907_),
    .C(_05948_),
    .X(_06017_));
 sg13g2_inv_1 _10931_ (.Y(_00088_),
    .A(_06017_));
 sg13g2_nor2_1 _10932_ (.A(_05469_),
    .B(\soc_inst.mem_ctrl.spi_done ),
    .Y(_06018_));
 sg13g2_a21oi_1 _10933_ (.A1(_05872_),
    .A2(_06018_),
    .Y(_06019_),
    .B1(net4015));
 sg13g2_o21ai_1 _10934_ (.B1(_06017_),
    .Y(_00008_),
    .A1(_05469_),
    .A2(_06019_));
 sg13g2_nor2_1 _10935_ (.A(net5120),
    .B(\soc_inst.i2c_inst.state[1] ),
    .Y(_06020_));
 sg13g2_or2_1 _10936_ (.X(_06021_),
    .B(\soc_inst.i2c_inst.state[1] ),
    .A(net5120));
 sg13g2_nor2_1 _10937_ (.A(net5115),
    .B(_06021_),
    .Y(_06022_));
 sg13g2_nor3_2 _10938_ (.A(net2936),
    .B(net5119),
    .C(_06021_),
    .Y(_06023_));
 sg13g2_inv_2 _10939_ (.Y(\soc_inst.i2c_ena ),
    .A(_06023_));
 sg13g2_o21ai_1 _10940_ (.B1(net4779),
    .Y(_06024_),
    .A1(_05946_),
    .A2(_06013_));
 sg13g2_inv_1 _10941_ (.Y(_06025_),
    .A(_06024_));
 sg13g2_nor2_1 _10942_ (.A(net2735),
    .B(_06024_),
    .Y(_06026_));
 sg13g2_nand2_1 _10943_ (.Y(_06027_),
    .A(net4772),
    .B(_06013_));
 sg13g2_and3_1 _10944_ (.X(_06028_),
    .A(net4772),
    .B(net403),
    .C(_06013_));
 sg13g2_o21ai_1 _10945_ (.B1(_05906_),
    .Y(_06029_),
    .A1(_06026_),
    .A2(_06028_));
 sg13g2_nand4_1 _10946_ (.B(net2566),
    .C(net2735),
    .A(net5074),
    .Y(_06030_),
    .D(_05869_));
 sg13g2_nand2_1 _10947_ (.Y(_06031_),
    .A(net4779),
    .B(net4015));
 sg13g2_nand3_1 _10948_ (.B(_06030_),
    .C(_06031_),
    .A(_06029_),
    .Y(_00006_));
 sg13g2_nor2_1 _10949_ (.A(net403),
    .B(_06027_),
    .Y(_06032_));
 sg13g2_a21o_1 _10950_ (.A2(_06025_),
    .A1(net2735),
    .B1(_06032_),
    .X(_06033_));
 sg13g2_nand2_1 _10951_ (.Y(_06034_),
    .A(_05872_),
    .B(_05946_));
 sg13g2_nand2_1 _10952_ (.Y(_06035_),
    .A(net4066),
    .B(_06034_));
 sg13g2_a22oi_1 _10953_ (.Y(_06036_),
    .B1(_06035_),
    .B2(net4772),
    .A2(_06033_),
    .A1(_05906_));
 sg13g2_inv_1 _10954_ (.Y(_00007_),
    .A(_06036_));
 sg13g2_nor2_1 _10955_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .B(_05492_),
    .Y(_06037_));
 sg13g2_nor2_2 _10956_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .B(net5059),
    .Y(_06038_));
 sg13g2_nor3_1 _10957_ (.A(net4782),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .C(net5059),
    .Y(_06039_));
 sg13g2_nor2_1 _10958_ (.A(net4782),
    .B(net4784),
    .Y(_06040_));
 sg13g2_nor3_2 _10959_ (.A(net4782),
    .B(net4784),
    .C(net2899),
    .Y(_06041_));
 sg13g2_nand3_1 _10960_ (.B(_06038_),
    .C(_06041_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .Y(_06042_));
 sg13g2_nand2_1 _10961_ (.Y(_06043_),
    .A(net5072),
    .B(_06042_));
 sg13g2_a21oi_1 _10962_ (.A1(net5072),
    .A2(_06042_),
    .Y(_06044_),
    .B1(net2215));
 sg13g2_and2_1 _10963_ (.A(_05434_),
    .B(_05878_),
    .X(_06045_));
 sg13g2_a21oi_2 _10964_ (.B1(net5074),
    .Y(_06046_),
    .A2(_06045_),
    .A1(_05879_));
 sg13g2_a21o_1 _10965_ (.A2(_06045_),
    .A1(_05879_),
    .B1(net5074),
    .X(_06047_));
 sg13g2_nand2_2 _10966_ (.Y(_06048_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .B(net408));
 sg13g2_nor3_2 _10967_ (.A(net5123),
    .B(net5073),
    .C(net409),
    .Y(_06049_));
 sg13g2_inv_1 _10968_ (.Y(_06050_),
    .A(_06049_));
 sg13g2_nand3b_1 _10969_ (.B(net4278),
    .C(net410),
    .Y(_06051_),
    .A_N(net334));
 sg13g2_o21ai_1 _10970_ (.B1(_06051_),
    .Y(_00013_),
    .A1(net5123),
    .A2(net2216));
 sg13g2_nand2b_1 _10971_ (.Y(_06052_),
    .B(net520),
    .A_N(\soc_inst.spi_inst.state[0] ));
 sg13g2_xor2_1 _10972_ (.B(net2298),
    .A(net520),
    .X(_00123_));
 sg13g2_nor2b_1 _10973_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .Y(_06053_));
 sg13g2_nor2_1 _10974_ (.A(_05376_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .Y(_06054_));
 sg13g2_nor2_1 _10975_ (.A(_05375_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .Y(_06055_));
 sg13g2_or4_1 _10976_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .B(_06053_),
    .C(_06054_),
    .D(_06055_),
    .X(_06056_));
 sg13g2_xnor2_1 _10977_ (.Y(_06057_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .B(_00329_));
 sg13g2_xnor2_1 _10978_ (.Y(_06058_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .B(_00327_));
 sg13g2_nor2_1 _10979_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .B(_05412_),
    .Y(_06059_));
 sg13g2_nor2b_1 _10980_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .B_N(net4759),
    .Y(_06060_));
 sg13g2_a221oi_1 _10981_ (.B2(_05376_),
    .C1(_06060_),
    .B1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .Y(_06061_),
    .A2(net4758));
 sg13g2_nor2_1 _10982_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .B(net4758),
    .Y(_06062_));
 sg13g2_nor2b_1 _10983_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .Y(_06063_));
 sg13g2_nor2_1 _10984_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .B(_00328_),
    .Y(_06064_));
 sg13g2_nor2b_1 _10985_ (.A(net4759),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .Y(_06065_));
 sg13g2_nor4_1 _10986_ (.A(_06062_),
    .B(_06063_),
    .C(_06064_),
    .D(_06065_),
    .Y(_06066_));
 sg13g2_nor2_1 _10987_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .B(_05413_),
    .Y(_06067_));
 sg13g2_a21oi_1 _10988_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .A2(_00328_),
    .Y(_06068_),
    .B1(_06067_));
 sg13g2_nor2_1 _10989_ (.A(_05374_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .Y(_06069_));
 sg13g2_nor2b_1 _10990_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .Y(_06070_));
 sg13g2_nor2_1 _10991_ (.A(_06069_),
    .B(_06070_),
    .Y(_06071_));
 sg13g2_nand4_1 _10992_ (.B(_06066_),
    .C(_06068_),
    .A(_06061_),
    .Y(_06072_),
    .D(_06071_));
 sg13g2_nor4_1 _10993_ (.A(_06056_),
    .B(_06057_),
    .C(_06058_),
    .D(_06072_),
    .Y(_06073_));
 sg13g2_xor2_1 _10994_ (.B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .X(_06074_));
 sg13g2_nand2b_1 _10995_ (.Y(_06075_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .A_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ));
 sg13g2_o21ai_1 _10996_ (.B1(_06075_),
    .Y(_06076_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .A2(_05411_));
 sg13g2_xnor2_1 _10997_ (.Y(_06077_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ));
 sg13g2_xor2_1 _10998_ (.B(_00329_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .X(_06078_));
 sg13g2_nand2_1 _10999_ (.Y(_06079_),
    .A(_06077_),
    .B(_06078_));
 sg13g2_a22oi_1 _11000_ (.Y(_06080_),
    .B1(net4759),
    .B2(_05374_),
    .A2(_00327_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ));
 sg13g2_a22oi_1 _11001_ (.Y(_06081_),
    .B1(_05413_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .A2(net4758),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ));
 sg13g2_nor2_1 _11002_ (.A(_05374_),
    .B(net4759),
    .Y(_06082_));
 sg13g2_nor2_1 _11003_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .B(_00328_),
    .Y(_06083_));
 sg13g2_or2_1 _11004_ (.X(_06084_),
    .B(_00327_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ));
 sg13g2_o21ai_1 _11005_ (.B1(_06084_),
    .Y(_06085_),
    .A1(_05375_),
    .A2(_05389_));
 sg13g2_nor3_1 _11006_ (.A(_06082_),
    .B(_06083_),
    .C(_06085_),
    .Y(_06086_));
 sg13g2_nor2b_1 _11007_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .Y(_06087_));
 sg13g2_nor2_1 _11008_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .B(net4758),
    .Y(_06088_));
 sg13g2_nor2_1 _11009_ (.A(_05376_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .Y(_06089_));
 sg13g2_nor2b_1 _11010_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .Y(_06090_));
 sg13g2_nor4_1 _11011_ (.A(_06087_),
    .B(_06088_),
    .C(_06089_),
    .D(_06090_),
    .Y(_06091_));
 sg13g2_nand4_1 _11012_ (.B(_06081_),
    .C(_06086_),
    .A(_06080_),
    .Y(_06092_),
    .D(_06091_));
 sg13g2_nor4_1 _11013_ (.A(_06074_),
    .B(_06076_),
    .C(_06079_),
    .D(_06092_),
    .Y(_06093_));
 sg13g2_xnor2_1 _11014_ (.Y(_06094_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .B(_00328_));
 sg13g2_nor4_1 _11015_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .B(_06057_),
    .C(_06069_),
    .D(_06094_),
    .Y(_06095_));
 sg13g2_nor3_1 _11016_ (.A(_06053_),
    .B(_06055_),
    .C(_06065_),
    .Y(_06096_));
 sg13g2_nor4_1 _11017_ (.A(_06054_),
    .B(_06060_),
    .C(_06067_),
    .D(_06070_),
    .Y(_06097_));
 sg13g2_xnor2_1 _11018_ (.Y(_06098_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .B(net4758));
 sg13g2_nor4_1 _11019_ (.A(_06058_),
    .B(_06059_),
    .C(_06063_),
    .D(_06098_),
    .Y(_06099_));
 sg13g2_and4_1 _11020_ (.A(_06095_),
    .B(_06096_),
    .C(_06097_),
    .D(_06099_),
    .X(_06100_));
 sg13g2_a22oi_1 _11021_ (.Y(_06101_),
    .B1(_05413_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .A2(net4759),
    .A1(_05374_));
 sg13g2_xor2_1 _11022_ (.B(_00328_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .X(_06102_));
 sg13g2_nand3_1 _11023_ (.B(_06101_),
    .C(_06102_),
    .A(_06077_),
    .Y(_06103_));
 sg13g2_nor3_1 _11024_ (.A(_06076_),
    .B(_06087_),
    .C(_06089_),
    .Y(_06104_));
 sg13g2_nor3_1 _11025_ (.A(_06082_),
    .B(_06088_),
    .C(_06090_),
    .Y(_06105_));
 sg13g2_nand2_1 _11026_ (.Y(_06106_),
    .A(_06104_),
    .B(_06105_));
 sg13g2_a22oi_1 _11027_ (.Y(_06107_),
    .B1(_00327_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .A2(net4758),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ));
 sg13g2_nand3_1 _11028_ (.B(_06084_),
    .C(_06107_),
    .A(_06078_),
    .Y(_06108_));
 sg13g2_nor4_1 _11029_ (.A(_06074_),
    .B(_06103_),
    .C(_06106_),
    .D(_06108_),
    .Y(_06109_));
 sg13g2_a21o_2 _11030_ (.A2(_06100_),
    .A1(net4762),
    .B1(_06109_),
    .X(_06110_));
 sg13g2_inv_1 _11031_ (.Y(_06111_),
    .A(_06110_));
 sg13g2_nand2_2 _11032_ (.Y(_06112_),
    .A(net5436),
    .B(_06111_));
 sg13g2_inv_1 _11033_ (.Y(_06113_),
    .A(_06112_));
 sg13g2_nor4_1 _11034_ (.A(_05377_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ),
    .C(net522),
    .D(net2124),
    .Y(_06114_));
 sg13g2_nand2_1 _11035_ (.Y(_06115_),
    .A(net5470),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ));
 sg13g2_nand3_1 _11036_ (.B(net1120),
    .C(net2125),
    .A(net5470),
    .Y(_06116_));
 sg13g2_o21ai_1 _11037_ (.B1(_06116_),
    .Y(_00022_),
    .A1(_05386_),
    .A2(_06112_));
 sg13g2_nor2b_1 _11038_ (.A(net1698),
    .B_N(net1114),
    .Y(_06117_));
 sg13g2_a22oi_1 _11039_ (.Y(_06118_),
    .B1(_06117_),
    .B2(net5470),
    .A2(_06113_),
    .A1(net938));
 sg13g2_inv_1 _11040_ (.Y(_00021_),
    .A(_06118_));
 sg13g2_nand3_1 _11041_ (.B(net938),
    .C(_06110_),
    .A(net5470),
    .Y(_06119_));
 sg13g2_o21ai_1 _11042_ (.B1(_06119_),
    .Y(_00020_),
    .A1(_06114_),
    .A2(_06115_));
 sg13g2_nand2_1 _11043_ (.Y(_06120_),
    .A(net1698),
    .B(net1114));
 sg13g2_o21ai_1 _11044_ (.B1(net4762),
    .Y(_06121_),
    .A1(_06073_),
    .A2(_06093_));
 sg13g2_nand3_1 _11045_ (.B(_06120_),
    .C(_06121_),
    .A(net5473),
    .Y(_00019_));
 sg13g2_nand2_1 _11046_ (.Y(_06122_),
    .A(net5064),
    .B(_06042_));
 sg13g2_a21oi_1 _11047_ (.A1(net5064),
    .A2(_06042_),
    .Y(_06123_),
    .B1(net504));
 sg13g2_nand3_1 _11048_ (.B(net4280),
    .C(net410),
    .A(net91),
    .Y(_06124_));
 sg13g2_o21ai_1 _11049_ (.B1(_06124_),
    .Y(_00011_),
    .A1(net5123),
    .A2(net505));
 sg13g2_nor2_1 _11050_ (.A(_05491_),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .Y(_06125_));
 sg13g2_nand3_1 _11051_ (.B(_06038_),
    .C(_06125_),
    .A(net2926),
    .Y(_06126_));
 sg13g2_nor2_1 _11052_ (.A(net4784),
    .B(_06126_),
    .Y(_06127_));
 sg13g2_o21ai_1 _11053_ (.B1(net5065),
    .Y(_06128_),
    .A1(net4784),
    .A2(_06126_));
 sg13g2_nand4_1 _11054_ (.B(_05493_),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ),
    .A(net2868),
    .Y(_06129_),
    .D(_06041_));
 sg13g2_nor2_1 _11055_ (.A(_05497_),
    .B(_06129_),
    .Y(_06130_));
 sg13g2_nand2_1 _11056_ (.Y(_06131_),
    .A(_05417_),
    .B(net2945));
 sg13g2_a21oi_1 _11057_ (.A1(net2953),
    .A2(_06131_),
    .Y(_00010_),
    .B1(net5123));
 sg13g2_nand4_1 _11058_ (.B(net4783),
    .C(_06038_),
    .A(net4782),
    .Y(_06132_),
    .D(_06125_));
 sg13g2_a21oi_1 _11059_ (.A1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .A2(_06132_),
    .Y(_06133_),
    .B1(net430));
 sg13g2_nand2b_1 _11060_ (.Y(_06134_),
    .B(net1034),
    .A_N(net5121));
 sg13g2_nor2_1 _11061_ (.A(net5121),
    .B(net431),
    .Y(_00018_));
 sg13g2_nand4_1 _11062_ (.B(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .C(net397),
    .A(net460),
    .Y(_06135_),
    .D(net401));
 sg13g2_nand4_1 _11063_ (.B(net368),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ),
    .A(net303),
    .Y(_06136_),
    .D(net144));
 sg13g2_nor2b_1 _11064_ (.A(net408),
    .B_N(net2740),
    .Y(_06137_));
 sg13g2_nand4_1 _11065_ (.B(net217),
    .C(net418),
    .A(net245),
    .Y(_06138_),
    .D(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ));
 sg13g2_or3_1 _11066_ (.A(_06135_),
    .B(_06136_),
    .C(_06138_),
    .X(_06139_));
 sg13g2_a22oi_1 _11067_ (.Y(_06140_),
    .B1(_06139_),
    .B2(net2578),
    .A2(_06137_),
    .A1(_05865_));
 sg13g2_nor2_1 _11068_ (.A(net5121),
    .B(_06140_),
    .Y(_00017_));
 sg13g2_nand3_1 _11069_ (.B(_06037_),
    .C(_06039_),
    .A(net4783),
    .Y(_06141_));
 sg13g2_nand2_1 _11070_ (.Y(_06142_),
    .A(net496),
    .B(_06141_));
 sg13g2_a21oi_1 _11071_ (.A1(_05499_),
    .A2(_06142_),
    .Y(_00016_),
    .B1(net5122));
 sg13g2_xnor2_1 _11072_ (.Y(_06143_),
    .A(net2373),
    .B(net2723));
 sg13g2_xnor2_1 _11073_ (.Y(_06144_),
    .A(net2868),
    .B(net2759));
 sg13g2_xnor2_1 _11074_ (.Y(_06145_),
    .A(net5059),
    .B(net2741));
 sg13g2_nand4_1 _11075_ (.B(_06143_),
    .C(_06144_),
    .A(_06041_),
    .Y(_06146_),
    .D(_06145_));
 sg13g2_nor3_1 _11076_ (.A(net5124),
    .B(net5076),
    .C(_05495_),
    .Y(_06147_));
 sg13g2_nand2_1 _11077_ (.Y(_06148_),
    .A(_06146_),
    .B(_06147_));
 sg13g2_and2_1 _11078_ (.A(net5076),
    .B(net5066),
    .X(_06149_));
 sg13g2_a221oi_1 _11079_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .C1(_06149_),
    .B1(net2945),
    .A1(net5065),
    .Y(_06150_),
    .A2(_06127_));
 sg13g2_o21ai_1 _11080_ (.B1(_06148_),
    .Y(_00015_),
    .A1(net5123),
    .A2(net2946));
 sg13g2_nor2_2 _11081_ (.A(_05491_),
    .B(_05492_),
    .Y(_06151_));
 sg13g2_nand3_1 _11082_ (.B(_06039_),
    .C(_06151_),
    .A(net4783),
    .Y(_06152_));
 sg13g2_nand3b_1 _11083_ (.B(net474),
    .C(_06152_),
    .Y(_06153_),
    .A_N(net5122));
 sg13g2_o21ai_1 _11084_ (.B1(_06153_),
    .Y(_00014_),
    .A1(_06132_),
    .A2(_06134_));
 sg13g2_or2_1 _11085_ (.X(_06154_),
    .B(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .A(_00292_));
 sg13g2_o21ai_1 _11086_ (.B1(_06154_),
    .Y(_06155_),
    .A1(_00291_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[46] ));
 sg13g2_or2_1 _11087_ (.X(_06156_),
    .B(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .A(_00290_));
 sg13g2_o21ai_1 _11088_ (.B1(_06156_),
    .Y(_06157_),
    .A1(_00289_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[44] ));
 sg13g2_a22oi_1 _11089_ (.Y(_06158_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .B2(_00288_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .A1(_00289_));
 sg13g2_or2_1 _11090_ (.X(_06159_),
    .B(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .A(_00288_));
 sg13g2_nand2_1 _11091_ (.Y(_06160_),
    .A(net1421),
    .B(\soc_inst.cpu_core.csr_file.mtime[42] ));
 sg13g2_a22oi_1 _11092_ (.Y(_06161_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .B2(_00285_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .A1(_00286_));
 sg13g2_or2_1 _11093_ (.X(_06162_),
    .B(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .A(_00286_));
 sg13g2_o21ai_1 _11094_ (.B1(_06162_),
    .Y(_06163_),
    .A1(_00287_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[42] ));
 sg13g2_o21ai_1 _11095_ (.B1(_06160_),
    .Y(_06164_),
    .A1(_06161_),
    .A2(_06163_));
 sg13g2_nand2_1 _11096_ (.Y(_06165_),
    .A(_06159_),
    .B(_06164_));
 sg13g2_a21oi_1 _11097_ (.A1(_06158_),
    .A2(_06165_),
    .Y(_06166_),
    .B1(_06157_));
 sg13g2_a221oi_1 _11098_ (.B2(net1786),
    .C1(_06166_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .A1(_00291_),
    .Y(_06167_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[46] ));
 sg13g2_nand2_1 _11099_ (.Y(_06168_),
    .A(net1758),
    .B(net694));
 sg13g2_nor2_1 _11100_ (.A(net1464),
    .B(net1715),
    .Y(_06169_));
 sg13g2_nor2_1 _11101_ (.A(_00280_),
    .B(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .Y(_06170_));
 sg13g2_and2_1 _11102_ (.A(net1304),
    .B(net2958),
    .X(_06171_));
 sg13g2_a21oi_1 _11103_ (.A1(_00279_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .Y(_06172_),
    .B1(_06171_));
 sg13g2_a21oi_1 _11104_ (.A1(net1621),
    .A2(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .Y(_06173_),
    .B1(_06170_));
 sg13g2_o21ai_1 _11105_ (.B1(_06173_),
    .Y(_06174_),
    .A1(net1621),
    .A2(net2587));
 sg13g2_a22oi_1 _11106_ (.Y(_06175_),
    .B1(net2769),
    .B2(net1718),
    .A2(net1892),
    .A1(net1917));
 sg13g2_nor2_1 _11107_ (.A(net1917),
    .B(net1892),
    .Y(_06176_));
 sg13g2_or3_1 _11108_ (.A(_06174_),
    .B(_06175_),
    .C(_06176_),
    .X(_06177_));
 sg13g2_o21ai_1 _11109_ (.B1(_06177_),
    .Y(_06178_),
    .A1(_06170_),
    .A2(_06172_));
 sg13g2_nand2b_1 _11110_ (.Y(_06179_),
    .B(_06178_),
    .A_N(_06169_));
 sg13g2_a22oi_1 _11111_ (.Y(_06180_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .B2(net1425),
    .A2(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .A1(_00284_));
 sg13g2_a22oi_1 _11112_ (.Y(_06181_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .B2(net1464),
    .A2(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .A1(_00282_));
 sg13g2_nand2_1 _11113_ (.Y(_06182_),
    .A(_06180_),
    .B(_06181_));
 sg13g2_a221oi_1 _11114_ (.B2(_00290_),
    .C1(_06157_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .A1(_00291_),
    .Y(_06183_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[46] ));
 sg13g2_nand3_1 _11115_ (.B(_06161_),
    .C(_06183_),
    .A(_06158_),
    .Y(_06184_));
 sg13g2_or2_1 _11116_ (.X(_06185_),
    .B(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .A(_00285_));
 sg13g2_nand4_1 _11117_ (.B(_06160_),
    .C(_06168_),
    .A(_06159_),
    .Y(_06186_),
    .D(_06185_));
 sg13g2_nor4_2 _11118_ (.A(_06155_),
    .B(_06163_),
    .C(_06184_),
    .Y(_06187_),
    .D(_06186_));
 sg13g2_nor2_1 _11119_ (.A(net1964),
    .B(net1653),
    .Y(_06188_));
 sg13g2_or2_1 _11120_ (.X(_06189_),
    .B(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .A(_00283_));
 sg13g2_o21ai_1 _11121_ (.B1(_06189_),
    .Y(_06190_),
    .A1(net1838),
    .A2(net1855));
 sg13g2_a21o_1 _11122_ (.A2(_06181_),
    .A1(_06179_),
    .B1(_06190_),
    .X(_06191_));
 sg13g2_a21oi_1 _11123_ (.A1(_06180_),
    .A2(_06191_),
    .Y(_06192_),
    .B1(_06188_));
 sg13g2_o21ai_1 _11124_ (.B1(_06168_),
    .Y(_06193_),
    .A1(_06155_),
    .A2(_06167_));
 sg13g2_a21oi_1 _11125_ (.A1(_06187_),
    .A2(_06192_),
    .Y(_06194_),
    .B1(_06193_));
 sg13g2_or2_1 _11126_ (.X(_06195_),
    .B(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .A(_00326_));
 sg13g2_o21ai_1 _11127_ (.B1(_06195_),
    .Y(_06196_),
    .A1(_00325_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[30] ));
 sg13g2_a21o_1 _11128_ (.A2(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .A1(_00325_),
    .B1(_06196_),
    .X(_06197_));
 sg13g2_a22oi_1 _11129_ (.Y(_06198_),
    .B1(_05513_),
    .B2(_05395_),
    .A2(_05512_),
    .A1(_05394_));
 sg13g2_a22oi_1 _11130_ (.Y(_06199_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .B2(_00319_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .A1(_00320_));
 sg13g2_nor2_1 _11131_ (.A(_00321_),
    .B(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .Y(_06200_));
 sg13g2_nor2_1 _11132_ (.A(_00322_),
    .B(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .Y(_06201_));
 sg13g2_nand2_1 _11133_ (.Y(_06202_),
    .A(_00321_),
    .B(\soc_inst.cpu_core.csr_file.mtime[26] ));
 sg13g2_o21ai_1 _11134_ (.B1(_06202_),
    .Y(_06203_),
    .A1(_00320_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[25] ));
 sg13g2_or3_1 _11135_ (.A(_06200_),
    .B(_06201_),
    .C(_06203_),
    .X(_06204_));
 sg13g2_a22oi_1 _11136_ (.Y(_06205_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .B2(_00322_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .A1(_00323_));
 sg13g2_o21ai_1 _11137_ (.B1(_06205_),
    .Y(_06206_),
    .A1(_06201_),
    .A2(_06202_));
 sg13g2_inv_1 _11138_ (.Y(_06207_),
    .A(_06206_));
 sg13g2_o21ai_1 _11139_ (.B1(_06207_),
    .Y(_06208_),
    .A1(_06199_),
    .A2(_06204_));
 sg13g2_a22oi_1 _11140_ (.Y(_06209_),
    .B1(_06198_),
    .B2(_06208_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .A1(_00324_));
 sg13g2_and3_1 _11141_ (.X(_06210_),
    .A(_00325_),
    .B(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .C(_06195_));
 sg13g2_a21oi_1 _11142_ (.A1(_00326_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .Y(_06211_),
    .B1(_06210_));
 sg13g2_o21ai_1 _11143_ (.B1(_06211_),
    .Y(_06212_),
    .A1(_06197_),
    .A2(_06209_));
 sg13g2_or2_1 _11144_ (.X(_06213_),
    .B(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .A(_00318_));
 sg13g2_and2_1 _11145_ (.A(_00317_),
    .B(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .X(_06214_));
 sg13g2_o21ai_1 _11146_ (.B1(_06213_),
    .Y(_06215_),
    .A1(_00317_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[22] ));
 sg13g2_nor2_1 _11147_ (.A(_06214_),
    .B(_06215_),
    .Y(_06216_));
 sg13g2_or2_1 _11148_ (.X(_06217_),
    .B(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .A(_00315_));
 sg13g2_o21ai_1 _11149_ (.B1(_06217_),
    .Y(_06218_),
    .A1(_00316_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[21] ));
 sg13g2_a22oi_1 _11150_ (.Y(_06219_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .B2(_00314_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .A1(_00315_));
 sg13g2_nor2_1 _11151_ (.A(_00313_),
    .B(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .Y(_06220_));
 sg13g2_nor2_1 _11152_ (.A(_00314_),
    .B(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .Y(_06221_));
 sg13g2_nor2_1 _11153_ (.A(_06220_),
    .B(_06221_),
    .Y(_06222_));
 sg13g2_nand2_1 _11154_ (.Y(_06223_),
    .A(_00313_),
    .B(\soc_inst.cpu_core.csr_file.mtime[18] ));
 sg13g2_a22oi_1 _11155_ (.Y(_06224_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .B2(_00311_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .A1(_00312_));
 sg13g2_nor2_1 _11156_ (.A(_00312_),
    .B(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .Y(_06225_));
 sg13g2_o21ai_1 _11157_ (.B1(_06223_),
    .Y(_06226_),
    .A1(_06224_),
    .A2(_06225_));
 sg13g2_nand2_1 _11158_ (.Y(_06227_),
    .A(_06222_),
    .B(_06226_));
 sg13g2_a21oi_1 _11159_ (.A1(_06219_),
    .A2(_06227_),
    .Y(_06228_),
    .B1(_06218_));
 sg13g2_a21o_1 _11160_ (.A2(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .A1(_00316_),
    .B1(_06228_),
    .X(_06229_));
 sg13g2_a21o_1 _11161_ (.A2(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .A1(_00318_),
    .B1(_06214_),
    .X(_06230_));
 sg13g2_a22oi_1 _11162_ (.Y(_06231_),
    .B1(_06230_),
    .B2(_06213_),
    .A2(_06229_),
    .A1(_06216_));
 sg13g2_nor2_1 _11163_ (.A(_00301_),
    .B(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .Y(_06232_));
 sg13g2_or2_1 _11164_ (.X(_06233_),
    .B(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .A(_00296_));
 sg13g2_o21ai_1 _11165_ (.B1(_06233_),
    .Y(_06234_),
    .A1(_00295_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[0] ));
 sg13g2_a22oi_1 _11166_ (.Y(_06235_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .B2(_00297_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .A1(_00296_));
 sg13g2_a22oi_1 _11167_ (.Y(_06236_),
    .B1(_06234_),
    .B2(_06235_),
    .A2(_05508_),
    .A1(_05396_));
 sg13g2_o21ai_1 _11168_ (.B1(_06236_),
    .Y(_06237_),
    .A1(_00298_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[3] ));
 sg13g2_a22oi_1 _11169_ (.Y(_06238_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .B2(_00299_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .A1(_00298_));
 sg13g2_or2_1 _11170_ (.X(_06239_),
    .B(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .A(_00300_));
 sg13g2_o21ai_1 _11171_ (.B1(_06239_),
    .Y(_06240_),
    .A1(_00299_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[4] ));
 sg13g2_a21oi_1 _11172_ (.A1(_06237_),
    .A2(_06238_),
    .Y(_06241_),
    .B1(_06240_));
 sg13g2_a21oi_1 _11173_ (.A1(_00300_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .Y(_06242_),
    .B1(_06241_));
 sg13g2_a22oi_1 _11174_ (.Y(_06243_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .B2(_00301_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .A1(_00302_));
 sg13g2_o21ai_1 _11175_ (.B1(_06243_),
    .Y(_06244_),
    .A1(_06232_),
    .A2(_06242_));
 sg13g2_nor2_1 _11176_ (.A(_00302_),
    .B(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .Y(_06245_));
 sg13g2_o21ai_1 _11177_ (.B1(_06244_),
    .Y(_06246_),
    .A1(_00303_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[8] ));
 sg13g2_a22oi_1 _11178_ (.Y(_06247_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .B2(_00303_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .A1(_00304_));
 sg13g2_o21ai_1 _11179_ (.B1(_06247_),
    .Y(_06248_),
    .A1(_06245_),
    .A2(_06246_));
 sg13g2_nor2_1 _11180_ (.A(_00305_),
    .B(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .Y(_06249_));
 sg13g2_o21ai_1 _11181_ (.B1(_06248_),
    .Y(_06250_),
    .A1(_00304_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[9] ));
 sg13g2_a22oi_1 _11182_ (.Y(_06251_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .B2(_00305_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .A1(_00306_));
 sg13g2_o21ai_1 _11183_ (.B1(_06251_),
    .Y(_06252_),
    .A1(_06249_),
    .A2(_06250_));
 sg13g2_a22oi_1 _11184_ (.Y(_06253_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .B2(_00309_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .A1(_00310_));
 sg13g2_nor2_1 _11185_ (.A(_00310_),
    .B(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .Y(_06254_));
 sg13g2_o21ai_1 _11186_ (.B1(_06253_),
    .Y(_06255_),
    .A1(_00309_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[14] ));
 sg13g2_nor2_1 _11187_ (.A(_06254_),
    .B(_06255_),
    .Y(_06256_));
 sg13g2_and2_1 _11188_ (.A(_00308_),
    .B(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .X(_06257_));
 sg13g2_nand2_1 _11189_ (.Y(_06258_),
    .A(_00308_),
    .B(\soc_inst.cpu_core.csr_file.mtime[13] ));
 sg13g2_nor2_1 _11190_ (.A(_00308_),
    .B(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .Y(_06259_));
 sg13g2_nand2_1 _11191_ (.Y(_06260_),
    .A(_00307_),
    .B(\soc_inst.cpu_core.csr_file.mtime[12] ));
 sg13g2_o21ai_1 _11192_ (.B1(_06260_),
    .Y(_06261_),
    .A1(_00306_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[11] ));
 sg13g2_o21ai_1 _11193_ (.B1(_06256_),
    .Y(_06262_),
    .A1(_00307_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[12] ));
 sg13g2_nor4_1 _11194_ (.A(_06257_),
    .B(_06259_),
    .C(_06261_),
    .D(_06262_),
    .Y(_06263_));
 sg13g2_o21ai_1 _11195_ (.B1(_06258_),
    .Y(_06264_),
    .A1(_06259_),
    .A2(_06260_));
 sg13g2_nor2_1 _11196_ (.A(_06253_),
    .B(_06254_),
    .Y(_06265_));
 sg13g2_a221oi_1 _11197_ (.B2(_06256_),
    .C1(_06265_),
    .B1(_06264_),
    .A1(_06252_),
    .Y(_06266_),
    .A2(_06263_));
 sg13g2_or2_1 _11198_ (.X(_06267_),
    .B(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .A(_00311_));
 sg13g2_a21oi_1 _11199_ (.A1(_00318_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .Y(_06268_),
    .B1(_06225_));
 sg13g2_a221oi_1 _11200_ (.B2(_00313_),
    .C1(_06218_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .A1(_00316_),
    .Y(_06269_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[21] ));
 sg13g2_and4_1 _11201_ (.A(_06216_),
    .B(_06267_),
    .C(_06268_),
    .D(_06269_),
    .X(_06270_));
 sg13g2_nand4_1 _11202_ (.B(_06222_),
    .C(_06224_),
    .A(_06219_),
    .Y(_06271_),
    .D(_06270_));
 sg13g2_o21ai_1 _11203_ (.B1(_06231_),
    .Y(_06272_),
    .A1(_06266_),
    .A2(_06271_));
 sg13g2_nand3_1 _11204_ (.B(_06199_),
    .C(_06205_),
    .A(_06198_),
    .Y(_06273_));
 sg13g2_a22oi_1 _11205_ (.Y(_06274_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .B2(_00324_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .A1(_00326_));
 sg13g2_o21ai_1 _11206_ (.B1(_06274_),
    .Y(_06275_),
    .A1(_00319_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[24] ));
 sg13g2_nor4_1 _11207_ (.A(_06197_),
    .B(_06204_),
    .C(_06273_),
    .D(_06275_),
    .Y(_06276_));
 sg13g2_a21oi_1 _11208_ (.A1(_06272_),
    .A2(_06276_),
    .Y(_06277_),
    .B1(_06212_));
 sg13g2_nor2_1 _11209_ (.A(net1718),
    .B(net2769),
    .Y(_06278_));
 sg13g2_nor4_1 _11210_ (.A(_06169_),
    .B(_06171_),
    .C(_06176_),
    .D(_06278_),
    .Y(_06279_));
 sg13g2_nor4_1 _11211_ (.A(_06174_),
    .B(_06182_),
    .C(_06188_),
    .D(_06190_),
    .Y(_06280_));
 sg13g2_nand4_1 _11212_ (.B(_06187_),
    .C(_06279_),
    .A(_06175_),
    .Y(_06281_),
    .D(_06280_));
 sg13g2_o21ai_1 _11213_ (.B1(_06194_),
    .Y(_00023_),
    .A1(_06277_),
    .A2(net2959));
 sg13g2_nand2_2 _11214_ (.Y(_06282_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .B(_06129_));
 sg13g2_nor2_1 _11215_ (.A(net5072),
    .B(net5064),
    .Y(_06283_));
 sg13g2_o21ai_1 _11216_ (.B1(_06282_),
    .Y(_06284_),
    .A1(_06042_),
    .A2(_06283_));
 sg13g2_inv_1 _11217_ (.Y(_06285_),
    .A(_06284_));
 sg13g2_nand3_1 _11218_ (.B(net4278),
    .C(net410),
    .A(net334),
    .Y(_06286_));
 sg13g2_o21ai_1 _11219_ (.B1(_06286_),
    .Y(_00012_),
    .A1(net5124),
    .A2(_06285_));
 sg13g2_nor3_2 _11220_ (.A(\soc_inst.core_mem_addr[5] ),
    .B(\soc_inst.core_mem_addr[6] ),
    .C(\soc_inst.core_mem_addr[7] ),
    .Y(_06287_));
 sg13g2_and2_1 _11221_ (.A(net4740),
    .B(_06287_),
    .X(_06288_));
 sg13g2_nand2_2 _11222_ (.Y(_06289_),
    .A(net4740),
    .B(_06287_));
 sg13g2_nor2_2 _11223_ (.A(\soc_inst.core_mem_addr[1] ),
    .B(\soc_inst.core_mem_addr[0] ),
    .Y(_06290_));
 sg13g2_and2_1 _11224_ (.A(net4797),
    .B(_06290_),
    .X(_06291_));
 sg13g2_nand2_2 _11225_ (.Y(_06292_),
    .A(net4798),
    .B(_06290_));
 sg13g2_and2_1 _11226_ (.A(net4795),
    .B(_06290_),
    .X(_06293_));
 sg13g2_nand2_1 _11227_ (.Y(_06294_),
    .A(net4795),
    .B(_06290_));
 sg13g2_nor2_2 _11228_ (.A(_05485_),
    .B(net4655),
    .Y(_06295_));
 sg13g2_nand2_2 _11229_ (.Y(_06296_),
    .A(net4795),
    .B(net4657));
 sg13g2_nor2_1 _11230_ (.A(_06289_),
    .B(_06296_),
    .Y(_06297_));
 sg13g2_nand2_2 _11231_ (.Y(_06298_),
    .A(_06288_),
    .B(_06295_));
 sg13g2_and4_1 _11232_ (.A(\soc_inst.core_mem_addr[12] ),
    .B(\soc_inst.core_mem_addr[14] ),
    .C(_05881_),
    .D(_05884_),
    .X(_06299_));
 sg13g2_nand2_1 _11233_ (.Y(_06300_),
    .A(net4786),
    .B(_06299_));
 sg13g2_or3_1 _11234_ (.A(\soc_inst.spi_inst.busy ),
    .B(_06298_),
    .C(_06300_),
    .X(_06301_));
 sg13g2_nor4_1 _11235_ (.A(\soc_inst.core_mem_addr[15] ),
    .B(_05425_),
    .C(_05887_),
    .D(_05890_),
    .Y(_06302_));
 sg13g2_nand2_2 _11236_ (.Y(_06303_),
    .A(net4786),
    .B(_06302_));
 sg13g2_nor3_2 _11237_ (.A(\soc_inst.spi_inst.busy ),
    .B(_06298_),
    .C(_06303_),
    .Y(_06304_));
 sg13g2_nand2_1 _11238_ (.Y(_06305_),
    .A(net4785),
    .B(_05899_));
 sg13g2_or3_1 _11239_ (.A(\soc_inst.spi_inst.busy ),
    .B(_06298_),
    .C(_06305_),
    .X(_06306_));
 sg13g2_nor2_1 _11240_ (.A(net224),
    .B(net4012),
    .Y(_06307_));
 sg13g2_nor2_1 _11241_ (.A(net962),
    .B(net4062),
    .Y(_06308_));
 sg13g2_xor2_1 _11242_ (.B(\soc_inst.spi_inst.clk_counter[4] ),
    .A(_00221_),
    .X(_06309_));
 sg13g2_xnor2_1 _11243_ (.Y(_06310_),
    .A(\soc_inst.spi_inst.clk_counter[6] ),
    .B(\soc_inst.spi_inst.clock_divider[6] ));
 sg13g2_xor2_1 _11244_ (.B(\soc_inst.spi_inst.clk_counter[3] ),
    .A(_00220_),
    .X(_06311_));
 sg13g2_xor2_1 _11245_ (.B(\soc_inst.spi_inst.clk_counter[1] ),
    .A(_00218_),
    .X(_06312_));
 sg13g2_o21ai_1 _11246_ (.B1(_06312_),
    .Y(_06313_),
    .A1(_00217_),
    .A2(\soc_inst.spi_inst.clk_counter[0] ));
 sg13g2_xnor2_1 _11247_ (.Y(_06314_),
    .A(\soc_inst.spi_inst.clk_counter[7] ),
    .B(\soc_inst.spi_inst.clock_divider[7] ));
 sg13g2_xor2_1 _11248_ (.B(\soc_inst.spi_inst.clock_divider[5] ),
    .A(\soc_inst.spi_inst.clk_counter[5] ),
    .X(_06315_));
 sg13g2_xor2_1 _11249_ (.B(\soc_inst.spi_inst.clk_counter[2] ),
    .A(_00219_),
    .X(_06316_));
 sg13g2_xor2_1 _11250_ (.B(\soc_inst.spi_inst.clk_counter[0] ),
    .A(_00217_),
    .X(_06317_));
 sg13g2_nand3_1 _11251_ (.B(_06312_),
    .C(_06316_),
    .A(_06309_),
    .Y(_06318_));
 sg13g2_nand4_1 _11252_ (.B(_06311_),
    .C(_06314_),
    .A(_06310_),
    .Y(_06319_),
    .D(_06317_));
 sg13g2_nor3_1 _11253_ (.A(_06315_),
    .B(_06318_),
    .C(_06319_),
    .Y(_06320_));
 sg13g2_nand2_1 _11254_ (.Y(_06321_),
    .A(\soc_inst.spi_inst.spi_clk_en ),
    .B(_06320_));
 sg13g2_inv_1 _11255_ (.Y(_06322_),
    .A(_06321_));
 sg13g2_nand3_1 _11256_ (.B(\soc_inst.spi_inst.spi_sclk ),
    .C(_06322_),
    .A(\soc_inst.spi_inst.cpol ),
    .Y(_06323_));
 sg13g2_or2_1 _11257_ (.X(_06324_),
    .B(_06321_),
    .A(net2277));
 sg13g2_o21ai_1 _11258_ (.B1(_06323_),
    .Y(_06325_),
    .A1(\soc_inst.spi_inst.cpol ),
    .A2(_06324_));
 sg13g2_nor2_1 _11259_ (.A(\soc_inst.spi_inst.cpha ),
    .B(_06325_),
    .Y(_06326_));
 sg13g2_a21oi_1 _11260_ (.A1(\soc_inst.spi_inst.spi_sclk ),
    .A2(_06322_),
    .Y(_06327_),
    .B1(\soc_inst.spi_inst.cpol ));
 sg13g2_a21o_1 _11261_ (.A2(_06324_),
    .A1(\soc_inst.spi_inst.cpol ),
    .B1(_06327_),
    .X(_06328_));
 sg13g2_and2_1 _11262_ (.A(\soc_inst.spi_inst.cpha ),
    .B(_06328_),
    .X(_06329_));
 sg13g2_nor3_1 _11263_ (.A(net4716),
    .B(_06326_),
    .C(_06329_),
    .Y(_06330_));
 sg13g2_nor3_2 _11264_ (.A(net4716),
    .B(_06326_),
    .C(_06329_),
    .Y(_06331_));
 sg13g2_nor3_1 _11265_ (.A(net4717),
    .B(_06326_),
    .C(_06329_),
    .Y(_06332_));
 sg13g2_nor3_1 _11266_ (.A(_06307_),
    .B(_06308_),
    .C(net3871),
    .Y(_00134_));
 sg13g2_nand2_1 _11267_ (.Y(_06333_),
    .A(_05551_),
    .B(net4062));
 sg13g2_o21ai_1 _11268_ (.B1(_06333_),
    .Y(_06334_),
    .A1(\soc_inst.core_mem_wdata[25] ),
    .A2(net4009));
 sg13g2_nand2_1 _11269_ (.Y(_06335_),
    .A(net224),
    .B(net3871));
 sg13g2_o21ai_1 _11270_ (.B1(_06335_),
    .Y(_00145_),
    .A1(net3871),
    .A2(_06334_));
 sg13g2_a221oi_1 _11271_ (.B2(\soc_inst.core_mem_wdata[26] ),
    .C1(net3879),
    .B1(net4012),
    .A1(net273),
    .Y(_06336_),
    .A2(net4062));
 sg13g2_a21oi_1 _11272_ (.A1(_05551_),
    .A2(net3871),
    .Y(_00156_),
    .B1(_06336_));
 sg13g2_or2_1 _11273_ (.X(_06337_),
    .B(net4012),
    .A(net238));
 sg13g2_o21ai_1 _11274_ (.B1(_06337_),
    .Y(_06338_),
    .A1(\soc_inst.core_mem_wdata[27] ),
    .A2(net4009));
 sg13g2_nand2_1 _11275_ (.Y(_06339_),
    .A(net273),
    .B(net3872));
 sg13g2_o21ai_1 _11276_ (.B1(_06339_),
    .Y(_00159_),
    .A1(net3872),
    .A2(_06338_));
 sg13g2_nand2_1 _11277_ (.Y(_06340_),
    .A(_05552_),
    .B(net4061));
 sg13g2_o21ai_1 _11278_ (.B1(_06340_),
    .Y(_06341_),
    .A1(\soc_inst.core_mem_wdata[28] ),
    .A2(net4009));
 sg13g2_nand2_1 _11279_ (.Y(_06342_),
    .A(net238),
    .B(net3871));
 sg13g2_o21ai_1 _11280_ (.B1(_06342_),
    .Y(_00160_),
    .A1(net3872),
    .A2(_06341_));
 sg13g2_a221oi_1 _11281_ (.B2(\soc_inst.core_mem_wdata[29] ),
    .C1(net3879),
    .B1(net4012),
    .A1(net243),
    .Y(_06343_),
    .A2(net4061));
 sg13g2_a21oi_1 _11282_ (.A1(_05552_),
    .A2(net3871),
    .Y(_00161_),
    .B1(_06343_));
 sg13g2_or2_1 _11283_ (.X(_06344_),
    .B(net4011),
    .A(net170));
 sg13g2_o21ai_1 _11284_ (.B1(_06344_),
    .Y(_06345_),
    .A1(\soc_inst.core_mem_wdata[30] ),
    .A2(net4009));
 sg13g2_nand2_1 _11285_ (.Y(_06346_),
    .A(net243),
    .B(net3871));
 sg13g2_o21ai_1 _11286_ (.B1(_06346_),
    .Y(_00162_),
    .A1(net3870),
    .A2(_06345_));
 sg13g2_nand2_1 _11287_ (.Y(_06347_),
    .A(_05553_),
    .B(net4061));
 sg13g2_o21ai_1 _11288_ (.B1(_06347_),
    .Y(_06348_),
    .A1(\soc_inst.core_mem_wdata[31] ),
    .A2(net4009));
 sg13g2_nand2_1 _11289_ (.Y(_06349_),
    .A(net170),
    .B(net3870));
 sg13g2_o21ai_1 _11290_ (.B1(_06349_),
    .Y(_00163_),
    .A1(net3870),
    .A2(_06348_));
 sg13g2_a221oi_1 _11291_ (.B2(\soc_inst.core_mem_wdata[16] ),
    .C1(net3879),
    .B1(net4011),
    .A1(net301),
    .Y(_06350_),
    .A2(net4061));
 sg13g2_a21oi_1 _11292_ (.A1(_05553_),
    .A2(net3870),
    .Y(_00164_),
    .B1(_06350_));
 sg13g2_a221oi_1 _11293_ (.B2(\soc_inst.core_mem_wdata[17] ),
    .C1(net3879),
    .B1(net4011),
    .A1(\soc_inst.spi_inst.tx_shift_reg[9] ),
    .Y(_06351_),
    .A2(net4061));
 sg13g2_a21oi_1 _11294_ (.A1(_05554_),
    .A2(net3870),
    .Y(_00165_),
    .B1(_06351_));
 sg13g2_a221oi_1 _11295_ (.B2(\soc_inst.core_mem_wdata[18] ),
    .C1(net3879),
    .B1(net4011),
    .A1(net215),
    .Y(_06352_),
    .A2(net4061));
 sg13g2_a21oi_1 _11296_ (.A1(_05555_),
    .A2(net3870),
    .Y(_00135_),
    .B1(_06352_));
 sg13g2_or2_1 _11297_ (.X(_06353_),
    .B(net4011),
    .A(net149));
 sg13g2_o21ai_1 _11298_ (.B1(_06353_),
    .Y(_06354_),
    .A1(\soc_inst.core_mem_wdata[19] ),
    .A2(net4009));
 sg13g2_nand2_1 _11299_ (.Y(_06355_),
    .A(net215),
    .B(net3869));
 sg13g2_o21ai_1 _11300_ (.B1(_06355_),
    .Y(_00136_),
    .A1(net3869),
    .A2(_06354_));
 sg13g2_or2_1 _11301_ (.X(_06356_),
    .B(net4011),
    .A(\soc_inst.spi_inst.tx_shift_reg[12] ));
 sg13g2_o21ai_1 _11302_ (.B1(_06356_),
    .Y(_06357_),
    .A1(\soc_inst.core_mem_wdata[20] ),
    .A2(net4009));
 sg13g2_nand2_1 _11303_ (.Y(_06358_),
    .A(net149),
    .B(net3869));
 sg13g2_o21ai_1 _11304_ (.B1(_06358_),
    .Y(_00137_),
    .A1(net3869),
    .A2(_06357_));
 sg13g2_nand2_1 _11305_ (.Y(_06359_),
    .A(_05556_),
    .B(net4061));
 sg13g2_o21ai_1 _11306_ (.B1(_06359_),
    .Y(_06360_),
    .A1(\soc_inst.core_mem_wdata[21] ),
    .A2(net4010));
 sg13g2_nand2_1 _11307_ (.Y(_06361_),
    .A(net438),
    .B(net3869));
 sg13g2_o21ai_1 _11308_ (.B1(_06361_),
    .Y(_00138_),
    .A1(net3873),
    .A2(_06360_));
 sg13g2_a221oi_1 _11309_ (.B2(\soc_inst.core_mem_wdata[22] ),
    .C1(net3879),
    .B1(net4011),
    .A1(net269),
    .Y(_06362_),
    .A2(net4061));
 sg13g2_a21oi_1 _11310_ (.A1(_05556_),
    .A2(net3869),
    .Y(_00139_),
    .B1(_06362_));
 sg13g2_or2_1 _11311_ (.X(_06363_),
    .B(net4011),
    .A(net118));
 sg13g2_o21ai_1 _11312_ (.B1(_06363_),
    .Y(_06364_),
    .A1(\soc_inst.core_mem_wdata[23] ),
    .A2(net4009));
 sg13g2_nand2_1 _11313_ (.Y(_06365_),
    .A(net269),
    .B(net3869));
 sg13g2_o21ai_1 _11314_ (.B1(_06365_),
    .Y(_00140_),
    .A1(net3871),
    .A2(_06364_));
 sg13g2_or2_1 _11315_ (.X(_06366_),
    .B(net4014),
    .A(\soc_inst.spi_inst.tx_shift_reg[16] ));
 sg13g2_o21ai_1 _11316_ (.B1(_06366_),
    .Y(_06367_),
    .A1(net5027),
    .A2(net4010));
 sg13g2_nand2_1 _11317_ (.Y(_06368_),
    .A(net118),
    .B(net3873));
 sg13g2_o21ai_1 _11318_ (.B1(_06368_),
    .Y(_00141_),
    .A1(net3874),
    .A2(_06367_));
 sg13g2_nand2_1 _11319_ (.Y(_06369_),
    .A(_05557_),
    .B(net4065));
 sg13g2_o21ai_1 _11320_ (.B1(_06369_),
    .Y(_06370_),
    .A1(net5024),
    .A2(net4010));
 sg13g2_nand2_1 _11321_ (.Y(_06371_),
    .A(net187),
    .B(net3874));
 sg13g2_o21ai_1 _11322_ (.B1(_06371_),
    .Y(_00142_),
    .A1(net3874),
    .A2(_06370_));
 sg13g2_a221oi_1 _11323_ (.B2(net5023),
    .C1(_06331_),
    .B1(net4014),
    .A1(net165),
    .Y(_06372_),
    .A2(net4065));
 sg13g2_a21oi_1 _11324_ (.A1(_05557_),
    .A2(net3874),
    .Y(_00143_),
    .B1(_06372_));
 sg13g2_or2_1 _11325_ (.X(_06373_),
    .B(net4014),
    .A(net113));
 sg13g2_o21ai_1 _11326_ (.B1(_06373_),
    .Y(_06374_),
    .A1(net5022),
    .A2(net4010));
 sg13g2_nand2_1 _11327_ (.Y(_06375_),
    .A(net165),
    .B(net3874));
 sg13g2_o21ai_1 _11328_ (.B1(_06375_),
    .Y(_00144_),
    .A1(net3877),
    .A2(_06374_));
 sg13g2_or2_1 _11329_ (.X(_06376_),
    .B(net4013),
    .A(\soc_inst.spi_inst.tx_shift_reg[20] ));
 sg13g2_o21ai_1 _11330_ (.B1(_06376_),
    .Y(_06377_),
    .A1(net5021),
    .A2(net4010));
 sg13g2_nand2_1 _11331_ (.Y(_06378_),
    .A(net113),
    .B(net3876));
 sg13g2_o21ai_1 _11332_ (.B1(_06378_),
    .Y(_00146_),
    .A1(net3876),
    .A2(_06377_));
 sg13g2_nand2_1 _11333_ (.Y(_06379_),
    .A(_05558_),
    .B(net4063));
 sg13g2_o21ai_1 _11334_ (.B1(_06379_),
    .Y(_06380_),
    .A1(net5020),
    .A2(net4010));
 sg13g2_nand2_1 _11335_ (.Y(_06381_),
    .A(net137),
    .B(net3876));
 sg13g2_o21ai_1 _11336_ (.B1(_06381_),
    .Y(_00147_),
    .A1(net3876),
    .A2(_06380_));
 sg13g2_a221oi_1 _11337_ (.B2(net5019),
    .C1(net3878),
    .B1(net4013),
    .A1(net329),
    .Y(_06382_),
    .A2(net4063));
 sg13g2_a21oi_1 _11338_ (.A1(_05558_),
    .A2(net3876),
    .Y(_00148_),
    .B1(_06382_));
 sg13g2_a221oi_1 _11339_ (.B2(net5018),
    .C1(net3878),
    .B1(net4013),
    .A1(net307),
    .Y(_06383_),
    .A2(net4063));
 sg13g2_a21oi_1 _11340_ (.A1(_05559_),
    .A2(net3876),
    .Y(_00149_),
    .B1(_06383_));
 sg13g2_a221oi_1 _11341_ (.B2(net5048),
    .C1(net3878),
    .B1(net4013),
    .A1(\soc_inst.spi_inst.tx_shift_reg[24] ),
    .Y(_06384_),
    .A2(net4063));
 sg13g2_a21oi_1 _11342_ (.A1(_05560_),
    .A2(net3876),
    .Y(_00150_),
    .B1(_06384_));
 sg13g2_a221oi_1 _11343_ (.B2(net5046),
    .C1(net3878),
    .B1(net4014),
    .A1(\soc_inst.spi_inst.tx_shift_reg[25] ),
    .Y(_06385_),
    .A2(net4064));
 sg13g2_a21oi_1 _11344_ (.A1(_05561_),
    .A2(net3875),
    .Y(_00151_),
    .B1(_06385_));
 sg13g2_a221oi_1 _11345_ (.B2(net5042),
    .C1(net3879),
    .B1(net4014),
    .A1(net232),
    .Y(_06386_),
    .A2(net4064));
 sg13g2_a21oi_1 _11346_ (.A1(_05562_),
    .A2(net3875),
    .Y(_00152_),
    .B1(_06386_));
 sg13g2_nand2_1 _11347_ (.Y(_06387_),
    .A(_05563_),
    .B(net4064));
 sg13g2_o21ai_1 _11348_ (.B1(_06387_),
    .Y(_06388_),
    .A1(net5039),
    .A2(net4010));
 sg13g2_nand2_1 _11349_ (.Y(_06389_),
    .A(net232),
    .B(net3875));
 sg13g2_o21ai_1 _11350_ (.B1(_06389_),
    .Y(_00153_),
    .A1(net3875),
    .A2(_06388_));
 sg13g2_a221oi_1 _11351_ (.B2(net5036),
    .C1(net3878),
    .B1(net4013),
    .A1(net339),
    .Y(_06390_),
    .A2(net4063));
 sg13g2_a21oi_1 _11352_ (.A1(_05563_),
    .A2(net3875),
    .Y(_00154_),
    .B1(_06390_));
 sg13g2_a221oi_1 _11353_ (.B2(net5033),
    .C1(net3878),
    .B1(net4013),
    .A1(\soc_inst.spi_inst.tx_shift_reg[29] ),
    .Y(_06391_),
    .A2(net4063));
 sg13g2_a21oi_1 _11354_ (.A1(_05564_),
    .A2(net3875),
    .Y(_00155_),
    .B1(_06391_));
 sg13g2_a221oi_1 _11355_ (.B2(net5031),
    .C1(net3878),
    .B1(net4013),
    .A1(\soc_inst.spi_inst.tx_shift_reg[30] ),
    .Y(_06392_),
    .A2(net4063));
 sg13g2_a21oi_1 _11356_ (.A1(_05565_),
    .A2(net3875),
    .Y(_00157_),
    .B1(_06392_));
 sg13g2_a221oi_1 _11357_ (.B2(net5028),
    .C1(net3878),
    .B1(net4013),
    .A1(\soc_inst.spi_inst.tx_shift_reg[31] ),
    .Y(_06393_),
    .A2(net4063));
 sg13g2_a21oi_1 _11358_ (.A1(_05566_),
    .A2(net3875),
    .Y(_00158_),
    .B1(_06393_));
 sg13g2_nand2b_2 _11359_ (.Y(_06394_),
    .B(\soc_inst.spi_inst.spi_clk_en ),
    .A_N(_06320_));
 sg13g2_inv_2 _11360_ (.Y(_06395_),
    .A(_06394_));
 sg13g2_nor2_1 _11361_ (.A(net490),
    .B(_06394_),
    .Y(_00124_));
 sg13g2_o21ai_1 _11362_ (.B1(_06395_),
    .Y(_06396_),
    .A1(net490),
    .A2(net494));
 sg13g2_a21oi_1 _11363_ (.A1(net490),
    .A2(net494),
    .Y(_00125_),
    .B1(_06396_));
 sg13g2_and3_1 _11364_ (.X(_06397_),
    .A(net490),
    .B(net494),
    .C(net584));
 sg13g2_a21oi_1 _11365_ (.A1(net490),
    .A2(net494),
    .Y(_06398_),
    .B1(net584));
 sg13g2_nor3_1 _11366_ (.A(_06394_),
    .B(_06397_),
    .C(_06398_),
    .Y(_00126_));
 sg13g2_and2_1 _11367_ (.A(net1918),
    .B(_06397_),
    .X(_06399_));
 sg13g2_nor2_1 _11368_ (.A(net1918),
    .B(_06397_),
    .Y(_06400_));
 sg13g2_nor3_1 _11369_ (.A(_06394_),
    .B(_06399_),
    .C(_06400_),
    .Y(_00127_));
 sg13g2_and2_1 _11370_ (.A(net1935),
    .B(_06399_),
    .X(_06401_));
 sg13g2_nor2_1 _11371_ (.A(net1935),
    .B(_06399_),
    .Y(_06402_));
 sg13g2_nor3_1 _11372_ (.A(_06394_),
    .B(_06401_),
    .C(_06402_),
    .Y(_00128_));
 sg13g2_nor2_1 _11373_ (.A(net2378),
    .B(_06401_),
    .Y(_06403_));
 sg13g2_and2_1 _11374_ (.A(net2378),
    .B(_06401_),
    .X(_06404_));
 sg13g2_nor3_1 _11375_ (.A(_06394_),
    .B(_06403_),
    .C(_06404_),
    .Y(_00129_));
 sg13g2_and2_1 _11376_ (.A(net1993),
    .B(_06404_),
    .X(_06405_));
 sg13g2_nor2_1 _11377_ (.A(net1993),
    .B(_06404_),
    .Y(_06406_));
 sg13g2_nor3_1 _11378_ (.A(_06394_),
    .B(_06405_),
    .C(net1994),
    .Y(_00130_));
 sg13g2_o21ai_1 _11379_ (.B1(_06395_),
    .Y(_06407_),
    .A1(net502),
    .A2(_06405_));
 sg13g2_a21oi_1 _11380_ (.A1(net502),
    .A2(_06405_),
    .Y(_00131_),
    .B1(_06407_));
 sg13g2_nand2_1 _11381_ (.Y(_06408_),
    .A(net2277),
    .B(_06395_));
 sg13g2_nand2b_1 _11382_ (.Y(_06409_),
    .B(\soc_inst.spi_inst.cpol ),
    .A_N(\soc_inst.spi_inst.spi_clk_en ));
 sg13g2_nand3_1 _11383_ (.B(net2278),
    .C(_06409_),
    .A(_06324_),
    .Y(_00132_));
 sg13g2_nor3_1 _11384_ (.A(\soc_inst.core_mem_addr[1] ),
    .B(\soc_inst.core_mem_addr[0] ),
    .C(net4796),
    .Y(_06410_));
 sg13g2_and2_1 _11385_ (.A(_05484_),
    .B(net4714),
    .X(_06411_));
 sg13g2_nand2_1 _11386_ (.Y(_06412_),
    .A(_05484_),
    .B(net4713));
 sg13g2_nand2_1 _11387_ (.Y(_06413_),
    .A(net4785),
    .B(_05902_));
 sg13g2_nor2_2 _11388_ (.A(net4651),
    .B(_06413_),
    .Y(_06414_));
 sg13g2_a21oi_1 _11389_ (.A1(net5045),
    .A2(_06414_),
    .Y(_06415_),
    .B1(net824));
 sg13g2_nor2b_1 _11390_ (.A(net5117),
    .B_N(net5116),
    .Y(_06416_));
 sg13g2_nand2b_1 _11391_ (.Y(_06417_),
    .B(net5116),
    .A_N(net5117));
 sg13g2_nand2_2 _11392_ (.Y(_06418_),
    .A(net5120),
    .B(_05471_));
 sg13g2_xnor2_1 _11393_ (.Y(_06419_),
    .A(_00222_),
    .B(\soc_inst.i2c_inst.clk_cnt[0] ));
 sg13g2_xnor2_1 _11394_ (.Y(_06420_),
    .A(\soc_inst.i2c_inst.prescale_reg[6] ),
    .B(\soc_inst.i2c_inst.clk_cnt[6] ));
 sg13g2_xnor2_1 _11395_ (.Y(_06421_),
    .A(_00227_),
    .B(\soc_inst.i2c_inst.clk_cnt[7] ));
 sg13g2_xnor2_1 _11396_ (.Y(_06422_),
    .A(_00223_),
    .B(\soc_inst.i2c_inst.clk_cnt[1] ));
 sg13g2_xor2_1 _11397_ (.B(\soc_inst.i2c_inst.clk_cnt[5] ),
    .A(\soc_inst.i2c_inst.prescale_reg[5] ),
    .X(_06423_));
 sg13g2_xnor2_1 _11398_ (.Y(_06424_),
    .A(_00224_),
    .B(\soc_inst.i2c_inst.clk_cnt[2] ));
 sg13g2_xnor2_1 _11399_ (.Y(_06425_),
    .A(_00226_),
    .B(\soc_inst.i2c_inst.clk_cnt[4] ));
 sg13g2_xnor2_1 _11400_ (.Y(_06426_),
    .A(_00225_),
    .B(\soc_inst.i2c_inst.clk_cnt[3] ));
 sg13g2_nor4_1 _11401_ (.A(_06419_),
    .B(_06421_),
    .C(_06423_),
    .D(_06425_),
    .Y(_06427_));
 sg13g2_nor3_1 _11402_ (.A(_06422_),
    .B(_06424_),
    .C(_06426_),
    .Y(_06428_));
 sg13g2_nand3_1 _11403_ (.B(_06427_),
    .C(_06428_),
    .A(_06420_),
    .Y(_06429_));
 sg13g2_inv_1 _11404_ (.Y(_06430_),
    .A(net4276));
 sg13g2_nor3_1 _11405_ (.A(_06417_),
    .B(_06418_),
    .C(net4274),
    .Y(_06431_));
 sg13g2_nor2_1 _11406_ (.A(_06415_),
    .B(_06431_),
    .Y(_00086_));
 sg13g2_nor2_1 _11407_ (.A(net4798),
    .B(_06294_),
    .Y(_06432_));
 sg13g2_nand2_2 _11408_ (.Y(_06433_),
    .A(_05484_),
    .B(_06293_));
 sg13g2_nor2_1 _11409_ (.A(_06413_),
    .B(net4270),
    .Y(_06434_));
 sg13g2_nand3_1 _11410_ (.B(_05902_),
    .C(net4272),
    .A(net4785),
    .Y(_06435_));
 sg13g2_nand2_1 _11411_ (.Y(_06436_),
    .A(net81),
    .B(net4060));
 sg13g2_a21oi_1 _11412_ (.A1(net5048),
    .A2(_06414_),
    .Y(_06437_),
    .B1(_06436_));
 sg13g2_nand2b_2 _11413_ (.Y(_06438_),
    .B(\soc_inst.i2c_inst.state[1] ),
    .A_N(\soc_inst.i2c_inst.state[0] ));
 sg13g2_nor2b_2 _11414_ (.A(net5116),
    .B_N(net5117),
    .Y(_06439_));
 sg13g2_nand2b_2 _11415_ (.Y(_06440_),
    .B(net5117),
    .A_N(net5115));
 sg13g2_nor2_1 _11416_ (.A(net5115),
    .B(_06438_),
    .Y(_06441_));
 sg13g2_or2_1 _11417_ (.X(_06442_),
    .B(_06438_),
    .A(net5115));
 sg13g2_nor2_1 _11418_ (.A(_06438_),
    .B(_06440_),
    .Y(_06443_));
 sg13g2_nand2_1 _11419_ (.Y(_06444_),
    .A(net5119),
    .B(_06441_));
 sg13g2_nor2_1 _11420_ (.A(net4276),
    .B(_06444_),
    .Y(_06445_));
 sg13g2_or2_1 _11421_ (.X(_00087_),
    .B(net4205),
    .A(_06437_));
 sg13g2_or2_1 _11422_ (.X(_06446_),
    .B(net4060),
    .A(net5048));
 sg13g2_o21ai_1 _11423_ (.B1(_06446_),
    .Y(_06447_),
    .A1(\soc_inst.i2c_inst.data_reg[0] ),
    .A2(net4008));
 sg13g2_nand2_1 _11424_ (.Y(_06448_),
    .A(net669),
    .B(net4204));
 sg13g2_o21ai_1 _11425_ (.B1(_06448_),
    .Y(_00078_),
    .A1(net4204),
    .A2(_06447_));
 sg13g2_nor2_1 _11426_ (.A(net5046),
    .B(net4060),
    .Y(_06449_));
 sg13g2_inv_1 _11427_ (.Y(_06450_),
    .A(_06449_));
 sg13g2_o21ai_1 _11428_ (.B1(_06450_),
    .Y(_06451_),
    .A1(\soc_inst.i2c_inst.data_reg[1] ),
    .A2(net4007));
 sg13g2_nand2_1 _11429_ (.Y(_06452_),
    .A(net545),
    .B(net4203));
 sg13g2_o21ai_1 _11430_ (.B1(_06452_),
    .Y(_00079_),
    .A1(net4203),
    .A2(_06451_));
 sg13g2_nor2_1 _11431_ (.A(\soc_inst.i2c_inst.data_reg[2] ),
    .B(net4007),
    .Y(_06453_));
 sg13g2_nor2_1 _11432_ (.A(net5041),
    .B(net4060),
    .Y(_06454_));
 sg13g2_nor3_1 _11433_ (.A(net4203),
    .B(_06453_),
    .C(_06454_),
    .Y(_06455_));
 sg13g2_a21o_1 _11434_ (.A2(net4203),
    .A1(net1523),
    .B1(_06455_),
    .X(_00080_));
 sg13g2_or2_1 _11435_ (.X(_06456_),
    .B(net4060),
    .A(net5038));
 sg13g2_o21ai_1 _11436_ (.B1(_06456_),
    .Y(_06457_),
    .A1(\soc_inst.i2c_inst.data_reg[3] ),
    .A2(net4007));
 sg13g2_nand2_1 _11437_ (.Y(_06458_),
    .A(net652),
    .B(net4203));
 sg13g2_o21ai_1 _11438_ (.B1(_06458_),
    .Y(_00081_),
    .A1(net4203),
    .A2(_06457_));
 sg13g2_or2_1 _11439_ (.X(_06459_),
    .B(net4060),
    .A(net5036));
 sg13g2_o21ai_1 _11440_ (.B1(_06459_),
    .Y(_06460_),
    .A1(\soc_inst.i2c_inst.data_reg[4] ),
    .A2(net4006));
 sg13g2_nand2_1 _11441_ (.Y(_06461_),
    .A(net492),
    .B(net4205));
 sg13g2_o21ai_1 _11442_ (.B1(_06461_),
    .Y(_00082_),
    .A1(net4205),
    .A2(_06460_));
 sg13g2_nor2_1 _11443_ (.A(net5034),
    .B(net4060),
    .Y(_06462_));
 sg13g2_inv_1 _11444_ (.Y(_06463_),
    .A(_06462_));
 sg13g2_o21ai_1 _11445_ (.B1(_06463_),
    .Y(_06464_),
    .A1(\soc_inst.i2c_inst.data_reg[5] ),
    .A2(net4006));
 sg13g2_nand2_1 _11446_ (.Y(_06465_),
    .A(net536),
    .B(net4203));
 sg13g2_o21ai_1 _11447_ (.B1(_06465_),
    .Y(_00083_),
    .A1(net4203),
    .A2(_06464_));
 sg13g2_nor2_1 _11448_ (.A(\soc_inst.i2c_inst.data_reg[6] ),
    .B(net4006),
    .Y(_06466_));
 sg13g2_nor2_1 _11449_ (.A(net5031),
    .B(net4060),
    .Y(_06467_));
 sg13g2_nor3_1 _11450_ (.A(net4205),
    .B(_06466_),
    .C(_06467_),
    .Y(_06468_));
 sg13g2_a21o_1 _11451_ (.A2(net4205),
    .A1(net1692),
    .B1(_06468_),
    .X(_00084_));
 sg13g2_nor2_1 _11452_ (.A(net1790),
    .B(net4008),
    .Y(_06469_));
 sg13g2_nor2_1 _11453_ (.A(net5028),
    .B(_06435_),
    .Y(_06470_));
 sg13g2_nor3_1 _11454_ (.A(net4204),
    .B(_06469_),
    .C(_06470_),
    .Y(_06471_));
 sg13g2_a21o_1 _11455_ (.A2(net4204),
    .A1(net1183),
    .B1(_06471_),
    .X(_00085_));
 sg13g2_nand2_1 _11456_ (.Y(_06472_),
    .A(\soc_inst.i2c_ena ),
    .B(net4276));
 sg13g2_nor2_1 _11457_ (.A(net315),
    .B(net4202),
    .Y(_00070_));
 sg13g2_xnor2_1 _11458_ (.Y(_06473_),
    .A(net315),
    .B(net2461));
 sg13g2_nor2_1 _11459_ (.A(net4202),
    .B(_06473_),
    .Y(_00071_));
 sg13g2_and3_1 _11460_ (.X(_06474_),
    .A(net315),
    .B(\soc_inst.i2c_inst.clk_cnt[1] ),
    .C(net710));
 sg13g2_a21oi_1 _11461_ (.A1(net315),
    .A2(\soc_inst.i2c_inst.clk_cnt[1] ),
    .Y(_06475_),
    .B1(net710));
 sg13g2_nor3_1 _11462_ (.A(net4202),
    .B(_06474_),
    .C(net711),
    .Y(_00072_));
 sg13g2_and2_1 _11463_ (.A(net1556),
    .B(_06474_),
    .X(_06476_));
 sg13g2_nor2_1 _11464_ (.A(net1556),
    .B(_06474_),
    .Y(_06477_));
 sg13g2_nor3_1 _11465_ (.A(net4202),
    .B(_06476_),
    .C(net1557),
    .Y(_00073_));
 sg13g2_and2_1 _11466_ (.A(net1701),
    .B(_06476_),
    .X(_06478_));
 sg13g2_nor2_1 _11467_ (.A(net1701),
    .B(_06476_),
    .Y(_06479_));
 sg13g2_nor3_1 _11468_ (.A(net4202),
    .B(_06478_),
    .C(net1702),
    .Y(_00074_));
 sg13g2_and2_1 _11469_ (.A(net2177),
    .B(_06478_),
    .X(_06480_));
 sg13g2_nor2_1 _11470_ (.A(net2177),
    .B(_06478_),
    .Y(_06481_));
 sg13g2_nor3_1 _11471_ (.A(net4202),
    .B(_06480_),
    .C(_06481_),
    .Y(_00075_));
 sg13g2_and2_1 _11472_ (.A(net2274),
    .B(_06480_),
    .X(_06482_));
 sg13g2_nor2_1 _11473_ (.A(net2274),
    .B(_06480_),
    .Y(_06483_));
 sg13g2_nor3_1 _11474_ (.A(net4202),
    .B(_06482_),
    .C(_06483_),
    .Y(_00076_));
 sg13g2_a21oi_1 _11475_ (.A1(net2604),
    .A2(_06482_),
    .Y(_06484_),
    .B1(_06472_));
 sg13g2_o21ai_1 _11476_ (.B1(_06484_),
    .Y(_06485_),
    .A1(net2604),
    .A2(_06482_));
 sg13g2_inv_1 _11477_ (.Y(_00077_),
    .A(_06485_));
 sg13g2_nor2_1 _11478_ (.A(_00251_),
    .B(\soc_inst.pwm_inst.channel_counter[1][5] ),
    .Y(_06486_));
 sg13g2_nand2_1 _11479_ (.Y(_06487_),
    .A(_00251_),
    .B(\soc_inst.pwm_inst.channel_counter[1][5] ));
 sg13g2_nor2_1 _11480_ (.A(_00247_),
    .B(\soc_inst.pwm_inst.channel_counter[1][1] ),
    .Y(_06488_));
 sg13g2_nor2_1 _11481_ (.A(_00246_),
    .B(\soc_inst.pwm_inst.channel_counter[1][0] ),
    .Y(_06489_));
 sg13g2_a22oi_1 _11482_ (.Y(_06490_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][1] ),
    .B2(_00247_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][2] ),
    .A1(_00248_));
 sg13g2_o21ai_1 _11483_ (.B1(_06490_),
    .Y(_06491_),
    .A1(_06488_),
    .A2(_06489_));
 sg13g2_nor2_1 _11484_ (.A(_00249_),
    .B(\soc_inst.pwm_inst.channel_counter[1][3] ),
    .Y(_06492_));
 sg13g2_o21ai_1 _11485_ (.B1(_06491_),
    .Y(_06493_),
    .A1(_00248_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][2] ));
 sg13g2_a22oi_1 _11486_ (.Y(_06494_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][3] ),
    .B2(_00249_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][4] ),
    .A1(_00250_));
 sg13g2_o21ai_1 _11487_ (.B1(_06494_),
    .Y(_06495_),
    .A1(_06492_),
    .A2(_06493_));
 sg13g2_o21ai_1 _11488_ (.B1(_06495_),
    .Y(_06496_),
    .A1(_00250_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][4] ));
 sg13g2_a21oi_1 _11489_ (.A1(_06487_),
    .A2(_06496_),
    .Y(_06497_),
    .B1(_06486_));
 sg13g2_o21ai_1 _11490_ (.B1(_06497_),
    .Y(_06498_),
    .A1(_00252_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][6] ));
 sg13g2_a22oi_1 _11491_ (.Y(_06499_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][6] ),
    .B2(_00252_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][7] ),
    .A1(_00253_));
 sg13g2_or2_1 _11492_ (.X(_06500_),
    .B(\soc_inst.pwm_inst.channel_counter[1][8] ),
    .A(_00254_));
 sg13g2_o21ai_1 _11493_ (.B1(_06500_),
    .Y(_06501_),
    .A1(_00253_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][7] ));
 sg13g2_a21oi_1 _11494_ (.A1(_06498_),
    .A2(_06499_),
    .Y(_06502_),
    .B1(_06501_));
 sg13g2_a221oi_1 _11495_ (.B2(_00254_),
    .C1(_06502_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][8] ),
    .A1(_00255_),
    .Y(_06503_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][9] ));
 sg13g2_nor2_1 _11496_ (.A(_00256_),
    .B(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .Y(_06504_));
 sg13g2_nor2_1 _11497_ (.A(_00255_),
    .B(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .Y(_06505_));
 sg13g2_nor2_1 _11498_ (.A(_00257_),
    .B(\soc_inst.pwm_inst.channel_counter[1][11] ),
    .Y(_06506_));
 sg13g2_nor4_1 _11499_ (.A(_06503_),
    .B(_06504_),
    .C(_06505_),
    .D(_06506_),
    .Y(_06507_));
 sg13g2_a221oi_1 _11500_ (.B2(_00256_),
    .C1(_06507_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .A1(_00257_),
    .Y(_06508_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][11] ));
 sg13g2_a22oi_1 _11501_ (.Y(_06509_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][12] ),
    .B2(_00258_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][13] ),
    .A1(_00259_));
 sg13g2_nor2_1 _11502_ (.A(_00261_),
    .B(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .Y(_06510_));
 sg13g2_a21oi_1 _11503_ (.A1(_05404_),
    .A2(_05569_),
    .Y(_06511_),
    .B1(_06510_));
 sg13g2_nand3_1 _11504_ (.B(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .C(_06506_),
    .A(_00256_),
    .Y(_06512_));
 sg13g2_or2_1 _11505_ (.X(_06513_),
    .B(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .A(_00260_));
 sg13g2_o21ai_1 _11506_ (.B1(_06513_),
    .Y(_06514_),
    .A1(_00259_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][13] ));
 sg13g2_a22oi_1 _11507_ (.Y(_06515_),
    .B1(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .B2(_00260_),
    .A2(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .A1(_00261_));
 sg13g2_nor2b_1 _11508_ (.A(_06514_),
    .B_N(_06515_),
    .Y(_06516_));
 sg13g2_nand4_1 _11509_ (.B(_06511_),
    .C(_06512_),
    .A(_06509_),
    .Y(_06517_),
    .D(_06516_));
 sg13g2_o21ai_1 _11510_ (.B1(_06515_),
    .Y(_06518_),
    .A1(_06509_),
    .A2(_06514_));
 sg13g2_nand2b_1 _11511_ (.Y(_06519_),
    .B(_06518_),
    .A_N(_06510_));
 sg13g2_nand2_1 _11512_ (.Y(_06520_),
    .A(\soc_inst.pwm_ena[1] ),
    .B(_06519_));
 sg13g2_nor2_1 _11513_ (.A(net4795),
    .B(net4655),
    .Y(_06521_));
 sg13g2_nand2_1 _11514_ (.Y(_06522_),
    .A(net4797),
    .B(net4714));
 sg13g2_nand2_2 _11515_ (.Y(_06523_),
    .A(net4794),
    .B(_06287_));
 sg13g2_nor2_2 _11516_ (.A(net4643),
    .B(_06523_),
    .Y(_06524_));
 sg13g2_or2_1 _11517_ (.X(_06525_),
    .B(_06523_),
    .A(net4643));
 sg13g2_nand3_1 _11518_ (.B(net4787),
    .C(_05896_),
    .A(net4785),
    .Y(_06526_));
 sg13g2_nor2_1 _11519_ (.A(_06525_),
    .B(_06526_),
    .Y(_06527_));
 sg13g2_nor2_1 _11520_ (.A(_06520_),
    .B(net4002),
    .Y(_06528_));
 sg13g2_o21ai_1 _11521_ (.B1(_06528_),
    .Y(_06529_),
    .A1(_06508_),
    .A2(_06517_));
 sg13g2_nor2_1 _11522_ (.A(net148),
    .B(net3738),
    .Y(_00107_));
 sg13g2_xnor2_1 _11523_ (.Y(_06530_),
    .A(net2356),
    .B(net148));
 sg13g2_nor2_1 _11524_ (.A(net3738),
    .B(_06530_),
    .Y(_00114_));
 sg13g2_nor3_1 _11525_ (.A(_05573_),
    .B(_05574_),
    .C(_05575_),
    .Y(_06531_));
 sg13g2_a21oi_1 _11526_ (.A1(\soc_inst.pwm_inst.channel_counter[1][1] ),
    .A2(net148),
    .Y(_06532_),
    .B1(net910));
 sg13g2_nor3_1 _11527_ (.A(net3738),
    .B(_06531_),
    .C(net911),
    .Y(_00115_));
 sg13g2_nor2_1 _11528_ (.A(net2242),
    .B(_06531_),
    .Y(_06533_));
 sg13g2_and2_1 _11529_ (.A(net2242),
    .B(_06531_),
    .X(_06534_));
 sg13g2_nor3_1 _11530_ (.A(net3738),
    .B(net2243),
    .C(_06534_),
    .Y(_00116_));
 sg13g2_and2_1 _11531_ (.A(net2321),
    .B(_06534_),
    .X(_06535_));
 sg13g2_nor2_1 _11532_ (.A(net2321),
    .B(_06534_),
    .Y(_06536_));
 sg13g2_nor3_1 _11533_ (.A(net3737),
    .B(_06535_),
    .C(_06536_),
    .Y(_00117_));
 sg13g2_nor2_1 _11534_ (.A(net2481),
    .B(_06535_),
    .Y(_06537_));
 sg13g2_and2_1 _11535_ (.A(net2481),
    .B(_06535_),
    .X(_06538_));
 sg13g2_nor3_1 _11536_ (.A(net3737),
    .B(_06537_),
    .C(_06538_),
    .Y(_00118_));
 sg13g2_and2_1 _11537_ (.A(net2446),
    .B(_06538_),
    .X(_06539_));
 sg13g2_nor2_1 _11538_ (.A(net2446),
    .B(_06538_),
    .Y(_06540_));
 sg13g2_nor3_1 _11539_ (.A(net3737),
    .B(_06539_),
    .C(net2447),
    .Y(_00119_));
 sg13g2_nor2_1 _11540_ (.A(net2644),
    .B(_06539_),
    .Y(_06541_));
 sg13g2_and2_1 _11541_ (.A(net2644),
    .B(_06539_),
    .X(_06542_));
 sg13g2_nor3_1 _11542_ (.A(net3737),
    .B(_06541_),
    .C(_06542_),
    .Y(_00120_));
 sg13g2_nor2_1 _11543_ (.A(net2390),
    .B(_06542_),
    .Y(_06543_));
 sg13g2_and2_1 _11544_ (.A(net2390),
    .B(_06542_),
    .X(_06544_));
 sg13g2_nor3_1 _11545_ (.A(net3737),
    .B(net2391),
    .C(_06544_),
    .Y(_00121_));
 sg13g2_xnor2_1 _11546_ (.Y(_06545_),
    .A(net2614),
    .B(_06544_));
 sg13g2_nor2_1 _11547_ (.A(net3737),
    .B(_06545_),
    .Y(_00122_));
 sg13g2_a21oi_1 _11548_ (.A1(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .A2(_06544_),
    .Y(_06546_),
    .B1(net2271));
 sg13g2_and3_1 _11549_ (.X(_06547_),
    .A(net2271),
    .B(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .C(_06544_));
 sg13g2_nor3_1 _11550_ (.A(net3737),
    .B(net2272),
    .C(_06547_),
    .Y(_00108_));
 sg13g2_and2_1 _11551_ (.A(net2467),
    .B(_06547_),
    .X(_06548_));
 sg13g2_nor2_1 _11552_ (.A(net2467),
    .B(_06547_),
    .Y(_06549_));
 sg13g2_nor3_1 _11553_ (.A(net3737),
    .B(_06548_),
    .C(net2468),
    .Y(_00109_));
 sg13g2_nor2_1 _11554_ (.A(net2392),
    .B(_06548_),
    .Y(_06550_));
 sg13g2_and2_1 _11555_ (.A(net2392),
    .B(_06548_),
    .X(_06551_));
 sg13g2_nor3_1 _11556_ (.A(net3738),
    .B(net2393),
    .C(_06551_),
    .Y(_00110_));
 sg13g2_and2_1 _11557_ (.A(net2300),
    .B(_06551_),
    .X(_06552_));
 sg13g2_nor2_1 _11558_ (.A(net2300),
    .B(_06551_),
    .Y(_06553_));
 sg13g2_nor3_1 _11559_ (.A(net3738),
    .B(_06552_),
    .C(net2301),
    .Y(_00111_));
 sg13g2_xnor2_1 _11560_ (.Y(_06554_),
    .A(net2549),
    .B(_06552_));
 sg13g2_nor2_1 _11561_ (.A(net3738),
    .B(_06554_),
    .Y(_00112_));
 sg13g2_a21oi_1 _11562_ (.A1(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .A2(_06552_),
    .Y(_06555_),
    .B1(net1235));
 sg13g2_nor2_1 _11563_ (.A(net3738),
    .B(net1236),
    .Y(_00113_));
 sg13g2_or2_1 _11564_ (.X(_06556_),
    .B(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .A(_00236_));
 sg13g2_nor2_1 _11565_ (.A(_00231_),
    .B(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .Y(_06557_));
 sg13g2_nor2_1 _11566_ (.A(_00230_),
    .B(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .Y(_06558_));
 sg13g2_a22oi_1 _11567_ (.Y(_06559_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .B2(_00231_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .A1(_00232_));
 sg13g2_o21ai_1 _11568_ (.B1(_06559_),
    .Y(_06560_),
    .A1(_06557_),
    .A2(_06558_));
 sg13g2_nor2_1 _11569_ (.A(_00232_),
    .B(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .Y(_06561_));
 sg13g2_o21ai_1 _11570_ (.B1(_06560_),
    .Y(_06562_),
    .A1(_00233_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][3] ));
 sg13g2_a22oi_1 _11571_ (.Y(_06563_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .B2(_00233_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .A1(_00234_));
 sg13g2_o21ai_1 _11572_ (.B1(_06563_),
    .Y(_06564_),
    .A1(_06561_),
    .A2(_06562_));
 sg13g2_nor2_1 _11573_ (.A(_00234_),
    .B(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .Y(_06565_));
 sg13g2_o21ai_1 _11574_ (.B1(_06564_),
    .Y(_06566_),
    .A1(_00235_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][5] ));
 sg13g2_a22oi_1 _11575_ (.Y(_06567_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .B2(_00235_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .A1(_00236_));
 sg13g2_o21ai_1 _11576_ (.B1(_06567_),
    .Y(_06568_),
    .A1(_06565_),
    .A2(_06566_));
 sg13g2_a22oi_1 _11577_ (.Y(_06569_),
    .B1(_06556_),
    .B2(_06568_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .A1(_00237_));
 sg13g2_nor2_1 _11578_ (.A(_00237_),
    .B(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .Y(_06570_));
 sg13g2_nor2_1 _11579_ (.A(_00239_),
    .B(net5127),
    .Y(_06571_));
 sg13g2_nor2_1 _11580_ (.A(_00238_),
    .B(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .Y(_06572_));
 sg13g2_nor4_1 _11581_ (.A(_06569_),
    .B(_06570_),
    .C(_06571_),
    .D(_06572_),
    .Y(_06573_));
 sg13g2_a221oi_1 _11582_ (.B2(_00238_),
    .C1(_06573_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .A1(_00239_),
    .Y(_06574_),
    .A2(net5127));
 sg13g2_nand3_1 _11583_ (.B(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .C(_06571_),
    .A(_00238_),
    .Y(_06575_));
 sg13g2_o21ai_1 _11584_ (.B1(_06575_),
    .Y(_06576_),
    .A1(_00240_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][10] ));
 sg13g2_nor2_1 _11585_ (.A(_06574_),
    .B(_06576_),
    .Y(_06577_));
 sg13g2_a221oi_1 _11586_ (.B2(_00240_),
    .C1(_06577_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .A1(_00241_),
    .Y(_06578_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][11] ));
 sg13g2_a22oi_1 _11587_ (.Y(_06579_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .B2(_00244_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .A1(_00245_));
 sg13g2_nor2_1 _11588_ (.A(_00244_),
    .B(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .Y(_06580_));
 sg13g2_nor2_1 _11589_ (.A(_00245_),
    .B(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .Y(_06581_));
 sg13g2_nand2b_1 _11590_ (.Y(_06582_),
    .B(_06579_),
    .A_N(_06581_));
 sg13g2_a22oi_1 _11591_ (.Y(_06583_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .B2(_00242_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .A1(_00243_));
 sg13g2_nor2_1 _11592_ (.A(_00243_),
    .B(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .Y(_06584_));
 sg13g2_nor2_1 _11593_ (.A(_00241_),
    .B(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .Y(_06585_));
 sg13g2_o21ai_1 _11594_ (.B1(_06583_),
    .Y(_06586_),
    .A1(_00242_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][12] ));
 sg13g2_or3_1 _11595_ (.A(_06584_),
    .B(_06585_),
    .C(_06586_),
    .X(_06587_));
 sg13g2_nor4_1 _11596_ (.A(_06578_),
    .B(_06580_),
    .C(_06582_),
    .D(_06587_),
    .Y(_06588_));
 sg13g2_nor4_1 _11597_ (.A(_06580_),
    .B(_06582_),
    .C(_06583_),
    .D(_06584_),
    .Y(_06589_));
 sg13g2_o21ai_1 _11598_ (.B1(net2984),
    .Y(_06590_),
    .A1(_06579_),
    .A2(_06581_));
 sg13g2_nor2_2 _11599_ (.A(_06289_),
    .B(net4643),
    .Y(_06591_));
 sg13g2_nand2_2 _11600_ (.Y(_06592_),
    .A(_06288_),
    .B(net4264));
 sg13g2_nor2_2 _11601_ (.A(_06526_),
    .B(_06592_),
    .Y(_06593_));
 sg13g2_or4_1 _11602_ (.A(_06588_),
    .B(_06589_),
    .C(_06590_),
    .D(net3997),
    .X(_06594_));
 sg13g2_nor2_1 _11603_ (.A(net186),
    .B(net3717),
    .Y(_00091_));
 sg13g2_xnor2_1 _11604_ (.Y(_06595_),
    .A(net2524),
    .B(net186));
 sg13g2_nor2_1 _11605_ (.A(net3717),
    .B(_06595_),
    .Y(_00098_));
 sg13g2_a21oi_1 _11606_ (.A1(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .A2(net186),
    .Y(_06596_),
    .B1(net1588));
 sg13g2_and3_1 _11607_ (.X(_06597_),
    .A(net1588),
    .B(net2524),
    .C(net186));
 sg13g2_nor3_1 _11608_ (.A(net3717),
    .B(net1589),
    .C(_06597_),
    .Y(_00099_));
 sg13g2_nor2_1 _11609_ (.A(net2568),
    .B(_06597_),
    .Y(_06598_));
 sg13g2_and2_1 _11610_ (.A(net2568),
    .B(_06597_),
    .X(_06599_));
 sg13g2_nor3_1 _11611_ (.A(net3717),
    .B(_06598_),
    .C(_06599_),
    .Y(_00100_));
 sg13g2_and2_1 _11612_ (.A(net2471),
    .B(_06599_),
    .X(_06600_));
 sg13g2_nor2_1 _11613_ (.A(net2471),
    .B(_06599_),
    .Y(_06601_));
 sg13g2_nor3_1 _11614_ (.A(net3717),
    .B(_06600_),
    .C(net2472),
    .Y(_00101_));
 sg13g2_nor2_1 _11615_ (.A(net2295),
    .B(_06600_),
    .Y(_06602_));
 sg13g2_and2_1 _11616_ (.A(net2295),
    .B(_06600_),
    .X(_06603_));
 sg13g2_nor3_1 _11617_ (.A(net3717),
    .B(net2296),
    .C(_06603_),
    .Y(_00102_));
 sg13g2_and2_1 _11618_ (.A(net2317),
    .B(_06603_),
    .X(_06604_));
 sg13g2_nor2_1 _11619_ (.A(net2317),
    .B(_06603_),
    .Y(_06605_));
 sg13g2_nor3_1 _11620_ (.A(_06594_),
    .B(_06604_),
    .C(net2318),
    .Y(_00103_));
 sg13g2_nor2_1 _11621_ (.A(net2492),
    .B(_06604_),
    .Y(_06606_));
 sg13g2_and2_1 _11622_ (.A(net2492),
    .B(_06604_),
    .X(_06607_));
 sg13g2_nor3_1 _11623_ (.A(net3716),
    .B(_06606_),
    .C(_06607_),
    .Y(_00104_));
 sg13g2_nor2_1 _11624_ (.A(net2626),
    .B(_06607_),
    .Y(_06608_));
 sg13g2_and2_1 _11625_ (.A(net2626),
    .B(_06607_),
    .X(_06609_));
 sg13g2_nor3_1 _11626_ (.A(net3716),
    .B(_06608_),
    .C(_06609_),
    .Y(_00105_));
 sg13g2_xnor2_1 _11627_ (.Y(_06610_),
    .A(net5127),
    .B(_06609_));
 sg13g2_nor2_1 _11628_ (.A(net3716),
    .B(_06610_),
    .Y(_00106_));
 sg13g2_a21oi_1 _11629_ (.A1(net5127),
    .A2(_06609_),
    .Y(_06611_),
    .B1(net1379));
 sg13g2_and3_1 _11630_ (.X(_06612_),
    .A(net1379),
    .B(net5127),
    .C(_06609_));
 sg13g2_nor3_1 _11631_ (.A(net3716),
    .B(net1380),
    .C(_06612_),
    .Y(_00092_));
 sg13g2_and2_1 _11632_ (.A(net2431),
    .B(_06612_),
    .X(_06613_));
 sg13g2_nor2_1 _11633_ (.A(net2431),
    .B(_06612_),
    .Y(_06614_));
 sg13g2_nor3_1 _11634_ (.A(net3716),
    .B(_06613_),
    .C(net2432),
    .Y(_00093_));
 sg13g2_nor2_1 _11635_ (.A(net2569),
    .B(_06613_),
    .Y(_06615_));
 sg13g2_and2_1 _11636_ (.A(net2569),
    .B(_06613_),
    .X(_06616_));
 sg13g2_nor3_1 _11637_ (.A(net3716),
    .B(_06615_),
    .C(_06616_),
    .Y(_00094_));
 sg13g2_and2_1 _11638_ (.A(net2544),
    .B(_06616_),
    .X(_06617_));
 sg13g2_nor2_1 _11639_ (.A(net2544),
    .B(_06616_),
    .Y(_06618_));
 sg13g2_nor3_1 _11640_ (.A(net3716),
    .B(_06617_),
    .C(net2545),
    .Y(_00095_));
 sg13g2_xnor2_1 _11641_ (.Y(_06619_),
    .A(net2658),
    .B(_06617_));
 sg13g2_nor2_1 _11642_ (.A(net3716),
    .B(_06619_),
    .Y(_00096_));
 sg13g2_a21oi_1 _11643_ (.A1(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .A2(_06617_),
    .Y(_06620_),
    .B1(net690));
 sg13g2_nor2_1 _11644_ (.A(net3717),
    .B(net691),
    .Y(_00097_));
 sg13g2_nand3b_1 _11645_ (.B(net4278),
    .C(_00262_),
    .Y(\soc_inst.flash_cs_n ),
    .A_N(net5123));
 sg13g2_nor2b_1 _11646_ (.A(\soc_inst.core_mem_addr[25] ),
    .B_N(_00262_),
    .Y(_06621_));
 sg13g2_nor4_1 _11647_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.stop ),
    .B(\soc_inst.core_mem_addr[27] ),
    .C(\soc_inst.core_mem_addr[26] ),
    .D(net5074),
    .Y(_06622_));
 sg13g2_nand4_1 _11648_ (.B(_06045_),
    .C(_06621_),
    .A(\soc_inst.core_mem_addr[24] ),
    .Y(\soc_inst.mem_ctrl.ram_cs_n ),
    .D(_06622_));
 sg13g2_nor2_1 _11649_ (.A(_00274_),
    .B(_00273_),
    .Y(_06623_));
 sg13g2_nand2b_1 _11650_ (.Y(_06624_),
    .B(_06623_),
    .A_N(\soc_inst.cpu_core.ex_instr[3] ));
 sg13g2_nand3_1 _11651_ (.B(\soc_inst.cpu_core.ex_instr[2] ),
    .C(_06623_),
    .A(\soc_inst.cpu_core.ex_instr[3] ),
    .Y(_06625_));
 sg13g2_nand2_1 _11652_ (.Y(_06626_),
    .A(_06624_),
    .B(_06625_));
 sg13g2_and4_1 _11653_ (.A(_00275_),
    .B(\soc_inst.cpu_core.ex_instr[5] ),
    .C(\soc_inst.cpu_core.ex_instr[6] ),
    .D(_06626_),
    .X(_06627_));
 sg13g2_nand4_1 _11654_ (.B(\soc_inst.cpu_core.ex_instr[5] ),
    .C(\soc_inst.cpu_core.ex_instr[6] ),
    .A(_00275_),
    .Y(_06628_),
    .D(_06626_));
 sg13g2_nand2b_1 _11655_ (.Y(_06629_),
    .B(_00275_),
    .A_N(\soc_inst.cpu_core.ex_instr[6] ));
 sg13g2_nor2_1 _11656_ (.A(net2014),
    .B(_06624_),
    .Y(_06630_));
 sg13g2_nor2_1 _11657_ (.A(\soc_inst.cpu_core.ex_instr[5] ),
    .B(_06629_),
    .Y(_06631_));
 sg13g2_nor2_1 _11658_ (.A(\soc_inst.cpu_core.ex_instr[5] ),
    .B(_06625_),
    .Y(_06632_));
 sg13g2_nor2_1 _11659_ (.A(_06630_),
    .B(_06632_),
    .Y(_06633_));
 sg13g2_o21ai_1 _11660_ (.B1(_06628_),
    .Y(_06634_),
    .A1(_06629_),
    .A2(_06633_));
 sg13g2_inv_1 _11661_ (.Y(_06635_),
    .A(_06634_));
 sg13g2_nand2_1 _11662_ (.Y(_06636_),
    .A(\soc_inst.cpu_core.ex_instr[5] ),
    .B(_06630_));
 sg13g2_nand2_1 _11663_ (.Y(_06637_),
    .A(\soc_inst.cpu_core.ex_instr[6] ),
    .B(_06636_));
 sg13g2_nor2_1 _11664_ (.A(_00275_),
    .B(_06624_),
    .Y(_06638_));
 sg13g2_a21oi_1 _11665_ (.A1(_06637_),
    .A2(_06638_),
    .Y(_06639_),
    .B1(_06634_));
 sg13g2_a21o_2 _11666_ (.A2(_06638_),
    .A1(_06637_),
    .B1(_06634_),
    .X(_06640_));
 sg13g2_and2_1 _11667_ (.A(\soc_inst.cpu_core.ex_branch_target[0] ),
    .B(net4196),
    .X(_06641_));
 sg13g2_nand2_1 _11668_ (.Y(_06642_),
    .A(\soc_inst.cpu_core.ex_branch_target[0] ),
    .B(net4196));
 sg13g2_nand2_1 _11669_ (.Y(_06643_),
    .A(net4055),
    .B(net4101));
 sg13g2_nand3b_1 _11670_ (.B(\soc_inst.cpu_core.ex_alu_result[0] ),
    .C(\soc_inst.cpu_core.ex_funct3[0] ),
    .Y(_06644_),
    .A_N(\soc_inst.cpu_core.ex_funct3[1] ));
 sg13g2_nor2b_1 _11671_ (.A(\soc_inst.cpu_core.ex_funct3[0] ),
    .B_N(\soc_inst.cpu_core.ex_funct3[1] ),
    .Y(_06645_));
 sg13g2_o21ai_1 _11672_ (.B1(_06645_),
    .Y(_06646_),
    .A1(\soc_inst.cpu_core.ex_alu_result[1] ),
    .A2(\soc_inst.cpu_core.ex_alu_result[0] ));
 sg13g2_a21o_1 _11673_ (.A2(_06646_),
    .A1(_06644_),
    .B1(\soc_inst.cpu_core.ex_funct3[2] ),
    .X(_06647_));
 sg13g2_nand2_1 _11674_ (.Y(_06648_),
    .A(_06644_),
    .B(_06647_));
 sg13g2_nand3_1 _11675_ (.B(_06631_),
    .C(_06648_),
    .A(_06630_),
    .Y(_06649_));
 sg13g2_or2_1 _11676_ (.X(_06650_),
    .B(_06647_),
    .A(_06629_));
 sg13g2_o21ai_1 _11677_ (.B1(_06649_),
    .Y(_06651_),
    .A1(_06636_),
    .A2(_06650_));
 sg13g2_nor2_1 _11678_ (.A(net3993),
    .B(net4052),
    .Y(_06652_));
 sg13g2_or2_1 _11679_ (.X(_06653_),
    .B(net4050),
    .A(net3995));
 sg13g2_nor3_1 _11680_ (.A(\soc_inst.cpu_core.ex_is_ecall ),
    .B(\soc_inst.cpu_core.ex_is_ebreak ),
    .C(_06653_),
    .Y(_06654_));
 sg13g2_or3_1 _11681_ (.A(\soc_inst.cpu_core.ex_is_ecall ),
    .B(\soc_inst.cpu_core.ex_is_ebreak ),
    .C(_06653_),
    .X(_06655_));
 sg13g2_nor3_1 _11682_ (.A(net4974),
    .B(_05720_),
    .C(net3859),
    .Y(_00024_));
 sg13g2_and3_1 _11683_ (.X(_00025_),
    .A(net4752),
    .B(net350),
    .C(net3862));
 sg13g2_nor2_1 _11684_ (.A(net4752),
    .B(net675),
    .Y(_06656_));
 sg13g2_or3_1 _11685_ (.A(_00024_),
    .B(_00025_),
    .C(_06656_),
    .X(_00026_));
 sg13g2_nor2_2 _11686_ (.A(\soc_inst.cpu_core.id_int_is_interrupt ),
    .B(net3858),
    .Y(_06657_));
 sg13g2_nand2_1 _11687_ (.Y(_06658_),
    .A(_05479_),
    .B(net3860));
 sg13g2_nor2_1 _11688_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .Y(_06659_));
 sg13g2_nor2_1 _11689_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .Y(_06660_));
 sg13g2_and2_1 _11690_ (.A(net4712),
    .B(_06660_),
    .X(_06661_));
 sg13g2_nand2_2 _11691_ (.Y(_06662_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[9] ));
 sg13g2_nor2_2 _11692_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .Y(_06663_));
 sg13g2_nor2b_2 _11693_ (.A(_06662_),
    .B_N(_06663_),
    .Y(_06664_));
 sg13g2_nand2b_1 _11694_ (.Y(_06665_),
    .B(_06663_),
    .A_N(_06662_));
 sg13g2_nor2_1 _11695_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .Y(_06666_));
 sg13g2_nor3_1 _11696_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .C(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .Y(_06667_));
 sg13g2_nor2_1 _11697_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .Y(_06668_));
 sg13g2_and2_1 _11698_ (.A(_06666_),
    .B(_06668_),
    .X(_06669_));
 sg13g2_nand2_2 _11699_ (.Y(_06670_),
    .A(_06664_),
    .B(_06669_));
 sg13g2_and3_1 _11700_ (.X(_06671_),
    .A(_06661_),
    .B(_06664_),
    .C(_06669_));
 sg13g2_nand3_1 _11701_ (.B(_06664_),
    .C(_06669_),
    .A(_06661_),
    .Y(_06672_));
 sg13g2_nor2_2 _11702_ (.A(net4871),
    .B(net4876),
    .Y(_06673_));
 sg13g2_or2_1 _11703_ (.X(_06674_),
    .B(net4876),
    .A(net4871));
 sg13g2_nor2_2 _11704_ (.A(net4872),
    .B(net4870),
    .Y(_06675_));
 sg13g2_nor2_2 _11705_ (.A(net4869),
    .B(net4711),
    .Y(_06676_));
 sg13g2_nand3_1 _11706_ (.B(\soc_inst.cpu_core.mem_instr[5] ),
    .C(\soc_inst.cpu_core.mem_instr[6] ),
    .A(_05403_),
    .Y(_06677_));
 sg13g2_or4_1 _11707_ (.A(_00271_),
    .B(_00270_),
    .C(\soc_inst.cpu_core.mem_instr[3] ),
    .D(\soc_inst.cpu_core.mem_instr[2] ),
    .X(_06678_));
 sg13g2_nor3_2 _11708_ (.A(_06676_),
    .B(_06677_),
    .C(_06678_),
    .Y(_06679_));
 sg13g2_or3_1 _11709_ (.A(_06676_),
    .B(_06677_),
    .C(_06678_),
    .X(_06680_));
 sg13g2_nand3_1 _11710_ (.B(net4712),
    .C(_06669_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .Y(_06681_));
 sg13g2_nor2b_1 _11711_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .B_N(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .Y(_06682_));
 sg13g2_nand3_1 _11712_ (.B(_06661_),
    .C(_06682_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .Y(_06683_));
 sg13g2_a21oi_1 _11713_ (.A1(_06681_),
    .A2(_06683_),
    .Y(_06684_),
    .B1(_06662_));
 sg13g2_nand4_1 _11714_ (.B(_06661_),
    .C(_06666_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .Y(_06685_),
    .D(_06682_));
 sg13g2_nor2_1 _11715_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .B(_06685_),
    .Y(_06686_));
 sg13g2_o21ai_1 _11716_ (.B1(_06663_),
    .Y(_06687_),
    .A1(_06684_),
    .A2(_06686_));
 sg13g2_nor2_1 _11717_ (.A(_05414_),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .Y(_06688_));
 sg13g2_nand2_1 _11718_ (.Y(_06689_),
    .A(net4712),
    .B(_06688_));
 sg13g2_and3_2 _11719_ (.X(_06690_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .B(_06664_),
    .C(_06667_));
 sg13g2_nor2b_1 _11720_ (.A(_06689_),
    .B_N(_06690_),
    .Y(_06691_));
 sg13g2_nand2b_2 _11721_ (.Y(_06692_),
    .B(_06690_),
    .A_N(_06689_));
 sg13g2_nor2b_1 _11722_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .B_N(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .Y(_06693_));
 sg13g2_nand2_1 _11723_ (.Y(_06694_),
    .A(_06660_),
    .B(_06693_));
 sg13g2_nor2_2 _11724_ (.A(_06670_),
    .B(_06694_),
    .Y(_06695_));
 sg13g2_nand2_1 _11725_ (.Y(_06696_),
    .A(_06688_),
    .B(_06693_));
 sg13g2_nor2_1 _11726_ (.A(_06670_),
    .B(_06696_),
    .Y(_06697_));
 sg13g2_nand3_1 _11727_ (.B(_06659_),
    .C(_06690_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .Y(_06698_));
 sg13g2_nand2b_1 _11728_ (.Y(_06699_),
    .B(_06698_),
    .A_N(net4185));
 sg13g2_nand2b_1 _11729_ (.Y(_06700_),
    .B(net4712),
    .A_N(_06660_));
 sg13g2_nand2_1 _11730_ (.Y(_06701_),
    .A(_06694_),
    .B(_06700_));
 sg13g2_nand2_2 _11731_ (.Y(_06702_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[11] ));
 sg13g2_nor2_1 _11732_ (.A(_06662_),
    .B(_06702_),
    .Y(_06703_));
 sg13g2_nor2b_1 _11733_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .B_N(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .Y(_06704_));
 sg13g2_nand4_1 _11734_ (.B(_06701_),
    .C(_06703_),
    .A(_06668_),
    .Y(_06705_),
    .D(_06704_));
 sg13g2_and2_1 _11735_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .X(_06706_));
 sg13g2_nor4_1 _11736_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .C(_06702_),
    .D(_06706_),
    .Y(_06707_));
 sg13g2_and4_1 _11737_ (.A(net4712),
    .B(_06666_),
    .C(_06682_),
    .D(_06707_),
    .X(_06708_));
 sg13g2_and3_1 _11738_ (.X(_06709_),
    .A(net4712),
    .B(_06669_),
    .C(_06707_));
 sg13g2_nor2_1 _11739_ (.A(net4239),
    .B(net4236),
    .Y(_06710_));
 sg13g2_and2_1 _11740_ (.A(_06661_),
    .B(_06690_),
    .X(_06711_));
 sg13g2_nor2_1 _11741_ (.A(_06670_),
    .B(_06689_),
    .Y(_06712_));
 sg13g2_and3_2 _11742_ (.X(_06713_),
    .A(_06660_),
    .B(_06690_),
    .C(_06693_));
 sg13g2_nor4_1 _11743_ (.A(net4251),
    .B(net4181),
    .C(_06712_),
    .D(_06713_),
    .Y(_06714_));
 sg13g2_nand3_1 _11744_ (.B(_06710_),
    .C(_06714_),
    .A(_06705_),
    .Y(_06715_));
 sg13g2_and3_2 _11745_ (.X(_06716_),
    .A(net4712),
    .B(_06669_),
    .C(_06707_));
 sg13g2_nor4_1 _11746_ (.A(net4189),
    .B(_06695_),
    .C(_06699_),
    .D(_06715_),
    .Y(_06717_));
 sg13g2_a21oi_2 _11747_ (.B1(net4240),
    .Y(_06718_),
    .A2(_06717_),
    .A1(_06687_));
 sg13g2_nand2_2 _11748_ (.Y(_06719_),
    .A(net4710),
    .B(net3946));
 sg13g2_nand3_1 _11749_ (.B(net4710),
    .C(net3946),
    .A(net4256),
    .Y(_06720_));
 sg13g2_or3_1 _11750_ (.A(_06676_),
    .B(_06677_),
    .C(_06678_),
    .X(_06721_));
 sg13g2_nand3_1 _11751_ (.B(_06661_),
    .C(_06667_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .Y(_06722_));
 sg13g2_nor2_2 _11752_ (.A(_06665_),
    .B(_06722_),
    .Y(_06723_));
 sg13g2_nand3_1 _11753_ (.B(net4712),
    .C(_06690_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .Y(_06724_));
 sg13g2_nand2b_1 _11754_ (.Y(_06725_),
    .B(_06724_),
    .A_N(net4185));
 sg13g2_nand4_1 _11755_ (.B(_06701_),
    .C(_06703_),
    .A(_06668_),
    .Y(_06726_),
    .D(_06704_));
 sg13g2_nor2_1 _11756_ (.A(net4254),
    .B(net4239),
    .Y(_06727_));
 sg13g2_nor4_1 _11757_ (.A(net4189),
    .B(_06695_),
    .C(net4236),
    .D(_06713_),
    .Y(_06728_));
 sg13g2_nand3_1 _11758_ (.B(_06727_),
    .C(_06728_),
    .A(_06726_),
    .Y(_06729_));
 sg13g2_nor4_1 _11759_ (.A(_06712_),
    .B(_06723_),
    .C(_06725_),
    .D(_06729_),
    .Y(_06730_));
 sg13g2_a21oi_1 _11760_ (.A1(_06687_),
    .A2(_06730_),
    .Y(_06731_),
    .B1(_06721_));
 sg13g2_nand2_1 _11761_ (.Y(_06732_),
    .A(net4710),
    .B(_06731_));
 sg13g2_nor2_2 _11762_ (.A(_06672_),
    .B(_06732_),
    .Y(_06733_));
 sg13g2_nor2_2 _11763_ (.A(net3796),
    .B(_06733_),
    .Y(_06734_));
 sg13g2_nand2_1 _11764_ (.Y(_06735_),
    .A(net5054),
    .B(net2084));
 sg13g2_o21ai_1 _11765_ (.B1(_06735_),
    .Y(_06736_),
    .A1(net5054),
    .A2(_05518_));
 sg13g2_nand2_1 _11766_ (.Y(_06737_),
    .A(_06734_),
    .B(_06736_));
 sg13g2_and2_1 _11767_ (.A(net4874),
    .B(net4877),
    .X(_06738_));
 sg13g2_or2_1 _11768_ (.X(_06739_),
    .B(\soc_inst.cpu_core.mem_rs1_data[3] ),
    .A(net4868));
 sg13g2_o21ai_1 _11769_ (.B1(_06739_),
    .Y(_06740_),
    .A1(net4753),
    .A2(\soc_inst.cpu_core.mem_instr[18] ));
 sg13g2_inv_1 _11770_ (.Y(_06741_),
    .A(_06740_));
 sg13g2_nor2_1 _11771_ (.A(net4707),
    .B(_06740_),
    .Y(_06742_));
 sg13g2_a21oi_1 _11772_ (.A1(net4871),
    .A2(_06740_),
    .Y(_06743_),
    .B1(_06742_));
 sg13g2_o21ai_1 _11773_ (.B1(_06733_),
    .Y(_06744_),
    .A1(net2864),
    .A2(_06742_));
 sg13g2_o21ai_1 _11774_ (.B1(_06737_),
    .Y(_00063_),
    .A1(_06743_),
    .A2(_06744_));
 sg13g2_nor2_1 _11775_ (.A(_06692_),
    .B(_06719_),
    .Y(_06745_));
 sg13g2_nand3_1 _11776_ (.B(net4192),
    .C(net3946),
    .A(net4710),
    .Y(_06746_));
 sg13g2_nand2_2 _11777_ (.Y(_06747_),
    .A(net3799),
    .B(net3851));
 sg13g2_nand2b_1 _11778_ (.Y(_06748_),
    .B(net4871),
    .A_N(net4877));
 sg13g2_nor2b_1 _11779_ (.A(net4871),
    .B_N(net4876),
    .Y(_06749_));
 sg13g2_nand2_2 _11780_ (.Y(_06750_),
    .A(net4755),
    .B(net4877));
 sg13g2_and2_1 _11781_ (.A(_06748_),
    .B(_06750_),
    .X(_06751_));
 sg13g2_o21ai_1 _11782_ (.B1(net3851),
    .Y(_06752_),
    .A1(_06719_),
    .A2(net4707));
 sg13g2_or2_1 _11783_ (.X(_06753_),
    .B(\soc_inst.cpu_core.mem_rs1_data[0] ),
    .A(net4868));
 sg13g2_o21ai_1 _11784_ (.B1(_06753_),
    .Y(_06754_),
    .A1(net4753),
    .A2(\soc_inst.cpu_core.mem_instr[15] ));
 sg13g2_inv_1 _11785_ (.Y(_06755_),
    .A(_06754_));
 sg13g2_a21oi_1 _11786_ (.A1(net4191),
    .A2(_06754_),
    .Y(_06756_),
    .B1(net4229));
 sg13g2_a21oi_2 _11787_ (.B1(net4756),
    .Y(_06757_),
    .A2(_06755_),
    .A1(net4876));
 sg13g2_a21oi_1 _11788_ (.A1(net2664),
    .A2(_06757_),
    .Y(_06758_),
    .B1(_06756_));
 sg13g2_nand2_2 _11789_ (.Y(_06759_),
    .A(net2786),
    .B(net3862));
 sg13g2_inv_1 _11790_ (.Y(_06760_),
    .A(_06759_));
 sg13g2_nor2_1 _11791_ (.A(\soc_inst.cpu_core.id_pc[0] ),
    .B(_06759_),
    .Y(_06761_));
 sg13g2_nor2_1 _11792_ (.A(net1296),
    .B(net3861),
    .Y(_06762_));
 sg13g2_o21ai_1 _11793_ (.B1(net3851),
    .Y(_06763_),
    .A1(_06761_),
    .A2(_06762_));
 sg13g2_o21ai_1 _11794_ (.B1(_06763_),
    .Y(_06764_),
    .A1(net2664),
    .A2(_06747_));
 sg13g2_a21oi_1 _11795_ (.A1(_06752_),
    .A2(_06758_),
    .Y(_00058_),
    .B1(_06764_));
 sg13g2_or2_1 _11796_ (.X(_06765_),
    .B(\soc_inst.cpu_core.mem_rs1_data[1] ),
    .A(net4868));
 sg13g2_o21ai_1 _11797_ (.B1(_06765_),
    .Y(_06766_),
    .A1(net4753),
    .A2(\soc_inst.cpu_core.mem_instr[16] ));
 sg13g2_inv_1 _11798_ (.Y(_06767_),
    .A(_06766_));
 sg13g2_a21oi_1 _11799_ (.A1(net4191),
    .A2(_06766_),
    .Y(_06768_),
    .B1(net4229));
 sg13g2_a21oi_2 _11800_ (.B1(net4757),
    .Y(_06769_),
    .A2(_06767_),
    .A1(net4876));
 sg13g2_a21oi_1 _11801_ (.A1(net2843),
    .A2(_06769_),
    .Y(_06770_),
    .B1(_06768_));
 sg13g2_a22oi_1 _11802_ (.Y(_06771_),
    .B1(net3798),
    .B2(_05612_),
    .A2(net3859),
    .A1(_05735_));
 sg13g2_o21ai_1 _11803_ (.B1(_06771_),
    .Y(_06772_),
    .A1(net2838),
    .A2(_06759_));
 sg13g2_a22oi_1 _11804_ (.Y(_00059_),
    .B1(_06772_),
    .B2(net3851),
    .A2(_06770_),
    .A1(_06752_));
 sg13g2_or2_1 _11805_ (.X(_06773_),
    .B(\soc_inst.cpu_core.mem_rs1_data[2] ),
    .A(net4868));
 sg13g2_o21ai_1 _11806_ (.B1(_06773_),
    .Y(_06774_),
    .A1(net4753),
    .A2(\soc_inst.cpu_core.mem_instr[17] ));
 sg13g2_inv_1 _11807_ (.Y(_06775_),
    .A(_06774_));
 sg13g2_a21oi_1 _11808_ (.A1(net4191),
    .A2(_06774_),
    .Y(_06776_),
    .B1(net4230));
 sg13g2_a21oi_2 _11809_ (.B1(net4756),
    .Y(_06777_),
    .A2(_06775_),
    .A1(net4876));
 sg13g2_a21oi_1 _11810_ (.A1(net2721),
    .A2(_06777_),
    .Y(_06778_),
    .B1(_06776_));
 sg13g2_a22oi_1 _11811_ (.Y(_06779_),
    .B1(net3752),
    .B2(_05679_),
    .A2(net3859),
    .A1(_05736_));
 sg13g2_o21ai_1 _11812_ (.B1(_06779_),
    .Y(_06780_),
    .A1(net2721),
    .A2(net3793));
 sg13g2_a22oi_1 _11813_ (.Y(_00060_),
    .B1(_06780_),
    .B2(net3851),
    .A2(_06778_),
    .A1(_06752_));
 sg13g2_a21oi_1 _11814_ (.A1(net4191),
    .A2(_06740_),
    .Y(_06781_),
    .B1(net4230));
 sg13g2_a21oi_1 _11815_ (.A1(net4876),
    .A2(_06741_),
    .Y(_06782_),
    .B1(net4756));
 sg13g2_a21oi_1 _11816_ (.A1(net2902),
    .A2(_06782_),
    .Y(_06783_),
    .B1(_06781_));
 sg13g2_a22oi_1 _11817_ (.Y(_06784_),
    .B1(net3798),
    .B2(_05615_),
    .A2(net3859),
    .A1(_05737_));
 sg13g2_o21ai_1 _11818_ (.B1(_06784_),
    .Y(_06785_),
    .A1(net2878),
    .A2(_06759_));
 sg13g2_a22oi_1 _11819_ (.Y(_00061_),
    .B1(_06785_),
    .B2(net3851),
    .A2(_06783_),
    .A1(_06752_));
 sg13g2_or2_1 _11820_ (.X(_06786_),
    .B(\soc_inst.cpu_core.mem_rs1_data[4] ),
    .A(net4868));
 sg13g2_o21ai_1 _11821_ (.B1(_06786_),
    .Y(_06787_),
    .A1(net4753),
    .A2(\soc_inst.cpu_core.mem_instr[19] ));
 sg13g2_inv_1 _11822_ (.Y(_06788_),
    .A(_06787_));
 sg13g2_a21oi_1 _11823_ (.A1(net4191),
    .A2(_06787_),
    .Y(_06789_),
    .B1(net4229));
 sg13g2_a21oi_2 _11824_ (.B1(net4757),
    .Y(_06790_),
    .A2(_06788_),
    .A1(net4877));
 sg13g2_a21oi_1 _11825_ (.A1(net2775),
    .A2(_06790_),
    .Y(_06791_),
    .B1(_06789_));
 sg13g2_a22oi_1 _11826_ (.Y(_06792_),
    .B1(net3752),
    .B2(_05681_),
    .A2(net3859),
    .A1(_05738_));
 sg13g2_o21ai_1 _11827_ (.B1(_06792_),
    .Y(_06793_),
    .A1(net2775),
    .A2(net3793));
 sg13g2_a22oi_1 _11828_ (.Y(_00062_),
    .B1(_06793_),
    .B2(net3851),
    .A2(_06791_),
    .A1(_06752_));
 sg13g2_o21ai_1 _11829_ (.B1(_06652_),
    .Y(_06794_),
    .A1(net2306),
    .A2(net3793));
 sg13g2_nor2_1 _11830_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(_06698_),
    .Y(_06795_));
 sg13g2_nand3_1 _11831_ (.B(net3946),
    .C(net4095),
    .A(net4710),
    .Y(_06796_));
 sg13g2_nor2_2 _11832_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(_06724_),
    .Y(_06797_));
 sg13g2_o21ai_1 _11833_ (.B1(net3849),
    .Y(_06798_),
    .A1(_06719_),
    .A2(net4707));
 sg13g2_a21oi_1 _11834_ (.A1(_06754_),
    .A2(net4095),
    .Y(_06799_),
    .B1(net4229));
 sg13g2_a21oi_1 _11835_ (.A1(net2306),
    .A2(_06757_),
    .Y(_06800_),
    .B1(_06799_));
 sg13g2_a22oi_1 _11836_ (.Y(_00027_),
    .B1(_06798_),
    .B2(_06800_),
    .A2(net3849),
    .A1(_06794_));
 sg13g2_nor2_1 _11837_ (.A(net4106),
    .B(net3798),
    .Y(_06801_));
 sg13g2_a22oi_1 _11838_ (.Y(_06802_),
    .B1(_06801_),
    .B2(_06649_),
    .A2(net3798),
    .A1(net2450));
 sg13g2_a21oi_1 _11839_ (.A1(_06766_),
    .A2(net4095),
    .Y(_06803_),
    .B1(net4229));
 sg13g2_a21oi_1 _11840_ (.A1(net2450),
    .A2(_06769_),
    .Y(_06804_),
    .B1(_06803_));
 sg13g2_a22oi_1 _11841_ (.Y(_00038_),
    .B1(_06804_),
    .B2(_06798_),
    .A2(_06802_),
    .A1(net3849));
 sg13g2_nand2_2 _11842_ (.Y(_06805_),
    .A(\soc_inst.cpu_core.csr_file.mie[7] ),
    .B(\soc_inst.cpu_core.csr_file.mip_tip ));
 sg13g2_a21oi_1 _11843_ (.A1(\soc_inst.cpu_core.id_int_is_interrupt ),
    .A2(_06805_),
    .Y(_06806_),
    .B1(_06655_));
 sg13g2_or2_1 _11844_ (.X(_06807_),
    .B(_06806_),
    .A(net4053));
 sg13g2_o21ai_1 _11845_ (.B1(_06807_),
    .Y(_06808_),
    .A1(net2452),
    .A2(net3795));
 sg13g2_a21oi_1 _11846_ (.A1(_06774_),
    .A2(net4095),
    .Y(_06809_),
    .B1(net4230));
 sg13g2_a21oi_1 _11847_ (.A1(net2452),
    .A2(_06777_),
    .Y(_06810_),
    .B1(_06809_));
 sg13g2_a22oi_1 _11848_ (.Y(_00049_),
    .B1(_06810_),
    .B2(_06798_),
    .A2(_06808_),
    .A1(net3849));
 sg13g2_nor2b_1 _11849_ (.A(net574),
    .B_N(net1911),
    .Y(_06811_));
 sg13g2_nor3_1 _11850_ (.A(_06653_),
    .B(_06806_),
    .C(_06811_),
    .Y(_06812_));
 sg13g2_a21oi_1 _11851_ (.A1(net2531),
    .A2(net3799),
    .Y(_06813_),
    .B1(_06812_));
 sg13g2_a21oi_1 _11852_ (.A1(_06740_),
    .A2(net4095),
    .Y(_06814_),
    .B1(net4230));
 sg13g2_a21oi_1 _11853_ (.A1(net2531),
    .A2(_06782_),
    .Y(_06815_),
    .B1(_06814_));
 sg13g2_a22oi_1 _11854_ (.Y(_00051_),
    .B1(_06815_),
    .B2(_06798_),
    .A2(_06813_),
    .A1(net3849));
 sg13g2_and3_1 _11855_ (.X(_00052_),
    .A(net441),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11856_ (.X(_00053_),
    .A(net117),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11857_ (.X(_00054_),
    .A(net169),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11858_ (.X(_00055_),
    .A(net105),
    .B(net3804),
    .C(net3848));
 sg13g2_and3_1 _11859_ (.X(_00056_),
    .A(net94),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11860_ (.X(_00057_),
    .A(net99),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11861_ (.X(_00028_),
    .A(net101),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11862_ (.X(_00029_),
    .A(net95),
    .B(net3804),
    .C(net3847));
 sg13g2_and3_1 _11863_ (.X(_00030_),
    .A(net268),
    .B(net3803),
    .C(net3848));
 sg13g2_and3_1 _11864_ (.X(_00031_),
    .A(net511),
    .B(net3805),
    .C(net3848));
 sg13g2_and3_1 _11865_ (.X(_00032_),
    .A(net178),
    .B(net3803),
    .C(net3848));
 sg13g2_and3_1 _11866_ (.X(_00033_),
    .A(net93),
    .B(net3803),
    .C(net3846));
 sg13g2_and3_1 _11867_ (.X(_00034_),
    .A(net421),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11868_ (.X(_00035_),
    .A(net440),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11869_ (.X(_00036_),
    .A(net102),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11870_ (.X(_00037_),
    .A(net426),
    .B(net3803),
    .C(net3846));
 sg13g2_and3_1 _11871_ (.X(_00039_),
    .A(net318),
    .B(net3803),
    .C(net3846));
 sg13g2_and3_1 _11872_ (.X(_00040_),
    .A(net103),
    .B(net3801),
    .C(net3849));
 sg13g2_and3_1 _11873_ (.X(_00041_),
    .A(net96),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11874_ (.X(_00042_),
    .A(net120),
    .B(net3801),
    .C(net3849));
 sg13g2_and3_1 _11875_ (.X(_00043_),
    .A(net128),
    .B(net3803),
    .C(net3846));
 sg13g2_and3_1 _11876_ (.X(_00044_),
    .A(net181),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11877_ (.X(_00045_),
    .A(net100),
    .B(net3805),
    .C(net3847));
 sg13g2_and3_1 _11878_ (.X(_00046_),
    .A(net110),
    .B(net3803),
    .C(net3846));
 sg13g2_and3_1 _11879_ (.X(_00047_),
    .A(net240),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11880_ (.X(_00048_),
    .A(net157),
    .B(net3802),
    .C(net3845));
 sg13g2_and3_1 _11881_ (.X(_00050_),
    .A(net338),
    .B(net3802),
    .C(net3845));
 sg13g2_nor2_2 _11882_ (.A(_05414_),
    .B(_06698_),
    .Y(_06816_));
 sg13g2_nor2b_1 _11883_ (.A(_06719_),
    .B_N(net4089),
    .Y(_06817_));
 sg13g2_nand3_1 _11884_ (.B(net3946),
    .C(net4089),
    .A(net4710),
    .Y(_06818_));
 sg13g2_o21ai_1 _11885_ (.B1(net3839),
    .Y(_06819_),
    .A1(_06719_),
    .A2(net4707));
 sg13g2_nor2_2 _11886_ (.A(_05414_),
    .B(_06724_),
    .Y(_06820_));
 sg13g2_a21oi_1 _11887_ (.A1(_06754_),
    .A2(net4088),
    .Y(_06821_),
    .B1(net4229));
 sg13g2_a21oi_1 _11888_ (.A1(net2674),
    .A2(_06757_),
    .Y(_06822_),
    .B1(_06821_));
 sg13g2_nor2b_1 _11889_ (.A(net4053),
    .B_N(_06811_),
    .Y(_06823_));
 sg13g2_a221oi_1 _11890_ (.B2(net1296),
    .C1(net4059),
    .B1(net3989),
    .A1(\soc_inst.cpu_core.ex_alu_result[0] ),
    .Y(_06824_),
    .A2(net4052));
 sg13g2_o21ai_1 _11891_ (.B1(_06801_),
    .Y(_06825_),
    .A1(_00273_),
    .A2(_06824_));
 sg13g2_o21ai_1 _11892_ (.B1(_06825_),
    .Y(_06826_),
    .A1(net2674),
    .A2(net3793));
 sg13g2_a22oi_1 _11893_ (.Y(_00064_),
    .B1(_06826_),
    .B2(net3839),
    .A2(_06822_),
    .A1(_06819_));
 sg13g2_a221oi_1 _11894_ (.B2(net2185),
    .C1(net3993),
    .B1(net3989),
    .A1(\soc_inst.cpu_core.ex_alu_result[1] ),
    .Y(_06827_),
    .A2(net4052));
 sg13g2_nor2_1 _11895_ (.A(net2441),
    .B(net4102),
    .Y(_06828_));
 sg13g2_nor3_1 _11896_ (.A(_00274_),
    .B(_06827_),
    .C(_06828_),
    .Y(_06829_));
 sg13g2_a21oi_1 _11897_ (.A1(net2478),
    .A2(net3798),
    .Y(_06830_),
    .B1(_06829_));
 sg13g2_a21oi_1 _11898_ (.A1(_06766_),
    .A2(net4088),
    .Y(_06831_),
    .B1(net4229));
 sg13g2_a21oi_1 _11899_ (.A1(net2478),
    .A2(_06769_),
    .Y(_06832_),
    .B1(_06831_));
 sg13g2_a22oi_1 _11900_ (.Y(_00065_),
    .B1(_06832_),
    .B2(_06819_),
    .A2(_06830_),
    .A1(net3839));
 sg13g2_a221oi_1 _11901_ (.B2(net1070),
    .C1(net3994),
    .B1(net3989),
    .A1(net2978),
    .Y(_06833_),
    .A2(net4053));
 sg13g2_a221oi_1 _11902_ (.B2(_05707_),
    .C1(_06833_),
    .B1(net4106),
    .A1(_05475_),
    .Y(_06834_),
    .A2(net4059));
 sg13g2_a21oi_1 _11903_ (.A1(net2556),
    .A2(net3798),
    .Y(_06835_),
    .B1(_06834_));
 sg13g2_a21oi_1 _11904_ (.A1(_06774_),
    .A2(net4088),
    .Y(_06836_),
    .B1(net4230));
 sg13g2_a21oi_1 _11905_ (.A1(net2556),
    .A2(_06777_),
    .Y(_06837_),
    .B1(_06836_));
 sg13g2_a22oi_1 _11906_ (.Y(_00066_),
    .B1(_06837_),
    .B2(_06819_),
    .A2(_06835_),
    .A1(net3839));
 sg13g2_a221oi_1 _11907_ (.B2(net2245),
    .C1(net3993),
    .B1(net3989),
    .A1(\soc_inst.cpu_core.ex_alu_result[3] ),
    .Y(_06838_),
    .A2(net4052));
 sg13g2_nor2_1 _11908_ (.A(net2442),
    .B(net4057),
    .Y(_06839_));
 sg13g2_nor2_1 _11909_ (.A(net2384),
    .B(net4103),
    .Y(_06840_));
 sg13g2_nor4_1 _11910_ (.A(net3861),
    .B(_06838_),
    .C(_06839_),
    .D(_06840_),
    .Y(_06841_));
 sg13g2_a21oi_1 _11911_ (.A1(net2475),
    .A2(net3798),
    .Y(_06842_),
    .B1(_06841_));
 sg13g2_a21oi_1 _11912_ (.A1(_06740_),
    .A2(net4088),
    .Y(_06843_),
    .B1(net4230));
 sg13g2_a21oi_1 _11913_ (.A1(net2475),
    .A2(_06782_),
    .Y(_06844_),
    .B1(_06843_));
 sg13g2_a22oi_1 _11914_ (.Y(_00067_),
    .B1(_06844_),
    .B2(_06819_),
    .A2(_06842_),
    .A1(net3839));
 sg13g2_nand2_1 _11915_ (.Y(_06845_),
    .A(\soc_inst.cpu_core.ex_alu_result[4] ),
    .B(net4053));
 sg13g2_a21oi_1 _11916_ (.A1(net1350),
    .A2(net3989),
    .Y(_06846_),
    .B1(net3993));
 sg13g2_nand2_1 _11917_ (.Y(_06847_),
    .A(_06845_),
    .B(_06846_));
 sg13g2_a221oi_1 _11918_ (.B2(_05709_),
    .C1(net3862),
    .B1(net4106),
    .A1(_00275_),
    .Y(_06848_),
    .A2(_06635_));
 sg13g2_a22oi_1 _11919_ (.Y(_06849_),
    .B1(_06847_),
    .B2(_06848_),
    .A2(net3798),
    .A1(net2696));
 sg13g2_a21oi_1 _11920_ (.A1(_06787_),
    .A2(net4088),
    .Y(_06850_),
    .B1(net4229));
 sg13g2_a21oi_1 _11921_ (.A1(net2696),
    .A2(_06790_),
    .Y(_06851_),
    .B1(_06850_));
 sg13g2_a22oi_1 _11922_ (.Y(_00068_),
    .B1(_06851_),
    .B2(_06819_),
    .A2(_06849_),
    .A1(net3839));
 sg13g2_nand2_1 _11923_ (.Y(_06852_),
    .A(\soc_inst.gpio_bidir_oe [0]),
    .B(_06023_));
 sg13g2_o21ai_1 _11924_ (.B1(_06852_),
    .Y(uio_oe[7]),
    .A1(_05405_),
    .A2(_06023_));
 sg13g2_and2_1 _11925_ (.A(\soc_inst.gpio_bidir_out [0]),
    .B(_06023_),
    .X(uio_out[7]));
 sg13g2_nor2_1 _11926_ (.A(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .B(_05606_),
    .Y(_06853_));
 sg13g2_nor2_1 _11927_ (.A(_05572_),
    .B(\soc_inst.pwm_inst.channel_duty[1][3] ),
    .Y(_06854_));
 sg13g2_a22oi_1 _11928_ (.Y(_06855_),
    .B1(\soc_inst.pwm_inst.channel_duty[1][1] ),
    .B2(_05574_),
    .A2(\soc_inst.pwm_inst.channel_duty[1][0] ),
    .A1(_05575_));
 sg13g2_a221oi_1 _11929_ (.B2(\soc_inst.pwm_inst.channel_counter[1][2] ),
    .C1(_06855_),
    .B1(_05593_),
    .A1(\soc_inst.pwm_inst.channel_counter[1][1] ),
    .Y(_06856_),
    .A2(_05590_));
 sg13g2_a221oi_1 _11930_ (.B2(_05572_),
    .C1(_06856_),
    .B1(\soc_inst.pwm_inst.channel_duty[1][3] ),
    .A1(_05573_),
    .Y(_06857_),
    .A2(\soc_inst.pwm_inst.channel_duty[1][2] ));
 sg13g2_nand2b_1 _11931_ (.Y(_06858_),
    .B(\soc_inst.pwm_inst.channel_duty[1][4] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[1][4] ));
 sg13g2_o21ai_1 _11932_ (.B1(_06858_),
    .Y(_06859_),
    .A1(_06854_),
    .A2(_06857_));
 sg13g2_nand2b_1 _11933_ (.Y(_06860_),
    .B(\soc_inst.pwm_inst.channel_duty[1][5] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[1][5] ));
 sg13g2_a22oi_1 _11934_ (.Y(_06861_),
    .B1(_05597_),
    .B2(\soc_inst.pwm_inst.channel_counter[1][5] ),
    .A2(_05595_),
    .A1(\soc_inst.pwm_inst.channel_counter[1][4] ));
 sg13g2_o21ai_1 _11935_ (.B1(_06860_),
    .Y(_06862_),
    .A1(\soc_inst.pwm_inst.channel_counter[1][6] ),
    .A2(_05600_));
 sg13g2_a21oi_1 _11936_ (.A1(_06859_),
    .A2(_06861_),
    .Y(_06863_),
    .B1(_06862_));
 sg13g2_a221oi_1 _11937_ (.B2(\soc_inst.pwm_inst.channel_counter[1][7] ),
    .C1(_06863_),
    .B1(_05602_),
    .A1(\soc_inst.pwm_inst.channel_counter[1][6] ),
    .Y(_06864_),
    .A2(_05600_));
 sg13g2_nor2b_1 _11938_ (.A(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .B_N(\soc_inst.pwm_inst.channel_duty[1][9] ),
    .Y(_06865_));
 sg13g2_nor2_1 _11939_ (.A(\soc_inst.pwm_inst.channel_counter[1][7] ),
    .B(_05602_),
    .Y(_06866_));
 sg13g2_xor2_1 _11940_ (.B(\soc_inst.pwm_inst.channel_duty[1][8] ),
    .A(\soc_inst.pwm_inst.channel_counter[1][8] ),
    .X(_06867_));
 sg13g2_nor4_1 _11941_ (.A(_06864_),
    .B(_06865_),
    .C(_06866_),
    .D(_06867_),
    .Y(_06868_));
 sg13g2_nor3_1 _11942_ (.A(_05571_),
    .B(\soc_inst.pwm_inst.channel_duty[1][8] ),
    .C(_06865_),
    .Y(_06869_));
 sg13g2_nor2b_1 _11943_ (.A(\soc_inst.pwm_inst.channel_duty[1][9] ),
    .B_N(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .Y(_06870_));
 sg13g2_nor3_1 _11944_ (.A(_06868_),
    .B(_06869_),
    .C(_06870_),
    .Y(_06871_));
 sg13g2_a22oi_1 _11945_ (.Y(_06872_),
    .B1(_05608_),
    .B2(\soc_inst.pwm_inst.channel_counter[1][11] ),
    .A2(_05606_),
    .A1(\soc_inst.pwm_inst.channel_counter[1][10] ));
 sg13g2_o21ai_1 _11946_ (.B1(_06872_),
    .Y(_06873_),
    .A1(_06853_),
    .A2(_06871_));
 sg13g2_nor2b_1 _11947_ (.A(\soc_inst.pwm_inst.channel_duty[1][15] ),
    .B_N(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .Y(_06874_));
 sg13g2_nor2b_1 _11948_ (.A(\soc_inst.pwm_inst.channel_duty[1][14] ),
    .B_N(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .Y(_06875_));
 sg13g2_nor2_1 _11949_ (.A(_06874_),
    .B(_06875_),
    .Y(_06876_));
 sg13g2_nor2b_1 _11950_ (.A(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .B_N(\soc_inst.pwm_inst.channel_duty[1][15] ),
    .Y(_06877_));
 sg13g2_nor2b_1 _11951_ (.A(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .B_N(\soc_inst.pwm_inst.channel_duty[1][14] ),
    .Y(_06878_));
 sg13g2_nand2b_1 _11952_ (.Y(_06879_),
    .B(\soc_inst.pwm_inst.channel_duty[1][13] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[1][13] ));
 sg13g2_nor4_1 _11953_ (.A(_06874_),
    .B(_06875_),
    .C(_06877_),
    .D(_06878_),
    .Y(_06880_));
 sg13g2_nand2b_1 _11954_ (.Y(_06881_),
    .B(\soc_inst.pwm_inst.channel_counter[1][13] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[1][13] ));
 sg13g2_o21ai_1 _11955_ (.B1(_06881_),
    .Y(_06882_),
    .A1(_05569_),
    .A2(\soc_inst.pwm_inst.channel_duty[1][12] ));
 sg13g2_a221oi_1 _11956_ (.B2(_05569_),
    .C1(_06882_),
    .B1(\soc_inst.pwm_inst.channel_duty[1][12] ),
    .A1(_05570_),
    .Y(_06883_),
    .A2(\soc_inst.pwm_inst.channel_duty[1][11] ));
 sg13g2_nand4_1 _11957_ (.B(_06879_),
    .C(_06880_),
    .A(_06873_),
    .Y(_06884_),
    .D(_06883_));
 sg13g2_nand3_1 _11958_ (.B(_06880_),
    .C(_06882_),
    .A(_06879_),
    .Y(_06885_));
 sg13g2_or2_1 _11959_ (.X(_06886_),
    .B(_06877_),
    .A(_06876_));
 sg13g2_nand4_1 _11960_ (.B(_06884_),
    .C(_06885_),
    .A(\soc_inst.pwm_ena[1] ),
    .Y(_06887_),
    .D(_06886_));
 sg13g2_o21ai_1 _11961_ (.B1(_06887_),
    .Y(uo_out[7]),
    .A1(\soc_inst.pwm_ena[1] ),
    .A2(_05598_));
 sg13g2_nand2b_1 _11962_ (.Y(_06888_),
    .B(\soc_inst.pwm_inst.channel_duty[0][4] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[0][4] ));
 sg13g2_nand2b_1 _11963_ (.Y(_06889_),
    .B(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[0][3] ));
 sg13g2_a22oi_1 _11964_ (.Y(_06890_),
    .B1(\soc_inst.pwm_inst.channel_duty[0][1] ),
    .B2(_05581_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .A1(_05582_));
 sg13g2_a221oi_1 _11965_ (.B2(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .C1(_06890_),
    .B1(_05592_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .Y(_06891_),
    .A2(_05589_));
 sg13g2_nand2b_1 _11966_ (.Y(_06892_),
    .B(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[0][3] ));
 sg13g2_o21ai_1 _11967_ (.B1(_06892_),
    .Y(_06893_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .A2(_05592_));
 sg13g2_o21ai_1 _11968_ (.B1(_06889_),
    .Y(_06894_),
    .A1(_06891_),
    .A2(_06893_));
 sg13g2_nand2b_1 _11969_ (.Y(_06895_),
    .B(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[0][4] ));
 sg13g2_o21ai_1 _11970_ (.B1(_06895_),
    .Y(_06896_),
    .A1(_05580_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][5] ));
 sg13g2_a21oi_1 _11971_ (.A1(_06888_),
    .A2(_06894_),
    .Y(_06897_),
    .B1(_06896_));
 sg13g2_a221oi_1 _11972_ (.B2(_05579_),
    .C1(_06897_),
    .B1(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .A1(_05580_),
    .Y(_06898_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][5] ));
 sg13g2_a221oi_1 _11973_ (.B2(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .C1(_06898_),
    .B1(_05601_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .Y(_06899_),
    .A2(_05599_));
 sg13g2_a22oi_1 _11974_ (.Y(_06900_),
    .B1(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .B2(_05577_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .A1(_05578_));
 sg13g2_o21ai_1 _11975_ (.B1(_06900_),
    .Y(_06901_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .A2(_05601_));
 sg13g2_a22oi_1 _11976_ (.Y(_06902_),
    .B1(_05605_),
    .B2(net5127),
    .A2(_05604_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][8] ));
 sg13g2_o21ai_1 _11977_ (.B1(_06902_),
    .Y(_06903_),
    .A1(_06899_),
    .A2(_06901_));
 sg13g2_nor3_1 _11978_ (.A(net5127),
    .B(_05578_),
    .C(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .Y(_06904_));
 sg13g2_nor2_1 _11979_ (.A(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .B(_05607_),
    .Y(_06905_));
 sg13g2_a221oi_1 _11980_ (.B2(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .C1(_06905_),
    .B1(_06904_),
    .A1(_05576_),
    .Y(_06906_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][10] ));
 sg13g2_nor2_1 _11981_ (.A(_05576_),
    .B(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .Y(_06907_));
 sg13g2_a221oi_1 _11982_ (.B2(_06906_),
    .C1(_06907_),
    .B1(_06903_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .Y(_06908_),
    .A2(_05607_));
 sg13g2_nand2b_1 _11983_ (.Y(_06909_),
    .B(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[0][15] ));
 sg13g2_nand2b_1 _11984_ (.Y(_06910_),
    .B(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[0][15] ));
 sg13g2_nor2b_1 _11985_ (.A(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .B_N(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .Y(_06911_));
 sg13g2_xnor2_1 _11986_ (.Y(_06912_),
    .A(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .B(\soc_inst.pwm_inst.channel_duty[0][14] ));
 sg13g2_nand3_1 _11987_ (.B(_06910_),
    .C(_06912_),
    .A(_06909_),
    .Y(_06913_));
 sg13g2_nand2_1 _11988_ (.Y(_06914_),
    .A(_06905_),
    .B(_06907_));
 sg13g2_a22oi_1 _11989_ (.Y(_06915_),
    .B1(_05610_),
    .B2(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .A2(_05609_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][12] ));
 sg13g2_nor2_1 _11990_ (.A(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .B(_05610_),
    .Y(_06916_));
 sg13g2_nand2b_1 _11991_ (.Y(_06917_),
    .B(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[0][13] ));
 sg13g2_o21ai_1 _11992_ (.B1(_06917_),
    .Y(_06918_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .A2(_05609_));
 sg13g2_nand2_1 _11993_ (.Y(_06919_),
    .A(_06914_),
    .B(_06915_));
 sg13g2_or4_1 _11994_ (.A(_06908_),
    .B(_06913_),
    .C(_06918_),
    .D(_06919_),
    .X(_06920_));
 sg13g2_nor3_1 _11995_ (.A(_06913_),
    .B(_06915_),
    .C(_06916_),
    .Y(_06921_));
 sg13g2_a21oi_1 _11996_ (.A1(_06910_),
    .A2(_06911_),
    .Y(_06922_),
    .B1(_06921_));
 sg13g2_nand4_1 _11997_ (.B(_06909_),
    .C(_06920_),
    .A(\soc_inst.pwm_ena[0] ),
    .Y(_06923_),
    .D(_06922_));
 sg13g2_o21ai_1 _11998_ (.B1(_06923_),
    .Y(uo_out[6]),
    .A1(\soc_inst.pwm_ena[0] ),
    .A2(_05596_));
 sg13g2_nor2_1 _11999_ (.A(\soc_inst.spi_ena ),
    .B(\soc_inst.gpio_inst.gpio_out[3] ),
    .Y(_06924_));
 sg13g2_a21oi_2 _12000_ (.B1(_06924_),
    .Y(uo_out[5]),
    .A2(_05784_),
    .A1(\soc_inst.spi_ena ));
 sg13g2_mux2_1 _12001_ (.A0(\soc_inst.gpio_inst.gpio_out[2] ),
    .A1(\soc_inst.spi_inst.spi_sclk ),
    .S(\soc_inst.spi_ena ),
    .X(uo_out[4]));
 sg13g2_nand2_1 _12002_ (.Y(_06925_),
    .A(\soc_inst.gpio_inst.gpio_out[0] ),
    .B(_06023_));
 sg13g2_o21ai_1 _12003_ (.B1(_06925_),
    .Y(uo_out[2]),
    .A1(_00229_),
    .A2(_06023_));
 sg13g2_nand2_1 _12004_ (.Y(_06926_),
    .A(net5035),
    .B(_06414_));
 sg13g2_and3_1 _12005_ (.X(_06927_),
    .A(net5115),
    .B(net5118),
    .C(_06020_));
 sg13g2_nand3_1 _12006_ (.B(net5117),
    .C(_06020_),
    .A(net5115),
    .Y(_06928_));
 sg13g2_a21o_1 _12007_ (.A2(net2404),
    .A1(net1558),
    .B1(_06928_),
    .X(_06929_));
 sg13g2_or4_1 _12008_ (.A(net5115),
    .B(net5117),
    .C(_06418_),
    .D(net4275),
    .X(_06930_));
 sg13g2_o21ai_1 _12009_ (.B1(_06930_),
    .Y(_06931_),
    .A1(net4274),
    .A2(_06928_));
 sg13g2_a22oi_1 _12010_ (.Y(_10277_[0]),
    .B1(_06929_),
    .B2(_06931_),
    .A2(_06926_),
    .A1(_05864_));
 sg13g2_nand2_1 _12011_ (.Y(_06932_),
    .A(_05468_),
    .B(net343));
 sg13g2_nand2_1 _12012_ (.Y(_06933_),
    .A(_00218_),
    .B(_00217_));
 sg13g2_nand3_1 _12013_ (.B(_00218_),
    .C(_00217_),
    .A(_00219_),
    .Y(_06934_));
 sg13g2_nor2_1 _12014_ (.A(_05406_),
    .B(_06934_),
    .Y(_06935_));
 sg13g2_nand2_1 _12015_ (.Y(_06936_),
    .A(_00221_),
    .B(_06935_));
 sg13g2_nor2_1 _12016_ (.A(\soc_inst.spi_inst.clock_divider[5] ),
    .B(_06936_),
    .Y(_06937_));
 sg13g2_nor3_1 _12017_ (.A(\soc_inst.spi_inst.bit_counter[0] ),
    .B(\soc_inst.spi_inst.bit_counter[1] ),
    .C(\soc_inst.spi_inst.bit_counter[2] ),
    .Y(_06938_));
 sg13g2_nor2b_1 _12018_ (.A(net5125),
    .B_N(\soc_inst.spi_inst.len_sel[0] ),
    .Y(_06939_));
 sg13g2_nand2b_2 _12019_ (.Y(_06940_),
    .B(\soc_inst.spi_inst.len_sel[0] ),
    .A_N(net5126));
 sg13g2_nand2_1 _12020_ (.Y(_06941_),
    .A(\soc_inst.spi_inst.bit_counter[4] ),
    .B(_06940_));
 sg13g2_nor2_1 _12021_ (.A(\soc_inst.spi_inst.bit_counter[4] ),
    .B(net5126),
    .Y(_06942_));
 sg13g2_o21ai_1 _12022_ (.B1(\soc_inst.spi_inst.bit_counter[3] ),
    .Y(_06943_),
    .A1(\soc_inst.spi_inst.bit_counter[4] ),
    .A2(net5126));
 sg13g2_o21ai_1 _12023_ (.B1(_06942_),
    .Y(_06944_),
    .A1(_05567_),
    .A2(\soc_inst.spi_inst.len_sel[0] ));
 sg13g2_nand4_1 _12024_ (.B(_06941_),
    .C(_06943_),
    .A(_06938_),
    .Y(_06945_),
    .D(_06944_));
 sg13g2_a21oi_1 _12025_ (.A1(_06309_),
    .A2(_06935_),
    .Y(_06946_),
    .B1(_06945_));
 sg13g2_o21ai_1 _12026_ (.B1(_06946_),
    .Y(_06947_),
    .A1(_06309_),
    .A2(_06935_));
 sg13g2_a21oi_1 _12027_ (.A1(_06310_),
    .A2(_06937_),
    .Y(_06948_),
    .B1(_06947_));
 sg13g2_o21ai_1 _12028_ (.B1(_06948_),
    .Y(_06949_),
    .A1(_06310_),
    .A2(_06937_));
 sg13g2_nor3_1 _12029_ (.A(\soc_inst.spi_inst.clock_divider[5] ),
    .B(\soc_inst.spi_inst.clock_divider[6] ),
    .C(_06936_),
    .Y(_06950_));
 sg13g2_and2_1 _12030_ (.A(_06314_),
    .B(_06950_),
    .X(_06951_));
 sg13g2_nor3_1 _12031_ (.A(\soc_inst.spi_inst.clk_counter[7] ),
    .B(_05502_),
    .C(_06950_),
    .Y(_06952_));
 sg13g2_xnor2_1 _12032_ (.Y(_06953_),
    .A(_06315_),
    .B(_06936_));
 sg13g2_xor2_1 _12033_ (.B(_06934_),
    .A(_06311_),
    .X(_06954_));
 sg13g2_a21oi_1 _12034_ (.A1(_00217_),
    .A2(\soc_inst.spi_inst.clk_counter[0] ),
    .Y(_06955_),
    .B1(_06312_));
 sg13g2_xnor2_1 _12035_ (.Y(_06956_),
    .A(_06316_),
    .B(_06933_));
 sg13g2_a21oi_1 _12036_ (.A1(\soc_inst.spi_inst.clk_counter[7] ),
    .A2(_05502_),
    .Y(_06957_),
    .B1(net4717));
 sg13g2_xnor2_1 _12037_ (.Y(_06958_),
    .A(\soc_inst.spi_inst.bit_counter[5] ),
    .B(net5126));
 sg13g2_nand4_1 _12038_ (.B(_06956_),
    .C(_06957_),
    .A(_06313_),
    .Y(_06959_),
    .D(_06958_));
 sg13g2_or4_1 _12039_ (.A(_06953_),
    .B(_06954_),
    .C(_06955_),
    .D(_06959_),
    .X(_06960_));
 sg13g2_or4_1 _12040_ (.A(_06949_),
    .B(_06951_),
    .C(_06952_),
    .D(_06960_),
    .X(_06961_));
 sg13g2_o21ai_1 _12041_ (.B1(_06961_),
    .Y(\soc_inst.spi_inst.next_state[0] ),
    .A1(\soc_inst.spi_inst.state[0] ),
    .A2(net344));
 sg13g2_and2_1 _12042_ (.A(_00123_),
    .B(_06961_),
    .X(_10279_[0]));
 sg13g2_a21oi_1 _12043_ (.A1(net5048),
    .A2(_06414_),
    .Y(_06962_),
    .B1(net1558));
 sg13g2_or3_1 _12044_ (.A(net1558),
    .B(net4274),
    .C(_06928_),
    .X(_06963_));
 sg13g2_a21oi_1 _12045_ (.A1(_06931_),
    .A2(_06963_),
    .Y(_10278_[0]),
    .B1(_06962_));
 sg13g2_nor2_2 _12046_ (.A(_06021_),
    .B(_06440_),
    .Y(_06964_));
 sg13g2_nand2_1 _12047_ (.Y(_06965_),
    .A(net4276),
    .B(_06964_));
 sg13g2_o21ai_1 _12048_ (.B1(_06965_),
    .Y(_06966_),
    .A1(\soc_inst.i2c_inst.start_pending ),
    .A2(\soc_inst.i2c_ena ));
 sg13g2_a21oi_1 _12049_ (.A1(net2661),
    .A2(_06430_),
    .Y(_06967_),
    .B1(_06928_));
 sg13g2_nand2_1 _12050_ (.Y(_06968_),
    .A(net5128),
    .B(_06964_));
 sg13g2_nor2_1 _12051_ (.A(_06021_),
    .B(_06416_),
    .Y(_06969_));
 sg13g2_nor4_1 _12052_ (.A(\soc_inst.i2c_inst.clk_cnt[4] ),
    .B(\soc_inst.i2c_inst.clk_cnt[5] ),
    .C(\soc_inst.i2c_inst.clk_cnt[6] ),
    .D(\soc_inst.i2c_inst.clk_cnt[7] ),
    .Y(_06970_));
 sg13g2_nor4_1 _12053_ (.A(\soc_inst.i2c_inst.clk_cnt[0] ),
    .B(\soc_inst.i2c_inst.clk_cnt[1] ),
    .C(\soc_inst.i2c_inst.clk_cnt[2] ),
    .D(\soc_inst.i2c_inst.clk_cnt[3] ),
    .Y(_06971_));
 sg13g2_and2_1 _12054_ (.A(_06970_),
    .B(_06971_),
    .X(_06972_));
 sg13g2_inv_1 _12055_ (.Y(_06973_),
    .A(_06972_));
 sg13g2_nand3b_1 _12056_ (.B(\soc_inst.i2c_inst.state[1] ),
    .C(net5120),
    .Y(_06974_),
    .A_N(net5118));
 sg13g2_or2_1 _12057_ (.X(_06975_),
    .B(_06974_),
    .A(net5115));
 sg13g2_nor3_1 _12058_ (.A(_05473_),
    .B(_06973_),
    .C(_06975_),
    .Y(_06976_));
 sg13g2_o21ai_1 _12059_ (.B1(_06968_),
    .Y(_06977_),
    .A1(_06969_),
    .A2(_06976_));
 sg13g2_nor3_2 _12060_ (.A(_06966_),
    .B(_06967_),
    .C(_06977_),
    .Y(_06978_));
 sg13g2_o21ai_1 _12061_ (.B1(_06446_),
    .Y(_06979_),
    .A1(net669),
    .A2(net4008));
 sg13g2_and3_1 _12062_ (.X(_06980_),
    .A(net1558),
    .B(_06440_),
    .C(_06969_));
 sg13g2_and2_1 _12063_ (.A(net2828),
    .B(_06980_),
    .X(_06981_));
 sg13g2_a22oi_1 _12064_ (.Y(_06982_),
    .B1(_06981_),
    .B2(net4202),
    .A2(_06976_),
    .A1(net13));
 sg13g2_o21ai_1 _12065_ (.B1(_06982_),
    .Y(_02148_),
    .A1(_06978_),
    .A2(_06979_));
 sg13g2_o21ai_1 _12066_ (.B1(_06450_),
    .Y(_06983_),
    .A1(net545),
    .A2(net4006));
 sg13g2_o21ai_1 _12067_ (.B1(\soc_inst.i2c_ena ),
    .Y(_06984_),
    .A1(net4276),
    .A2(_06928_));
 sg13g2_and2_1 _12068_ (.A(\soc_inst.i2c_inst.start_pending ),
    .B(_06984_),
    .X(_06985_));
 sg13g2_nor4_1 _12069_ (.A(net5128),
    .B(_06021_),
    .C(net4274),
    .D(_06440_),
    .Y(_06986_));
 sg13g2_or2_1 _12070_ (.X(_06987_),
    .B(_06986_),
    .A(_06976_));
 sg13g2_a22oi_1 _12071_ (.Y(_06988_),
    .B1(_06987_),
    .B2(net669),
    .A2(_06985_),
    .A1(net2146));
 sg13g2_o21ai_1 _12072_ (.B1(net2147),
    .Y(_02149_),
    .A1(_06978_),
    .A2(_06983_));
 sg13g2_nor2_1 _12073_ (.A(net1523),
    .B(net4006),
    .Y(_06989_));
 sg13g2_nor3_1 _12074_ (.A(_06454_),
    .B(_06978_),
    .C(_06989_),
    .Y(_06990_));
 sg13g2_a221oi_1 _12075_ (.B2(net545),
    .C1(_06990_),
    .B1(_06987_),
    .A1(net2712),
    .Y(_06991_),
    .A2(_06985_));
 sg13g2_inv_1 _12076_ (.Y(_02150_),
    .A(_06991_));
 sg13g2_o21ai_1 _12077_ (.B1(_06456_),
    .Y(_06992_),
    .A1(net652),
    .A2(net4007));
 sg13g2_a22oi_1 _12078_ (.Y(_06993_),
    .B1(_06987_),
    .B2(net1523),
    .A2(_06985_),
    .A1(net2054));
 sg13g2_o21ai_1 _12079_ (.B1(net2055),
    .Y(_02151_),
    .A1(_06978_),
    .A2(_06992_));
 sg13g2_o21ai_1 _12080_ (.B1(_06459_),
    .Y(_06994_),
    .A1(net492),
    .A2(net4006));
 sg13g2_a22oi_1 _12081_ (.Y(_06995_),
    .B1(_06987_),
    .B2(net652),
    .A2(_06985_),
    .A1(net2308));
 sg13g2_o21ai_1 _12082_ (.B1(net2309),
    .Y(_02152_),
    .A1(_06978_),
    .A2(_06994_));
 sg13g2_o21ai_1 _12083_ (.B1(_06463_),
    .Y(_06996_),
    .A1(net536),
    .A2(net4006));
 sg13g2_a22oi_1 _12084_ (.Y(_06997_),
    .B1(_06987_),
    .B2(net492),
    .A2(_06985_),
    .A1(net2155));
 sg13g2_o21ai_1 _12085_ (.B1(net2156),
    .Y(_02153_),
    .A1(_06978_),
    .A2(_06996_));
 sg13g2_nor2_1 _12086_ (.A(net1692),
    .B(net4006),
    .Y(_06998_));
 sg13g2_nor3_1 _12087_ (.A(_06467_),
    .B(_06978_),
    .C(_06998_),
    .Y(_06999_));
 sg13g2_a221oi_1 _12088_ (.B2(net536),
    .C1(_06999_),
    .B1(_06987_),
    .A1(net2645),
    .Y(_07000_),
    .A2(_06985_));
 sg13g2_inv_1 _12089_ (.Y(_02154_),
    .A(_07000_));
 sg13g2_nor2_1 _12090_ (.A(net1183),
    .B(net4008),
    .Y(_07001_));
 sg13g2_nor3_1 _12091_ (.A(_06470_),
    .B(_06978_),
    .C(_07001_),
    .Y(_07002_));
 sg13g2_a221oi_1 _12092_ (.B2(net1692),
    .C1(_07002_),
    .B1(_06987_),
    .A1(net1790),
    .Y(_07003_),
    .A2(_06985_));
 sg13g2_inv_1 _12093_ (.Y(_02155_),
    .A(_07003_));
 sg13g2_and2_1 _12094_ (.A(_05882_),
    .B(_05892_),
    .X(_07004_));
 sg13g2_nand4_1 _12095_ (.B(net4785),
    .C(net4206),
    .A(net5041),
    .Y(_07005_),
    .D(_07004_));
 sg13g2_nor3_1 _12096_ (.A(net938),
    .B(net1120),
    .C(_06117_),
    .Y(_07006_));
 sg13g2_nand2b_2 _12097_ (.Y(_07007_),
    .B(_07006_),
    .A_N(_06121_));
 sg13g2_nor4_1 _12098_ (.A(net655),
    .B(net1019),
    .C(net620),
    .D(net605),
    .Y(_07008_));
 sg13g2_nor4_1 _12099_ (.A(net1276),
    .B(net1299),
    .C(net1991),
    .D(net597),
    .Y(_07009_));
 sg13g2_and2_1 _12100_ (.A(_07008_),
    .B(_07009_),
    .X(_07010_));
 sg13g2_nand2_2 _12101_ (.Y(_07011_),
    .A(net4786),
    .B(_05901_));
 sg13g2_o21ai_1 _12102_ (.B1(_07010_),
    .Y(_07012_),
    .A1(_06298_),
    .A2(_07011_));
 sg13g2_o21ai_1 _12103_ (.B1(_07005_),
    .Y(_00166_),
    .A1(_07007_),
    .A2(_07012_));
 sg13g2_nand4_1 _12104_ (.B(_05891_),
    .C(_05892_),
    .A(net4785),
    .Y(_07013_),
    .D(net4206));
 sg13g2_nand3_1 _12105_ (.B(_06110_),
    .C(_07006_),
    .A(net1584),
    .Y(_07014_));
 sg13g2_nand2b_1 _12106_ (.Y(_07015_),
    .B(_07014_),
    .A_N(net2933));
 sg13g2_mux2_1 _12107_ (.A0(net5047),
    .A1(_07015_),
    .S(_07013_),
    .X(_00167_));
 sg13g2_nand3_1 _12108_ (.B(net2687),
    .C(net4259),
    .A(net5049),
    .Y(_07016_));
 sg13g2_or3_1 _12109_ (.A(net2913),
    .B(_06300_),
    .C(_07016_),
    .X(_07017_));
 sg13g2_inv_2 _12110_ (.Y(_00133_),
    .A(_07017_));
 sg13g2_nor3_1 _12111_ (.A(net5121),
    .B(_05506_),
    .C(_06139_),
    .Y(_00000_));
 sg13g2_nor2b_1 _12112_ (.A(net97),
    .B_N(\soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ),
    .Y(_00090_));
 sg13g2_xor2_1 _12113_ (.B(net761),
    .A(net556),
    .X(_00180_));
 sg13g2_nand3_1 _12114_ (.B(net761),
    .C(net2898),
    .A(net556),
    .Y(_07018_));
 sg13g2_a21o_1 _12115_ (.A2(net761),
    .A1(net556),
    .B1(net2898),
    .X(_07019_));
 sg13g2_and2_1 _12116_ (.A(_07018_),
    .B(_07019_),
    .X(_00191_));
 sg13g2_and4_1 _12117_ (.A(net556),
    .B(net761),
    .C(net967),
    .D(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .X(_07020_));
 sg13g2_xnor2_1 _12118_ (.Y(_00202_),
    .A(net967),
    .B(_07018_));
 sg13g2_xor2_1 _12119_ (.B(_07020_),
    .A(net1660),
    .X(_00211_));
 sg13g2_nand3_1 _12120_ (.B(net1660),
    .C(_07020_),
    .A(net2925),
    .Y(_07021_));
 sg13g2_a21o_1 _12121_ (.A2(_07020_),
    .A1(net1660),
    .B1(net2925),
    .X(_07022_));
 sg13g2_and2_1 _12122_ (.A(_07021_),
    .B(_07022_),
    .X(_00212_));
 sg13g2_nand4_1 _12123_ (.B(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .C(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .A(net826),
    .Y(_07023_),
    .D(_07020_));
 sg13g2_xnor2_1 _12124_ (.Y(_00213_),
    .A(net826),
    .B(_07021_));
 sg13g2_nor2_2 _12125_ (.A(_05509_),
    .B(_07023_),
    .Y(_07024_));
 sg13g2_xnor2_1 _12126_ (.Y(_00214_),
    .A(net1262),
    .B(_07023_));
 sg13g2_xor2_1 _12127_ (.B(_07024_),
    .A(net884),
    .X(_00215_));
 sg13g2_nand3_1 _12128_ (.B(net884),
    .C(_07024_),
    .A(net2885),
    .Y(_07025_));
 sg13g2_a21o_1 _12129_ (.A2(_07024_),
    .A1(net884),
    .B1(net2885),
    .X(_07026_));
 sg13g2_and2_1 _12130_ (.A(_07025_),
    .B(net2886),
    .X(_00216_));
 sg13g2_and4_1 _12131_ (.A(net645),
    .B(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .C(net884),
    .D(_07024_),
    .X(_07027_));
 sg13g2_xnor2_1 _12132_ (.Y(_00170_),
    .A(net645),
    .B(_07025_));
 sg13g2_xor2_1 _12133_ (.B(_07027_),
    .A(net1168),
    .X(_00171_));
 sg13g2_and3_2 _12134_ (.X(_07028_),
    .A(net2192),
    .B(net1168),
    .C(_07027_));
 sg13g2_a21oi_1 _12135_ (.A1(net1168),
    .A2(_07027_),
    .Y(_07029_),
    .B1(net2192));
 sg13g2_nor2_1 _12136_ (.A(_07028_),
    .B(net2193),
    .Y(_00172_));
 sg13g2_and2_1 _12137_ (.A(net1611),
    .B(_07028_),
    .X(_07030_));
 sg13g2_xor2_1 _12138_ (.B(_07028_),
    .A(net1611),
    .X(_00173_));
 sg13g2_xor2_1 _12139_ (.B(_07030_),
    .A(net1833),
    .X(_00174_));
 sg13g2_nand4_1 _12140_ (.B(net1833),
    .C(net1611),
    .A(net2928),
    .Y(_07031_),
    .D(_07028_));
 sg13g2_a21o_1 _12141_ (.A2(_07030_),
    .A1(net1833),
    .B1(net2928),
    .X(_07032_));
 sg13g2_and2_1 _12142_ (.A(_07031_),
    .B(_07032_),
    .X(_00175_));
 sg13g2_nand4_1 _12143_ (.B(net1833),
    .C(net2424),
    .A(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .Y(_07033_),
    .D(_07030_));
 sg13g2_xnor2_1 _12144_ (.Y(_00176_),
    .A(net2424),
    .B(_07031_));
 sg13g2_nand2_2 _12145_ (.Y(_07034_),
    .A(net2438),
    .B(net2424));
 sg13g2_nor2_1 _12146_ (.A(_07031_),
    .B(_07034_),
    .Y(_07035_));
 sg13g2_xnor2_1 _12147_ (.Y(_00177_),
    .A(net2438),
    .B(_07033_));
 sg13g2_xor2_1 _12148_ (.B(_07035_),
    .A(net2126),
    .X(_00178_));
 sg13g2_a21oi_1 _12149_ (.A1(net2126),
    .A2(_07035_),
    .Y(_07036_),
    .B1(net2602));
 sg13g2_nand2_1 _12150_ (.Y(_07037_),
    .A(net2602),
    .B(net2126));
 sg13g2_nor3_2 _12151_ (.A(_07031_),
    .B(_07034_),
    .C(_07037_),
    .Y(_07038_));
 sg13g2_nor2_1 _12152_ (.A(_07036_),
    .B(_07038_),
    .Y(_00179_));
 sg13g2_xor2_1 _12153_ (.B(_07038_),
    .A(net2419),
    .X(_00181_));
 sg13g2_a21oi_1 _12154_ (.A1(net2419),
    .A2(_07038_),
    .Y(_07039_),
    .B1(net2698));
 sg13g2_and3_2 _12155_ (.X(_07040_),
    .A(net2698),
    .B(net2419),
    .C(_07038_));
 sg13g2_nor2_1 _12156_ (.A(_07039_),
    .B(_07040_),
    .Y(_00182_));
 sg13g2_xor2_1 _12157_ (.B(_07040_),
    .A(net1527),
    .X(_00183_));
 sg13g2_a21oi_1 _12158_ (.A1(net1527),
    .A2(_07040_),
    .Y(_07041_),
    .B1(net2540));
 sg13g2_nand4_1 _12159_ (.B(net1527),
    .C(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .A(net2540),
    .Y(_07042_),
    .D(net2419));
 sg13g2_nor4_2 _12160_ (.A(_07031_),
    .B(_07034_),
    .C(_07037_),
    .Y(_07043_),
    .D(_07042_));
 sg13g2_nor2_1 _12161_ (.A(net2541),
    .B(_07043_),
    .Y(_00184_));
 sg13g2_xor2_1 _12162_ (.B(_07043_),
    .A(net2227),
    .X(_00185_));
 sg13g2_a21oi_1 _12163_ (.A1(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .A2(_07043_),
    .Y(_07044_),
    .B1(net2218));
 sg13g2_and3_2 _12164_ (.X(_07045_),
    .A(net2218),
    .B(net2227),
    .C(_07043_));
 sg13g2_nor2_1 _12165_ (.A(net2219),
    .B(_07045_),
    .Y(_00186_));
 sg13g2_nand2_1 _12166_ (.Y(_07046_),
    .A(net1656),
    .B(_07045_));
 sg13g2_xor2_1 _12167_ (.B(_07045_),
    .A(net1656),
    .X(_00187_));
 sg13g2_xnor2_1 _12168_ (.Y(_00188_),
    .A(net2266),
    .B(_07046_));
 sg13g2_nand3_1 _12169_ (.B(net1656),
    .C(_07045_),
    .A(net2266),
    .Y(_07047_));
 sg13g2_or2_1 _12170_ (.X(_07048_),
    .B(_07047_),
    .A(_05513_));
 sg13g2_xnor2_1 _12171_ (.Y(_00189_),
    .A(net1772),
    .B(_07047_));
 sg13g2_nor3_2 _12172_ (.A(_05512_),
    .B(_05513_),
    .C(_07047_),
    .Y(_07049_));
 sg13g2_a21oi_1 _12173_ (.A1(_05512_),
    .A2(_07048_),
    .Y(_00190_),
    .B1(_07049_));
 sg13g2_nand2_1 _12174_ (.Y(_07050_),
    .A(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .B(_07049_));
 sg13g2_xor2_1 _12175_ (.B(_07049_),
    .A(net2049),
    .X(_00192_));
 sg13g2_xnor2_1 _12176_ (.Y(_00193_),
    .A(net1900),
    .B(_07050_));
 sg13g2_and3_2 _12177_ (.X(_07051_),
    .A(net1900),
    .B(net2049),
    .C(_07049_));
 sg13g2_xnor2_1 _12178_ (.Y(_00194_),
    .A(_05516_),
    .B(_07051_));
 sg13g2_a21oi_1 _12179_ (.A1(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .A2(_07051_),
    .Y(_07052_),
    .B1(net1892));
 sg13g2_nand3_1 _12180_ (.B(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .C(_07051_),
    .A(net1892),
    .Y(_07053_));
 sg13g2_nor2b_1 _12181_ (.A(net1893),
    .B_N(_07053_),
    .Y(_00195_));
 sg13g2_and4_1 _12182_ (.A(net2587),
    .B(net1892),
    .C(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .D(_07051_),
    .X(_07054_));
 sg13g2_a21oi_1 _12183_ (.A1(_05515_),
    .A2(_07053_),
    .Y(_00196_),
    .B1(_07054_));
 sg13g2_nand2_1 _12184_ (.Y(_07055_),
    .A(net1244),
    .B(_07054_));
 sg13g2_inv_1 _12185_ (.Y(_07056_),
    .A(_07055_));
 sg13g2_xor2_1 _12186_ (.B(_07054_),
    .A(net1244),
    .X(_00197_));
 sg13g2_xnor2_1 _12187_ (.Y(_00198_),
    .A(net1715),
    .B(_07055_));
 sg13g2_a21oi_1 _12188_ (.A1(net1715),
    .A2(_07056_),
    .Y(_07057_),
    .B1(net1855));
 sg13g2_and4_1 _12189_ (.A(net1855),
    .B(net1715),
    .C(net1244),
    .D(_07054_),
    .X(_07058_));
 sg13g2_nor2_1 _12190_ (.A(_07057_),
    .B(_07058_),
    .Y(_00199_));
 sg13g2_and2_1 _12191_ (.A(net793),
    .B(_07058_),
    .X(_07059_));
 sg13g2_xor2_1 _12192_ (.B(_07058_),
    .A(net793),
    .X(_00200_));
 sg13g2_xor2_1 _12193_ (.B(_07059_),
    .A(net1653),
    .X(_00201_));
 sg13g2_a21oi_1 _12194_ (.A1(net1653),
    .A2(_07059_),
    .Y(_07060_),
    .B1(net1756));
 sg13g2_nand3_1 _12195_ (.B(net1653),
    .C(_07059_),
    .A(net1756),
    .Y(_07061_));
 sg13g2_nor2b_1 _12196_ (.A(_07060_),
    .B_N(_07061_),
    .Y(_00203_));
 sg13g2_and4_1 _12197_ (.A(net1932),
    .B(net1756),
    .C(net1653),
    .D(_07059_),
    .X(_07062_));
 sg13g2_a21oi_1 _12198_ (.A1(_05514_),
    .A2(_07061_),
    .Y(_00204_),
    .B1(_07062_));
 sg13g2_xor2_1 _12199_ (.B(_07062_),
    .A(net724),
    .X(_00205_));
 sg13g2_and3_2 _12200_ (.X(_07063_),
    .A(net1025),
    .B(net724),
    .C(_07062_));
 sg13g2_a21oi_1 _12201_ (.A1(net724),
    .A2(_07062_),
    .Y(_07064_),
    .B1(net1025));
 sg13g2_nor2_1 _12202_ (.A(_07063_),
    .B(net1026),
    .Y(_00206_));
 sg13g2_and2_1 _12203_ (.A(net1093),
    .B(_07063_),
    .X(_07065_));
 sg13g2_xor2_1 _12204_ (.B(_07063_),
    .A(net1093),
    .X(_00207_));
 sg13g2_xor2_1 _12205_ (.B(_07065_),
    .A(net1407),
    .X(_00208_));
 sg13g2_nand3_1 _12206_ (.B(net1407),
    .C(_07065_),
    .A(net2916),
    .Y(_07066_));
 sg13g2_a21o_1 _12207_ (.A2(_07065_),
    .A1(net1407),
    .B1(net2916),
    .X(_07067_));
 sg13g2_and2_1 _12208_ (.A(_07066_),
    .B(_07067_),
    .X(_00209_));
 sg13g2_xnor2_1 _12209_ (.Y(_00210_),
    .A(net694),
    .B(_07066_));
 sg13g2_nor2b_1 _12210_ (.A(net5122),
    .B_N(net486),
    .Y(_00001_));
 sg13g2_or2_1 _12211_ (.X(_07068_),
    .B(_06141_),
    .A(_05496_));
 sg13g2_nor2_1 _12212_ (.A(net5122),
    .B(_07068_),
    .Y(_00005_));
 sg13g2_nor4_1 _12213_ (.A(net5124),
    .B(net5076),
    .C(_05495_),
    .D(_06146_),
    .Y(_00004_));
 sg13g2_nor3_1 _12214_ (.A(net5121),
    .B(_05498_),
    .C(_06152_),
    .Y(_00003_));
 sg13g2_nor3_1 _12215_ (.A(net91),
    .B(net4278),
    .C(_06050_),
    .Y(_00002_));
 sg13g2_and4_1 _12216_ (.A(net5045),
    .B(net4786),
    .C(net4259),
    .D(_07004_),
    .X(_00168_));
 sg13g2_or2_1 _12217_ (.X(_07069_),
    .B(_06523_),
    .A(net4269));
 sg13g2_nor2_2 _12218_ (.A(_06526_),
    .B(_07069_),
    .Y(_07070_));
 sg13g2_mux2_1 _12219_ (.A0(net2118),
    .A1(net5047),
    .S(_07070_),
    .X(_00333_));
 sg13g2_mux2_1 _12220_ (.A0(net1728),
    .A1(net5044),
    .S(net3987),
    .X(_00334_));
 sg13g2_mux2_1 _12221_ (.A0(net1939),
    .A1(net5041),
    .S(net3987),
    .X(_00335_));
 sg13g2_mux2_1 _12222_ (.A0(net2292),
    .A1(net5038),
    .S(net3987),
    .X(_00336_));
 sg13g2_mux2_1 _12223_ (.A0(net1744),
    .A1(net5035),
    .S(net3986),
    .X(_00337_));
 sg13g2_mux2_1 _12224_ (.A0(net1966),
    .A1(net5033),
    .S(net3986),
    .X(_00338_));
 sg13g2_mux2_1 _12225_ (.A0(net1867),
    .A1(net5032),
    .S(net3987),
    .X(_00339_));
 sg13g2_mux2_1 _12226_ (.A0(net1709),
    .A1(net5028),
    .S(net3986),
    .X(_00340_));
 sg13g2_mux2_1 _12227_ (.A0(net2210),
    .A1(net5026),
    .S(net3986),
    .X(_00341_));
 sg13g2_mux2_1 _12228_ (.A0(net2415),
    .A1(net5024),
    .S(net3986),
    .X(_00342_));
 sg13g2_mux2_1 _12229_ (.A0(net1188),
    .A1(net5023),
    .S(net3986),
    .X(_00343_));
 sg13g2_mux2_1 _12230_ (.A0(net2202),
    .A1(net5022),
    .S(net3986),
    .X(_00344_));
 sg13g2_mux2_1 _12231_ (.A0(net2179),
    .A1(net5021),
    .S(net3986),
    .X(_00345_));
 sg13g2_mux2_1 _12232_ (.A0(net2313),
    .A1(net5020),
    .S(net3987),
    .X(_00346_));
 sg13g2_mux2_1 _12233_ (.A0(net2407),
    .A1(net5019),
    .S(net3987),
    .X(_00347_));
 sg13g2_mux2_1 _12234_ (.A0(net2197),
    .A1(net5018),
    .S(net3987),
    .X(_00348_));
 sg13g2_a21oi_1 _12235_ (.A1(\soc_inst.spi_inst.cpha ),
    .A2(_06325_),
    .Y(_07071_),
    .B1(net4717));
 sg13g2_o21ai_1 _12236_ (.B1(_07071_),
    .Y(_07072_),
    .A1(\soc_inst.spi_inst.cpha ),
    .A2(_06328_));
 sg13g2_nand2_1 _12237_ (.Y(_07073_),
    .A(\soc_inst.spi_inst.state[0] ),
    .B(\soc_inst.spi_inst.cpha ));
 sg13g2_nand4_1 _12238_ (.B(_00123_),
    .C(_07072_),
    .A(net748),
    .Y(_07074_),
    .D(_07073_));
 sg13g2_o21ai_1 _12239_ (.B1(net749),
    .Y(_00349_),
    .A1(_05784_),
    .A2(_07072_));
 sg13g2_xnor2_1 _12240_ (.Y(_07075_),
    .A(net2320),
    .B(net3874));
 sg13g2_nor2_1 _12241_ (.A(net4716),
    .B(_07075_),
    .Y(_00350_));
 sg13g2_a21oi_1 _12242_ (.A1(\soc_inst.spi_inst.bit_counter[0] ),
    .A2(net3874),
    .Y(_07076_),
    .B1(net817));
 sg13g2_and3_1 _12243_ (.X(_07077_),
    .A(\soc_inst.spi_inst.bit_counter[0] ),
    .B(net817),
    .C(net3874));
 sg13g2_nor3_1 _12244_ (.A(net4716),
    .B(net818),
    .C(_07077_),
    .Y(_00351_));
 sg13g2_and4_1 _12245_ (.A(net2320),
    .B(net817),
    .C(net1710),
    .D(_06330_),
    .X(_07078_));
 sg13g2_xnor2_1 _12246_ (.Y(_07079_),
    .A(net1710),
    .B(_07077_));
 sg13g2_nor2_1 _12247_ (.A(net4716),
    .B(net1711),
    .Y(_00352_));
 sg13g2_nor2_1 _12248_ (.A(net1983),
    .B(_07078_),
    .Y(_07080_));
 sg13g2_and2_1 _12249_ (.A(net1983),
    .B(_07078_),
    .X(_07081_));
 sg13g2_nor3_1 _12250_ (.A(net4716),
    .B(net1984),
    .C(_07081_),
    .Y(_00353_));
 sg13g2_nor2_1 _12251_ (.A(net2376),
    .B(_07081_),
    .Y(_07082_));
 sg13g2_and2_1 _12252_ (.A(net2376),
    .B(_07081_),
    .X(_07083_));
 sg13g2_nor3_1 _12253_ (.A(net4716),
    .B(_07082_),
    .C(_07083_),
    .Y(_00354_));
 sg13g2_a21oi_1 _12254_ (.A1(net2539),
    .A2(_07083_),
    .Y(_07084_),
    .B1(net4716));
 sg13g2_o21ai_1 _12255_ (.B1(_07084_),
    .Y(_07085_),
    .A1(net2539),
    .A2(_07083_));
 sg13g2_inv_1 _12256_ (.Y(_00355_),
    .A(_07085_));
 sg13g2_a21oi_1 _12257_ (.A1(_05468_),
    .A2(\soc_inst.spi_inst.state[0] ),
    .Y(_07086_),
    .B1(_06330_));
 sg13g2_a22oi_1 _12258_ (.Y(_07087_),
    .B1(net3783),
    .B2(net2353),
    .A2(net3869),
    .A1(net2));
 sg13g2_inv_1 _12259_ (.Y(_00356_),
    .A(_07087_));
 sg13g2_a22oi_1 _12260_ (.Y(_07088_),
    .B1(net3784),
    .B2(net2337),
    .A2(net3867),
    .A1(\soc_inst.spi_inst.rx_shift_reg[0] ));
 sg13g2_inv_1 _12261_ (.Y(_00357_),
    .A(net2338));
 sg13g2_a22oi_1 _12262_ (.Y(_07089_),
    .B1(net3783),
    .B2(net1730),
    .A2(net3866),
    .A1(\soc_inst.spi_inst.rx_shift_reg[1] ));
 sg13g2_inv_1 _12263_ (.Y(_00358_),
    .A(net1731));
 sg13g2_a22oi_1 _12264_ (.Y(_07090_),
    .B1(net3781),
    .B2(net1924),
    .A2(net3865),
    .A1(net1730));
 sg13g2_inv_1 _12265_ (.Y(_00359_),
    .A(_07090_));
 sg13g2_a22oi_1 _12266_ (.Y(_07091_),
    .B1(net3781),
    .B2(net1552),
    .A2(net3865),
    .A1(\soc_inst.spi_inst.rx_shift_reg[3] ));
 sg13g2_inv_1 _12267_ (.Y(_00360_),
    .A(net1553));
 sg13g2_a22oi_1 _12268_ (.Y(_07092_),
    .B1(net3780),
    .B2(net1663),
    .A2(net3864),
    .A1(net1552));
 sg13g2_inv_1 _12269_ (.Y(_00361_),
    .A(_07092_));
 sg13g2_a22oi_1 _12270_ (.Y(_07093_),
    .B1(net3780),
    .B2(net2160),
    .A2(net3866),
    .A1(net1663));
 sg13g2_inv_1 _12271_ (.Y(_00362_),
    .A(_07093_));
 sg13g2_a22oi_1 _12272_ (.Y(_07094_),
    .B1(net3780),
    .B2(net2140),
    .A2(net3866),
    .A1(\soc_inst.spi_inst.rx_shift_reg[6] ));
 sg13g2_inv_1 _12273_ (.Y(_00363_),
    .A(net2141));
 sg13g2_a22oi_1 _12274_ (.Y(_07095_),
    .B1(net3779),
    .B2(net1635),
    .A2(net3865),
    .A1(\soc_inst.spi_inst.rx_shift_reg[7] ));
 sg13g2_inv_1 _12275_ (.Y(_00364_),
    .A(net1636));
 sg13g2_a22oi_1 _12276_ (.Y(_07096_),
    .B1(net3779),
    .B2(net1789),
    .A2(net3864),
    .A1(net1635));
 sg13g2_inv_1 _12277_ (.Y(_00365_),
    .A(_07096_));
 sg13g2_a22oi_1 _12278_ (.Y(_07097_),
    .B1(net3779),
    .B2(net1948),
    .A2(net3865),
    .A1(net1789));
 sg13g2_inv_1 _12279_ (.Y(_00366_),
    .A(_07097_));
 sg13g2_a22oi_1 _12280_ (.Y(_07098_),
    .B1(net3779),
    .B2(net1920),
    .A2(net3864),
    .A1(\soc_inst.spi_inst.rx_shift_reg[10] ));
 sg13g2_inv_1 _12281_ (.Y(_00367_),
    .A(net1921));
 sg13g2_a22oi_1 _12282_ (.Y(_07099_),
    .B1(net3779),
    .B2(net1762),
    .A2(net3864),
    .A1(\soc_inst.spi_inst.rx_shift_reg[11] ));
 sg13g2_inv_1 _12283_ (.Y(_00368_),
    .A(net1763));
 sg13g2_a22oi_1 _12284_ (.Y(_07100_),
    .B1(net3779),
    .B2(net2087),
    .A2(net3864),
    .A1(net1762));
 sg13g2_inv_1 _12285_ (.Y(_00369_),
    .A(_07100_));
 sg13g2_a22oi_1 _12286_ (.Y(_07101_),
    .B1(net3779),
    .B2(net1977),
    .A2(net3864),
    .A1(\soc_inst.spi_inst.rx_shift_reg[13] ));
 sg13g2_inv_1 _12287_ (.Y(_00370_),
    .A(net1978));
 sg13g2_a22oi_1 _12288_ (.Y(_07102_),
    .B1(net3781),
    .B2(net1733),
    .A2(net3865),
    .A1(\soc_inst.spi_inst.rx_shift_reg[14] ));
 sg13g2_inv_1 _12289_ (.Y(_00371_),
    .A(net1734));
 sg13g2_a22oi_1 _12290_ (.Y(_07103_),
    .B1(net3783),
    .B2(net1664),
    .A2(net3867),
    .A1(\soc_inst.spi_inst.rx_shift_reg[15] ));
 sg13g2_inv_1 _12291_ (.Y(_00372_),
    .A(net1665));
 sg13g2_a22oi_1 _12292_ (.Y(_07104_),
    .B1(net3784),
    .B2(net1667),
    .A2(net3867),
    .A1(net1664));
 sg13g2_inv_1 _12293_ (.Y(_00373_),
    .A(net1668));
 sg13g2_a22oi_1 _12294_ (.Y(_07105_),
    .B1(net3783),
    .B2(net1203),
    .A2(net3867),
    .A1(\soc_inst.spi_inst.rx_shift_reg[17] ));
 sg13g2_inv_1 _12295_ (.Y(_00374_),
    .A(net1204));
 sg13g2_a22oi_1 _12296_ (.Y(_07106_),
    .B1(net3783),
    .B2(net1470),
    .A2(net3867),
    .A1(net1203));
 sg13g2_inv_1 _12297_ (.Y(_00375_),
    .A(_07106_));
 sg13g2_a22oi_1 _12298_ (.Y(_07107_),
    .B1(net3781),
    .B2(net776),
    .A2(net3865),
    .A1(\soc_inst.spi_inst.rx_shift_reg[19] ));
 sg13g2_inv_1 _12299_ (.Y(_00376_),
    .A(net777));
 sg13g2_a22oi_1 _12300_ (.Y(_07108_),
    .B1(net3780),
    .B2(net608),
    .A2(net3864),
    .A1(\soc_inst.spi_inst.rx_shift_reg[20] ));
 sg13g2_inv_1 _12301_ (.Y(_00377_),
    .A(net609));
 sg13g2_a22oi_1 _12302_ (.Y(_07109_),
    .B1(net3779),
    .B2(net788),
    .A2(net3864),
    .A1(net608));
 sg13g2_inv_1 _12303_ (.Y(_00378_),
    .A(_07109_));
 sg13g2_a22oi_1 _12304_ (.Y(_07110_),
    .B1(net3780),
    .B2(net1024),
    .A2(net3865),
    .A1(net788));
 sg13g2_inv_1 _12305_ (.Y(_00379_),
    .A(_07110_));
 sg13g2_a22oi_1 _12306_ (.Y(_07111_),
    .B1(net3782),
    .B2(net649),
    .A2(net3868),
    .A1(\soc_inst.spi_inst.rx_shift_reg[23] ));
 sg13g2_inv_1 _12307_ (.Y(_00380_),
    .A(net650));
 sg13g2_a22oi_1 _12308_ (.Y(_07112_),
    .B1(net3782),
    .B2(net709),
    .A2(net3868),
    .A1(net649));
 sg13g2_inv_1 _12309_ (.Y(_00381_),
    .A(_07112_));
 sg13g2_a22oi_1 _12310_ (.Y(_07113_),
    .B1(net3782),
    .B2(net1078),
    .A2(net3867),
    .A1(net709));
 sg13g2_inv_1 _12311_ (.Y(_00382_),
    .A(_07113_));
 sg13g2_a22oi_1 _12312_ (.Y(_07114_),
    .B1(net3782),
    .B2(net974),
    .A2(net3867),
    .A1(\soc_inst.spi_inst.rx_shift_reg[26] ));
 sg13g2_inv_1 _12313_ (.Y(_00383_),
    .A(net975));
 sg13g2_a22oi_1 _12314_ (.Y(_07115_),
    .B1(net3783),
    .B2(net681),
    .A2(net3868),
    .A1(\soc_inst.spi_inst.rx_shift_reg[27] ));
 sg13g2_inv_1 _12315_ (.Y(_00384_),
    .A(net682));
 sg13g2_a22oi_1 _12316_ (.Y(_07116_),
    .B1(net3783),
    .B2(net890),
    .A2(net3868),
    .A1(net681));
 sg13g2_inv_1 _12317_ (.Y(_00385_),
    .A(_07116_));
 sg13g2_a22oi_1 _12318_ (.Y(_07117_),
    .B1(net3783),
    .B2(net1249),
    .A2(net3867),
    .A1(net890));
 sg13g2_inv_1 _12319_ (.Y(_00386_),
    .A(_07117_));
 sg13g2_a22oi_1 _12320_ (.Y(_07118_),
    .B1(net3784),
    .B2(net432),
    .A2(net3868),
    .A1(\soc_inst.spi_inst.rx_shift_reg[30] ));
 sg13g2_inv_1 _12321_ (.Y(_00387_),
    .A(net433));
 sg13g2_nor2_1 _12322_ (.A(_06305_),
    .B(_06525_),
    .Y(_07119_));
 sg13g2_mux2_1 _12323_ (.A0(net2682),
    .A1(net5026),
    .S(net3985),
    .X(_00388_));
 sg13g2_nand2_2 _12324_ (.Y(_07120_),
    .A(_06288_),
    .B(_06411_));
 sg13g2_nor2_1 _12325_ (.A(_06300_),
    .B(_07120_),
    .Y(_07121_));
 sg13g2_mux2_1 _12326_ (.A0(net2687),
    .A1(net5049),
    .S(_07121_),
    .X(_00389_));
 sg13g2_nor2_1 _12327_ (.A(net2521),
    .B(net3983),
    .Y(_07122_));
 sg13g2_a21oi_1 _12328_ (.A1(net5048),
    .A2(net3983),
    .Y(_00390_),
    .B1(_07122_));
 sg13g2_nor2_1 _12329_ (.A(net2088),
    .B(net3983),
    .Y(_07123_));
 sg13g2_a21oi_1 _12330_ (.A1(net5045),
    .A2(net3983),
    .Y(_00391_),
    .B1(_07123_));
 sg13g2_nor2_1 _12331_ (.A(net1683),
    .B(net3983),
    .Y(_07124_));
 sg13g2_a21oi_1 _12332_ (.A1(net5042),
    .A2(net3983),
    .Y(_00392_),
    .B1(_07124_));
 sg13g2_nor2_1 _12333_ (.A(net1433),
    .B(net3983),
    .Y(_07125_));
 sg13g2_a21oi_1 _12334_ (.A1(net5039),
    .A2(net3984),
    .Y(_00393_),
    .B1(_07125_));
 sg13g2_nor2_1 _12335_ (.A(net1869),
    .B(net3983),
    .Y(_07126_));
 sg13g2_a21oi_1 _12336_ (.A1(net5036),
    .A2(net3984),
    .Y(_00394_),
    .B1(_07126_));
 sg13g2_mux2_1 _12337_ (.A0(net2477),
    .A1(net5034),
    .S(net3984),
    .X(_00395_));
 sg13g2_mux2_1 _12338_ (.A0(net2303),
    .A1(net5031),
    .S(net3984),
    .X(_00396_));
 sg13g2_mux2_1 _12339_ (.A0(net2237),
    .A1(net5029),
    .S(net3985),
    .X(_00397_));
 sg13g2_a22oi_1 _12340_ (.Y(_07127_),
    .B1(net622),
    .B2(_07017_),
    .A2(\soc_inst.spi_inst.state[0] ),
    .A1(net520));
 sg13g2_inv_1 _12341_ (.Y(_00398_),
    .A(net623));
 sg13g2_mux2_1 _12342_ (.A0(net2630),
    .A1(net5025),
    .S(net3985),
    .X(_00399_));
 sg13g2_nor2b_1 _12343_ (.A(\soc_inst.gpio_inst.gpio_sync2[0] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[0] ),
    .Y(_07128_));
 sg13g2_a21oi_1 _12344_ (.A1(net87),
    .A2(_07128_),
    .Y(_07129_),
    .B1(net467));
 sg13g2_nand2_2 _12345_ (.Y(_07130_),
    .A(net4785),
    .B(_05897_));
 sg13g2_nor2_2 _12346_ (.A(_07069_),
    .B(_07130_),
    .Y(_07131_));
 sg13g2_a21oi_1 _12347_ (.A1(net5049),
    .A2(_07131_),
    .Y(_00400_),
    .B1(net468));
 sg13g2_mux2_1 _12348_ (.A0(net5128),
    .A1(net5042),
    .S(_06414_),
    .X(_00401_));
 sg13g2_mux2_1 _12349_ (.A0(net2149),
    .A1(net5038),
    .S(_06414_),
    .X(_00402_));
 sg13g2_mux2_1 _12350_ (.A0(net933),
    .A1(net5036),
    .S(_06414_),
    .X(_00403_));
 sg13g2_nor4_1 _12351_ (.A(net158),
    .B(net13),
    .C(net5128),
    .D(_06975_),
    .Y(_07132_));
 sg13g2_a21o_1 _12352_ (.A2(net159),
    .A1(_06972_),
    .B1(net89),
    .X(_00404_));
 sg13g2_nor2_1 _12353_ (.A(_06296_),
    .B(_06413_),
    .Y(_07133_));
 sg13g2_nor2_1 _12354_ (.A(net2065),
    .B(net3982),
    .Y(_07134_));
 sg13g2_a21oi_1 _12355_ (.A1(net5050),
    .A2(net3982),
    .Y(_00405_),
    .B1(_07134_));
 sg13g2_nor2_1 _12356_ (.A(net1725),
    .B(net3981),
    .Y(_07135_));
 sg13g2_a21oi_1 _12357_ (.A1(net5046),
    .A2(net3981),
    .Y(_00406_),
    .B1(_07135_));
 sg13g2_nor2_1 _12358_ (.A(net1618),
    .B(net3981),
    .Y(_07136_));
 sg13g2_a21oi_1 _12359_ (.A1(net5042),
    .A2(net3981),
    .Y(_00407_),
    .B1(_07136_));
 sg13g2_nor2_1 _12360_ (.A(net1952),
    .B(net3981),
    .Y(_07137_));
 sg13g2_a21oi_1 _12361_ (.A1(net5039),
    .A2(net3981),
    .Y(_00408_),
    .B1(_07137_));
 sg13g2_nor2_1 _12362_ (.A(net1729),
    .B(net3981),
    .Y(_07138_));
 sg13g2_a21oi_1 _12363_ (.A1(net5036),
    .A2(net3981),
    .Y(_00409_),
    .B1(_07138_));
 sg13g2_mux2_1 _12364_ (.A0(net2357),
    .A1(net5034),
    .S(net3982),
    .X(_00410_));
 sg13g2_mux2_1 _12365_ (.A0(net2137),
    .A1(net5032),
    .S(net3982),
    .X(_00411_));
 sg13g2_nor2_1 _12366_ (.A(net1890),
    .B(net3982),
    .Y(_07139_));
 sg13g2_a21oi_1 _12367_ (.A1(net5029),
    .A2(net3982),
    .Y(_00412_),
    .B1(_07139_));
 sg13g2_nand2_1 _12368_ (.Y(_07140_),
    .A(_06442_),
    .B(_06928_));
 sg13g2_o21ai_1 _12369_ (.B1(_06965_),
    .Y(_07141_),
    .A1(_06441_),
    .A2(_06969_));
 sg13g2_a21o_1 _12370_ (.A2(_07140_),
    .A1(net4274),
    .B1(_07141_),
    .X(_07142_));
 sg13g2_nand2b_2 _12371_ (.Y(_07143_),
    .B(_06963_),
    .A_N(_07142_));
 sg13g2_nand3b_1 _12372_ (.B(_06963_),
    .C(_06964_),
    .Y(_07144_),
    .A_N(_07142_));
 sg13g2_nand2_1 _12373_ (.Y(_07145_),
    .A(net592),
    .B(_07143_));
 sg13g2_o21ai_1 _12374_ (.B1(_07145_),
    .Y(_00413_),
    .A1(net592),
    .A2(_07144_));
 sg13g2_nand2_1 _12375_ (.Y(_07146_),
    .A(net952),
    .B(_07143_));
 sg13g2_nand2_1 _12376_ (.Y(_07147_),
    .A(net592),
    .B(net952));
 sg13g2_xnor2_1 _12377_ (.Y(_07148_),
    .A(net592),
    .B(net952));
 sg13g2_o21ai_1 _12378_ (.B1(_07146_),
    .Y(_00414_),
    .A1(_07144_),
    .A2(_07148_));
 sg13g2_nand3_1 _12379_ (.B(net952),
    .C(net1482),
    .A(net592),
    .Y(_07149_));
 sg13g2_a21oi_1 _12380_ (.A1(_06964_),
    .A2(_07149_),
    .Y(_07150_),
    .B1(_07143_));
 sg13g2_nor2_1 _12381_ (.A(_07143_),
    .B(_07147_),
    .Y(_07151_));
 sg13g2_nor2_1 _12382_ (.A(net1482),
    .B(_07151_),
    .Y(_07152_));
 sg13g2_nor2_1 _12383_ (.A(_07150_),
    .B(_07152_),
    .Y(_00415_));
 sg13g2_or3_1 _12384_ (.A(net1122),
    .B(_07144_),
    .C(_07149_),
    .X(_07153_));
 sg13g2_o21ai_1 _12385_ (.B1(_07153_),
    .Y(_00416_),
    .A1(_05568_),
    .A2(_07150_));
 sg13g2_nor2_2 _12386_ (.A(net5117),
    .B(_06418_),
    .Y(_07154_));
 sg13g2_nand2_1 _12387_ (.Y(_07155_),
    .A(_06418_),
    .B(_06438_));
 sg13g2_nand2_1 _12388_ (.Y(_07156_),
    .A(net2662),
    .B(_06439_));
 sg13g2_a21oi_1 _12389_ (.A1(_06417_),
    .A2(_07156_),
    .Y(_07157_),
    .B1(_07155_));
 sg13g2_nor2_1 _12390_ (.A(\soc_inst.i2c_inst.state[1] ),
    .B(_06440_),
    .Y(_07158_));
 sg13g2_nor2_1 _12391_ (.A(_07154_),
    .B(_07158_),
    .Y(_07159_));
 sg13g2_nand2_1 _12392_ (.Y(_07160_),
    .A(\soc_inst.i2c_ena ),
    .B(_07159_));
 sg13g2_a22oi_1 _12393_ (.Y(_07161_),
    .B1(_07158_),
    .B2(_06973_),
    .A2(_07157_),
    .A1(net4274));
 sg13g2_o21ai_1 _12394_ (.B1(_07161_),
    .Y(_07162_),
    .A1(_07157_),
    .A2(_07160_));
 sg13g2_a21oi_1 _12395_ (.A1(net4274),
    .A2(_07154_),
    .Y(_07163_),
    .B1(_07162_));
 sg13g2_nand2_1 _12396_ (.Y(_07164_),
    .A(net5120),
    .B(_07158_));
 sg13g2_a21oi_1 _12397_ (.A1(net5128),
    .A2(\soc_inst.i2c_inst.ack_enable ),
    .Y(_07165_),
    .B1(_07164_));
 sg13g2_o21ai_1 _12398_ (.B1(_06964_),
    .Y(_07166_),
    .A1(\soc_inst.i2c_inst.ctrl_reg[2] ),
    .A2(net1183));
 sg13g2_nor2_1 _12399_ (.A(_07159_),
    .B(_07165_),
    .Y(_07167_));
 sg13g2_nand3_1 _12400_ (.B(net1184),
    .C(_07167_),
    .A(_07163_),
    .Y(_07168_));
 sg13g2_o21ai_1 _12401_ (.B1(net1185),
    .Y(_00417_),
    .A1(_05405_),
    .A2(_07163_));
 sg13g2_nand3_1 _12402_ (.B(\soc_inst.i2c_inst.state[1] ),
    .C(_06439_),
    .A(net5120),
    .Y(_07169_));
 sg13g2_nor2_1 _12403_ (.A(net5120),
    .B(_06417_),
    .Y(_07170_));
 sg13g2_o21ai_1 _12404_ (.B1(_07169_),
    .Y(_07171_),
    .A1(net5117),
    .A2(_06442_));
 sg13g2_or2_1 _12405_ (.X(_07172_),
    .B(_07171_),
    .A(_07170_));
 sg13g2_nor2_1 _12406_ (.A(net5120),
    .B(net5118),
    .Y(_07173_));
 sg13g2_nor3_1 _12407_ (.A(_06020_),
    .B(_06439_),
    .C(_07173_),
    .Y(_07174_));
 sg13g2_a22oi_1 _12408_ (.Y(_07175_),
    .B1(_07174_),
    .B2(_06975_),
    .A2(_07172_),
    .A1(net4275));
 sg13g2_and2_1 _12409_ (.A(net4275),
    .B(_07174_),
    .X(_07176_));
 sg13g2_nor4_1 _12410_ (.A(_06023_),
    .B(_06443_),
    .C(_07170_),
    .D(_07176_),
    .Y(_07177_));
 sg13g2_mux2_1 _12411_ (.A0(net1054),
    .A1(_07177_),
    .S(_07175_),
    .X(_00418_));
 sg13g2_nand2b_1 _12412_ (.Y(_00419_),
    .B(_07068_),
    .A_N(net91));
 sg13g2_nor2_1 _12413_ (.A(net1306),
    .B(net3999),
    .Y(_07178_));
 sg13g2_a21oi_1 _12414_ (.A1(net5047),
    .A2(net3999),
    .Y(_00420_),
    .B1(_07178_));
 sg13g2_nor2_1 _12415_ (.A(net1501),
    .B(net3999),
    .Y(_07179_));
 sg13g2_a21oi_1 _12416_ (.A1(net5044),
    .A2(net3999),
    .Y(_00421_),
    .B1(_07179_));
 sg13g2_nor2_1 _12417_ (.A(net1598),
    .B(net3999),
    .Y(_07180_));
 sg13g2_a21oi_1 _12418_ (.A1(net5041),
    .A2(net3999),
    .Y(_00422_),
    .B1(_07180_));
 sg13g2_nor2_1 _12419_ (.A(net1376),
    .B(net3999),
    .Y(_07181_));
 sg13g2_a21oi_1 _12420_ (.A1(net5038),
    .A2(net3999),
    .Y(_00423_),
    .B1(_07181_));
 sg13g2_nor2_1 _12421_ (.A(net1632),
    .B(net3998),
    .Y(_07182_));
 sg13g2_a21oi_1 _12422_ (.A1(net5035),
    .A2(net3998),
    .Y(_00424_),
    .B1(_07182_));
 sg13g2_nor2_1 _12423_ (.A(net1343),
    .B(net3998),
    .Y(_07183_));
 sg13g2_a21oi_1 _12424_ (.A1(net5033),
    .A2(net3998),
    .Y(_00425_),
    .B1(_07183_));
 sg13g2_nor2_1 _12425_ (.A(net1829),
    .B(net3998),
    .Y(_07184_));
 sg13g2_a21oi_1 _12426_ (.A1(net5032),
    .A2(net3998),
    .Y(_00426_),
    .B1(_07184_));
 sg13g2_nor2_1 _12427_ (.A(net1544),
    .B(net3998),
    .Y(_07185_));
 sg13g2_a21oi_1 _12428_ (.A1(net5028),
    .A2(net3998),
    .Y(_00427_),
    .B1(_07185_));
 sg13g2_nor2_1 _12429_ (.A(net2129),
    .B(net3996),
    .Y(_07186_));
 sg13g2_a21oi_1 _12430_ (.A1(net5026),
    .A2(net3996),
    .Y(_00428_),
    .B1(_07186_));
 sg13g2_nor2_1 _12431_ (.A(net2119),
    .B(net3996),
    .Y(_07187_));
 sg13g2_a21oi_1 _12432_ (.A1(net5024),
    .A2(net3996),
    .Y(_00429_),
    .B1(_07187_));
 sg13g2_nor2_1 _12433_ (.A(net1671),
    .B(net3996),
    .Y(_07188_));
 sg13g2_a21oi_1 _12434_ (.A1(net5023),
    .A2(net3996),
    .Y(_00430_),
    .B1(_07188_));
 sg13g2_nor2_1 _12435_ (.A(net1563),
    .B(net3996),
    .Y(_07189_));
 sg13g2_a21oi_1 _12436_ (.A1(net5022),
    .A2(net3996),
    .Y(_00431_),
    .B1(_07189_));
 sg13g2_nor2_1 _12437_ (.A(net1485),
    .B(net3997),
    .Y(_07190_));
 sg13g2_a21oi_1 _12438_ (.A1(net5021),
    .A2(net3997),
    .Y(_00432_),
    .B1(_07190_));
 sg13g2_nor2_1 _12439_ (.A(net1765),
    .B(net3997),
    .Y(_07191_));
 sg13g2_a21oi_1 _12440_ (.A1(net5020),
    .A2(net3997),
    .Y(_00433_),
    .B1(_07191_));
 sg13g2_nor2_1 _12441_ (.A(net1831),
    .B(net3997),
    .Y(_07192_));
 sg13g2_a21oi_1 _12442_ (.A1(net5019),
    .A2(net4000),
    .Y(_00434_),
    .B1(_07192_));
 sg13g2_nor2_1 _12443_ (.A(net1222),
    .B(net3997),
    .Y(_07193_));
 sg13g2_a21oi_1 _12444_ (.A1(net5018),
    .A2(net4000),
    .Y(_00435_),
    .B1(_07193_));
 sg13g2_nor2_1 _12445_ (.A(net1942),
    .B(net4003),
    .Y(_07194_));
 sg13g2_a21oi_1 _12446_ (.A1(net5047),
    .A2(net4003),
    .Y(_00436_),
    .B1(_07194_));
 sg13g2_nor2_1 _12447_ (.A(net1866),
    .B(net4003),
    .Y(_07195_));
 sg13g2_a21oi_1 _12448_ (.A1(net5044),
    .A2(net4003),
    .Y(_00437_),
    .B1(_07195_));
 sg13g2_nor2_1 _12449_ (.A(net1754),
    .B(net4003),
    .Y(_07196_));
 sg13g2_a21oi_1 _12450_ (.A1(net5041),
    .A2(net4003),
    .Y(_00438_),
    .B1(_07196_));
 sg13g2_nor2_1 _12451_ (.A(net1745),
    .B(net4005),
    .Y(_07197_));
 sg13g2_a21oi_1 _12452_ (.A1(net5038),
    .A2(net4005),
    .Y(_00439_),
    .B1(_07197_));
 sg13g2_nor2_1 _12453_ (.A(net1397),
    .B(net4004),
    .Y(_07198_));
 sg13g2_a21oi_1 _12454_ (.A1(net5035),
    .A2(net4004),
    .Y(_00440_),
    .B1(_07198_));
 sg13g2_nor2_1 _12455_ (.A(net1279),
    .B(net4004),
    .Y(_07199_));
 sg13g2_a21oi_1 _12456_ (.A1(net5033),
    .A2(net4004),
    .Y(_00441_),
    .B1(_07199_));
 sg13g2_nor2_1 _12457_ (.A(net1695),
    .B(net4004),
    .Y(_07200_));
 sg13g2_a21oi_1 _12458_ (.A1(net5032),
    .A2(net4004),
    .Y(_00442_),
    .B1(_07200_));
 sg13g2_nor2_1 _12459_ (.A(net1639),
    .B(net4004),
    .Y(_07201_));
 sg13g2_a21oi_1 _12460_ (.A1(net5028),
    .A2(net4004),
    .Y(_00443_),
    .B1(_07201_));
 sg13g2_nor2_1 _12461_ (.A(net1603),
    .B(net4001),
    .Y(_07202_));
 sg13g2_a21oi_1 _12462_ (.A1(net5026),
    .A2(net4001),
    .Y(_00444_),
    .B1(_07202_));
 sg13g2_nor2_1 _12463_ (.A(net1743),
    .B(net4001),
    .Y(_07203_));
 sg13g2_a21oi_1 _12464_ (.A1(net5024),
    .A2(net4001),
    .Y(_00445_),
    .B1(_07203_));
 sg13g2_nor2_1 _12465_ (.A(net2024),
    .B(net4001),
    .Y(_07204_));
 sg13g2_a21oi_1 _12466_ (.A1(net5023),
    .A2(net4001),
    .Y(_00446_),
    .B1(_07204_));
 sg13g2_nor2_1 _12467_ (.A(net1850),
    .B(net4001),
    .Y(_07205_));
 sg13g2_a21oi_1 _12468_ (.A1(net5022),
    .A2(net4001),
    .Y(_00447_),
    .B1(_07205_));
 sg13g2_nor2_1 _12469_ (.A(net1330),
    .B(net4002),
    .Y(_07206_));
 sg13g2_a21oi_1 _12470_ (.A1(net5021),
    .A2(net4002),
    .Y(_00448_),
    .B1(_07206_));
 sg13g2_nor2_1 _12471_ (.A(net1644),
    .B(net4002),
    .Y(_07207_));
 sg13g2_a21oi_1 _12472_ (.A1(net5020),
    .A2(net4002),
    .Y(_00449_),
    .B1(_07207_));
 sg13g2_nor2_1 _12473_ (.A(net1554),
    .B(net4003),
    .Y(_07208_));
 sg13g2_a21oi_1 _12474_ (.A1(net5019),
    .A2(net4003),
    .Y(_00450_),
    .B1(_07208_));
 sg13g2_nor2_1 _12475_ (.A(net1970),
    .B(net4002),
    .Y(_07209_));
 sg13g2_a21oi_1 _12476_ (.A1(net5018),
    .A2(net4002),
    .Y(_00451_),
    .B1(_07209_));
 sg13g2_nor2_2 _12477_ (.A(_06289_),
    .B(net4269),
    .Y(_07210_));
 sg13g2_nor2b_2 _12478_ (.A(_06526_),
    .B_N(net4178),
    .Y(_07211_));
 sg13g2_mux2_1 _12479_ (.A0(net1990),
    .A1(net5047),
    .S(_07211_),
    .X(_00452_));
 sg13g2_mux2_1 _12480_ (.A0(net1757),
    .A1(net5044),
    .S(net3980),
    .X(_00453_));
 sg13g2_mux2_1 _12481_ (.A0(net1631),
    .A1(net5041),
    .S(net3980),
    .X(_00454_));
 sg13g2_mux2_1 _12482_ (.A0(net2365),
    .A1(net5038),
    .S(net3980),
    .X(_00455_));
 sg13g2_mux2_1 _12483_ (.A0(net2262),
    .A1(net5035),
    .S(net3979),
    .X(_00456_));
 sg13g2_mux2_1 _12484_ (.A0(net2161),
    .A1(net5033),
    .S(net3979),
    .X(_00457_));
 sg13g2_mux2_1 _12485_ (.A0(net2322),
    .A1(net5032),
    .S(net3980),
    .X(_00458_));
 sg13g2_mux2_1 _12486_ (.A0(net882),
    .A1(net5028),
    .S(net3980),
    .X(_00459_));
 sg13g2_mux2_1 _12487_ (.A0(net2363),
    .A1(net5026),
    .S(net3979),
    .X(_00460_));
 sg13g2_mux2_1 _12488_ (.A0(net2449),
    .A1(net5024),
    .S(net3979),
    .X(_00461_));
 sg13g2_mux2_1 _12489_ (.A0(net2080),
    .A1(net5023),
    .S(net3979),
    .X(_00462_));
 sg13g2_mux2_1 _12490_ (.A0(net1904),
    .A1(net5022),
    .S(net3979),
    .X(_00463_));
 sg13g2_mux2_1 _12491_ (.A0(net1839),
    .A1(net5021),
    .S(net3979),
    .X(_00464_));
 sg13g2_mux2_1 _12492_ (.A0(net2293),
    .A1(net5020),
    .S(net3979),
    .X(_00465_));
 sg13g2_mux2_1 _12493_ (.A0(net2094),
    .A1(net5019),
    .S(net3980),
    .X(_00466_));
 sg13g2_mux2_1 _12494_ (.A0(net2375),
    .A1(net5018),
    .S(net3980),
    .X(_00467_));
 sg13g2_mux2_1 _12495_ (.A0(net2482),
    .A1(net5045),
    .S(_00133_),
    .X(_00468_));
 sg13g2_mux2_1 _12496_ (.A0(net5126),
    .A1(net5043),
    .S(_00133_),
    .X(_00469_));
 sg13g2_nand3_1 _12497_ (.B(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .C(\soc_inst.cpu_core.mem_reg_we ),
    .A(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .Y(_07212_));
 sg13g2_nand2_2 _12498_ (.Y(_07213_),
    .A(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[3] ));
 sg13g2_nor2_2 _12499_ (.A(_07212_),
    .B(_07213_),
    .Y(_07214_));
 sg13g2_nor4_1 _12500_ (.A(_05403_),
    .B(\soc_inst.cpu_core.mem_instr[5] ),
    .C(\soc_inst.cpu_core.mem_instr[6] ),
    .D(_06678_),
    .Y(_07215_));
 sg13g2_or4_1 _12501_ (.A(_05403_),
    .B(\soc_inst.cpu_core.mem_instr[5] ),
    .C(\soc_inst.cpu_core.mem_instr[6] ),
    .D(_06678_),
    .X(_07216_));
 sg13g2_nor2_2 _12502_ (.A(net4755),
    .B(net4754),
    .Y(_07217_));
 sg13g2_nand2_2 _12503_ (.Y(_07218_),
    .A(net4871),
    .B(net4866));
 sg13g2_nor3_2 _12504_ (.A(_06738_),
    .B(_07216_),
    .C(_07217_),
    .Y(_07219_));
 sg13g2_a21oi_1 _12505_ (.A1(_05483_),
    .A2(net4242),
    .Y(_07220_),
    .B1(net4626));
 sg13g2_a22oi_1 _12506_ (.Y(_07221_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[0] ),
    .A2(net4191),
    .A1(\soc_inst.cpu_core.csr_file.mepc[0] ));
 sg13g2_a22oi_1 _12507_ (.Y(_07222_),
    .B1(net4186),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[0] ),
    .A2(net4255),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[0] ));
 sg13g2_a221oi_1 _12508_ (.B2(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .C1(net4245),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .Y(_07223_),
    .A2(net4237));
 sg13g2_inv_4 _12509_ (.A(_07223_),
    .Y(_07224_));
 sg13g2_a221oi_1 _12510_ (.B2(\soc_inst.cpu_core.csr_file.mtval[0] ),
    .C1(_07224_),
    .B1(net4088),
    .A1(\soc_inst.cpu_core.csr_file.mcause[0] ),
    .Y(_07225_),
    .A2(net4095));
 sg13g2_nand3_1 _12511_ (.B(_07222_),
    .C(_07225_),
    .A(_07221_),
    .Y(_07226_));
 sg13g2_a22oi_1 _12512_ (.Y(_07227_),
    .B1(_07220_),
    .B2(_07226_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[0] ));
 sg13g2_nor2_1 _12513_ (.A(net1146),
    .B(net4637),
    .Y(_07228_));
 sg13g2_a21oi_1 _12514_ (.A1(net4637),
    .A2(net3944),
    .Y(_00470_),
    .B1(_07228_));
 sg13g2_a21oi_1 _12515_ (.A1(_05482_),
    .A2(net4242),
    .Y(_07229_),
    .B1(net4626));
 sg13g2_a22oi_1 _12516_ (.Y(_07230_),
    .B1(net4191),
    .B2(\soc_inst.cpu_core.csr_file.mepc[1] ),
    .A2(net4255),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[1] ));
 sg13g2_a22oi_1 _12517_ (.Y(_07231_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[1] ),
    .A2(net4186),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[1] ));
 sg13g2_a221oi_1 _12518_ (.B2(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .C1(net4245),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .Y(_07232_),
    .A2(net4237));
 sg13g2_inv_4 _12519_ (.A(_07232_),
    .Y(_07233_));
 sg13g2_a221oi_1 _12520_ (.B2(\soc_inst.cpu_core.csr_file.mtval[1] ),
    .C1(_07233_),
    .B1(net4088),
    .A1(\soc_inst.cpu_core.csr_file.mcause[1] ),
    .Y(_07234_),
    .A2(net4095));
 sg13g2_nand3_1 _12521_ (.B(_07231_),
    .C(_07234_),
    .A(_07230_),
    .Y(_07235_));
 sg13g2_a22oi_1 _12522_ (.Y(_07236_),
    .B1(_07229_),
    .B2(_07235_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[1] ));
 sg13g2_nor2_1 _12523_ (.A(net2145),
    .B(net4636),
    .Y(_07237_));
 sg13g2_a21oi_1 _12524_ (.A1(net4636),
    .A2(net3943),
    .Y(_00471_),
    .B1(_07237_));
 sg13g2_a21oi_1 _12525_ (.A1(_05484_),
    .A2(net4242),
    .Y(_07238_),
    .B1(net4626));
 sg13g2_a22oi_1 _12526_ (.Y(_07239_),
    .B1(net4183),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[2] ),
    .A2(net4255),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[2] ));
 sg13g2_nor2_2 _12527_ (.A(net4240),
    .B(_06712_),
    .Y(_07240_));
 sg13g2_nand2_1 _12528_ (.Y(_07241_),
    .A(\soc_inst.cpu_core.csr_file.mtvec[2] ),
    .B(net4186));
 sg13g2_a22oi_1 _12529_ (.Y(_07242_),
    .B1(net4234),
    .B2(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .A2(net4237),
    .A1(\soc_inst.cpu_core.csr_file.mtime[34] ));
 sg13g2_o21ai_1 _12530_ (.B1(_07242_),
    .Y(_07243_),
    .A1(_05614_),
    .A2(_06692_));
 sg13g2_a221oi_1 _12531_ (.B2(\soc_inst.cpu_core.csr_file.mtval[2] ),
    .C1(_07243_),
    .B1(net4089),
    .A1(\soc_inst.cpu_core.csr_file.mcause[2] ),
    .Y(_07244_),
    .A2(net4096));
 sg13g2_nand4_1 _12532_ (.B(_07240_),
    .C(_07241_),
    .A(_07239_),
    .Y(_07245_),
    .D(_07244_));
 sg13g2_a22oi_1 _12533_ (.Y(_07246_),
    .B1(_07238_),
    .B2(_07245_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[2] ));
 sg13g2_nor2_1 _12534_ (.A(net981),
    .B(net4640),
    .Y(_07247_));
 sg13g2_a21oi_1 _12535_ (.A1(net4637),
    .A2(net3940),
    .Y(_00472_),
    .B1(_07247_));
 sg13g2_a21oi_1 _12536_ (.A1(_05485_),
    .A2(net4242),
    .Y(_07248_),
    .B1(net4627));
 sg13g2_a22oi_1 _12537_ (.Y(_07249_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[3] ),
    .A2(net4256),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[3] ));
 sg13g2_a22oi_1 _12538_ (.Y(_07250_),
    .B1(net4186),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[3] ),
    .A2(net4191),
    .A1(\soc_inst.cpu_core.csr_file.mepc[3] ));
 sg13g2_a221oi_1 _12539_ (.B2(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .C1(net4245),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .Y(_07251_),
    .A2(net4237));
 sg13g2_inv_4 _12540_ (.A(_07251_),
    .Y(_07252_));
 sg13g2_a221oi_1 _12541_ (.B2(\soc_inst.cpu_core.csr_file.mtval[3] ),
    .C1(_07252_),
    .B1(net4088),
    .A1(\soc_inst.cpu_core.csr_file.mcause[3] ),
    .Y(_07253_),
    .A2(net4095));
 sg13g2_nand3_1 _12542_ (.B(_07250_),
    .C(_07253_),
    .A(_07249_),
    .Y(_07254_));
 sg13g2_a22oi_1 _12543_ (.Y(_07255_),
    .B1(_07248_),
    .B2(_07254_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[3] ));
 sg13g2_nor2_1 _12544_ (.A(net1547),
    .B(net4636),
    .Y(_07256_));
 sg13g2_a21oi_1 _12545_ (.A1(net4636),
    .A2(net3938),
    .Y(_00473_),
    .B1(_07256_));
 sg13g2_a21oi_1 _12546_ (.A1(_05487_),
    .A2(net4243),
    .Y(_07257_),
    .B1(net4628));
 sg13g2_a22oi_1 _12547_ (.Y(_07258_),
    .B1(net4192),
    .B2(\soc_inst.cpu_core.csr_file.mepc[4] ),
    .A2(net4255),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[4] ));
 sg13g2_a22oi_1 _12548_ (.Y(_07259_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[4] ),
    .A2(net4186),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[4] ));
 sg13g2_a22oi_1 _12549_ (.Y(_07260_),
    .B1(net4233),
    .B2(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .A2(net4237),
    .A1(\soc_inst.cpu_core.csr_file.mtime[36] ));
 sg13g2_nand2_1 _12550_ (.Y(_07261_),
    .A(_07240_),
    .B(_07260_));
 sg13g2_a221oi_1 _12551_ (.B2(\soc_inst.cpu_core.csr_file.mtval[4] ),
    .C1(_07261_),
    .B1(net4090),
    .A1(\soc_inst.cpu_core.csr_file.mcause[4] ),
    .Y(_07262_),
    .A2(net4096));
 sg13g2_nand3_1 _12552_ (.B(_07259_),
    .C(_07262_),
    .A(_07258_),
    .Y(_07263_));
 sg13g2_a22oi_1 _12553_ (.Y(_07264_),
    .B1(_07257_),
    .B2(_07263_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[4] ));
 sg13g2_nor2_1 _12554_ (.A(net1013),
    .B(net4639),
    .Y(_07265_));
 sg13g2_a21oi_1 _12555_ (.A1(net4639),
    .A2(net3835),
    .Y(_00474_),
    .B1(_07265_));
 sg13g2_a21oi_1 _12556_ (.A1(_05486_),
    .A2(net4243),
    .Y(_07266_),
    .B1(net4628));
 sg13g2_a22oi_1 _12557_ (.Y(_07267_),
    .B1(net4187),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[5] ),
    .A2(net4193),
    .A1(\soc_inst.cpu_core.csr_file.mepc[5] ));
 sg13g2_a22oi_1 _12558_ (.Y(_07268_),
    .B1(net4183),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[5] ),
    .A2(net4256),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[5] ));
 sg13g2_a221oi_1 _12559_ (.B2(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .C1(net4245),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .Y(_07269_),
    .A2(net4238));
 sg13g2_inv_1 _12560_ (.Y(_07270_),
    .A(_07269_));
 sg13g2_a221oi_1 _12561_ (.B2(\soc_inst.cpu_core.csr_file.mtval[5] ),
    .C1(_07270_),
    .B1(net4093),
    .A1(\soc_inst.cpu_core.csr_file.mcause[5] ),
    .Y(_07271_),
    .A2(net4098));
 sg13g2_nand3_1 _12562_ (.B(_07268_),
    .C(_07271_),
    .A(_07267_),
    .Y(_07272_));
 sg13g2_a22oi_1 _12563_ (.Y(_07273_),
    .B1(_07266_),
    .B2(_07272_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[5] ));
 sg13g2_nor2_1 _12564_ (.A(net1438),
    .B(net4639),
    .Y(_07274_));
 sg13g2_a21oi_1 _12565_ (.A1(net4639),
    .A2(net3935),
    .Y(_00475_),
    .B1(_07274_));
 sg13g2_a21oi_1 _12566_ (.A1(_05488_),
    .A2(net4243),
    .Y(_07275_),
    .B1(net4628));
 sg13g2_a22oi_1 _12567_ (.Y(_07276_),
    .B1(net4183),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[6] ),
    .A2(net4193),
    .A1(\soc_inst.cpu_core.csr_file.mepc[6] ));
 sg13g2_a22oi_1 _12568_ (.Y(_07277_),
    .B1(net4187),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[6] ),
    .A2(net4257),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[6] ));
 sg13g2_a221oi_1 _12569_ (.B2(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .C1(net4245),
    .B1(net4234),
    .A1(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .Y(_07278_),
    .A2(net4238));
 sg13g2_inv_1 _12570_ (.Y(_07279_),
    .A(_07278_));
 sg13g2_a221oi_1 _12571_ (.B2(\soc_inst.cpu_core.csr_file.mtval[6] ),
    .C1(_07279_),
    .B1(net4093),
    .A1(\soc_inst.cpu_core.csr_file.mcause[6] ),
    .Y(_07280_),
    .A2(net4098));
 sg13g2_nand3_1 _12572_ (.B(_07277_),
    .C(_07280_),
    .A(_07276_),
    .Y(_07281_));
 sg13g2_a22oi_1 _12573_ (.Y(_07282_),
    .B1(_07275_),
    .B2(_07281_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[6] ));
 sg13g2_nor2_1 _12574_ (.A(net703),
    .B(net4639),
    .Y(_07283_));
 sg13g2_a21oi_1 _12575_ (.A1(net4640),
    .A2(net3932),
    .Y(_00476_),
    .B1(_07283_));
 sg13g2_a21oi_1 _12576_ (.A1(_05489_),
    .A2(net4243),
    .Y(_07284_),
    .B1(net4628));
 sg13g2_a22oi_1 _12577_ (.Y(_07285_),
    .B1(_06713_),
    .B2(\soc_inst.cpu_core.csr_file.mip_tip ),
    .A2(net4256),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[7] ));
 sg13g2_a22oi_1 _12578_ (.Y(_07286_),
    .B1(net4182),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[7] ),
    .A2(net4186),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[7] ));
 sg13g2_a221oi_1 _12579_ (.B2(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .C1(net4245),
    .B1(net4234),
    .A1(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .Y(_07287_),
    .A2(net4237));
 sg13g2_a22oi_1 _12580_ (.Y(_07288_),
    .B1(_06695_),
    .B2(\soc_inst.cpu_core.csr_file.mie[7] ),
    .A2(net4193),
    .A1(\soc_inst.cpu_core.csr_file.mepc[7] ));
 sg13g2_and2_1 _12581_ (.A(_07287_),
    .B(_07288_),
    .X(_07289_));
 sg13g2_a22oi_1 _12582_ (.Y(_07290_),
    .B1(net4093),
    .B2(\soc_inst.cpu_core.csr_file.mtval[7] ),
    .A2(net4098),
    .A1(\soc_inst.cpu_core.csr_file.mcause[7] ));
 sg13g2_nand4_1 _12583_ (.B(_07286_),
    .C(_07289_),
    .A(_07285_),
    .Y(_07291_),
    .D(_07290_));
 sg13g2_a22oi_1 _12584_ (.Y(_07292_),
    .B1(_07284_),
    .B2(_07291_),
    .A2(_07219_),
    .A1(\soc_inst.core_mem_rdata[7] ));
 sg13g2_nor2_1 _12585_ (.A(net921),
    .B(net4636),
    .Y(_07293_));
 sg13g2_a21oi_1 _12586_ (.A1(net4636),
    .A2(net3931),
    .Y(_00477_),
    .B1(_07293_));
 sg13g2_nand2_2 _12587_ (.Y(_07294_),
    .A(\soc_inst.core_mem_rdata[7] ),
    .B(_06676_));
 sg13g2_nor2_2 _12588_ (.A(net4231),
    .B(_07217_),
    .Y(_07295_));
 sg13g2_nand2_1 _12589_ (.Y(_07296_),
    .A(\soc_inst.core_mem_rdata[8] ),
    .B(net4177));
 sg13g2_nand2_1 _12590_ (.Y(_07297_),
    .A(net4228),
    .B(_07296_));
 sg13g2_a21oi_1 _12591_ (.A1(_05418_),
    .A2(net4246),
    .Y(_07298_),
    .B1(net4629));
 sg13g2_a22oi_1 _12592_ (.Y(_07299_),
    .B1(net4194),
    .B2(\soc_inst.cpu_core.csr_file.mepc[8] ),
    .A2(net4257),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[8] ));
 sg13g2_a22oi_1 _12593_ (.Y(_07300_),
    .B1(net4182),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[8] ),
    .A2(net4187),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[8] ));
 sg13g2_a221oi_1 _12594_ (.B2(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .C1(net4246),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .Y(_07301_),
    .A2(net4237));
 sg13g2_inv_1 _12595_ (.Y(_07302_),
    .A(_07301_));
 sg13g2_a221oi_1 _12596_ (.B2(\soc_inst.cpu_core.csr_file.mtval[8] ),
    .C1(_07302_),
    .B1(net4093),
    .A1(\soc_inst.cpu_core.csr_file.mcause[8] ),
    .Y(_07303_),
    .A2(net4098));
 sg13g2_nand3_1 _12597_ (.B(_07300_),
    .C(_07303_),
    .A(_07299_),
    .Y(_07304_));
 sg13g2_a22oi_1 _12598_ (.Y(_07305_),
    .B1(_07298_),
    .B2(_07304_),
    .A2(_07297_),
    .A1(net4629));
 sg13g2_nor2_1 _12599_ (.A(net1288),
    .B(net4632),
    .Y(_07306_));
 sg13g2_a21oi_1 _12600_ (.A1(net4632),
    .A2(net3928),
    .Y(_00478_),
    .B1(_07306_));
 sg13g2_nand2_1 _12601_ (.Y(_07307_),
    .A(\soc_inst.core_mem_rdata[9] ),
    .B(net4177));
 sg13g2_nand2_1 _12602_ (.Y(_07308_),
    .A(net4228),
    .B(_07307_));
 sg13g2_a21oi_1 _12603_ (.A1(_05419_),
    .A2(net4242),
    .Y(_07309_),
    .B1(net4626));
 sg13g2_a22oi_1 _12604_ (.Y(_07310_),
    .B1(net4193),
    .B2(\soc_inst.cpu_core.csr_file.mepc[9] ),
    .A2(net4256),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[9] ));
 sg13g2_a22oi_1 _12605_ (.Y(_07311_),
    .B1(net4182),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[9] ),
    .A2(net4187),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[9] ));
 sg13g2_a221oi_1 _12606_ (.B2(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .C1(net4244),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .Y(_07312_),
    .A2(net4237));
 sg13g2_inv_1 _12607_ (.Y(_07313_),
    .A(_07312_));
 sg13g2_a221oi_1 _12608_ (.B2(\soc_inst.cpu_core.csr_file.mtval[9] ),
    .C1(_07313_),
    .B1(net4093),
    .A1(\soc_inst.cpu_core.csr_file.mcause[9] ),
    .Y(_07314_),
    .A2(net4098));
 sg13g2_nand3_1 _12609_ (.B(_07311_),
    .C(_07314_),
    .A(_07310_),
    .Y(_07315_));
 sg13g2_a22oi_1 _12610_ (.Y(_07316_),
    .B1(_07309_),
    .B2(_07315_),
    .A2(_07308_),
    .A1(net4628));
 sg13g2_nor2_1 _12611_ (.A(net901),
    .B(net4638),
    .Y(_07317_));
 sg13g2_a21oi_1 _12612_ (.A1(net4638),
    .A2(net3926),
    .Y(_00479_),
    .B1(_07317_));
 sg13g2_nand2_1 _12613_ (.Y(_07318_),
    .A(\soc_inst.core_mem_rdata[10] ),
    .B(net4177));
 sg13g2_nand2_1 _12614_ (.Y(_07319_),
    .A(net4228),
    .B(_07318_));
 sg13g2_a21oi_1 _12615_ (.A1(_05421_),
    .A2(net4242),
    .Y(_07320_),
    .B1(net4626));
 sg13g2_a22oi_1 _12616_ (.Y(_07321_),
    .B1(net4183),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[10] ),
    .A2(net4257),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[10] ));
 sg13g2_a22oi_1 _12617_ (.Y(_07322_),
    .B1(net4187),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[10] ),
    .A2(net4193),
    .A1(\soc_inst.cpu_core.csr_file.mepc[10] ));
 sg13g2_a221oi_1 _12618_ (.B2(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .C1(net4244),
    .B1(net4233),
    .A1(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .Y(_07323_),
    .A2(net4238));
 sg13g2_inv_1 _12619_ (.Y(_07324_),
    .A(_07323_));
 sg13g2_a221oi_1 _12620_ (.B2(\soc_inst.cpu_core.csr_file.mtval[10] ),
    .C1(_07324_),
    .B1(net4093),
    .A1(\soc_inst.cpu_core.csr_file.mcause[10] ),
    .Y(_07325_),
    .A2(net4098));
 sg13g2_nand3_1 _12621_ (.B(_07322_),
    .C(_07325_),
    .A(_07321_),
    .Y(_07326_));
 sg13g2_a22oi_1 _12622_ (.Y(_07327_),
    .B1(_07320_),
    .B2(_07326_),
    .A2(_07319_),
    .A1(net4626));
 sg13g2_nor2_1 _12623_ (.A(net1707),
    .B(net4637),
    .Y(_07328_));
 sg13g2_a21oi_1 _12624_ (.A1(net4637),
    .A2(net3925),
    .Y(_00480_),
    .B1(_07328_));
 sg13g2_nand2_1 _12625_ (.Y(_07329_),
    .A(\soc_inst.core_mem_rdata[11] ),
    .B(net4177));
 sg13g2_nand2_1 _12626_ (.Y(_07330_),
    .A(net4228),
    .B(_07329_));
 sg13g2_a22oi_1 _12627_ (.Y(_07331_),
    .B1(net4182),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[11] ),
    .A2(net4186),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[11] ));
 sg13g2_a22oi_1 _12628_ (.Y(_07332_),
    .B1(_06713_),
    .B2(\soc_inst.cpu_core.csr_file.mip_eip ),
    .A2(net4257),
    .A1(_05398_));
 sg13g2_and2_1 _12629_ (.A(_07331_),
    .B(_07332_),
    .X(_07333_));
 sg13g2_a22oi_1 _12630_ (.Y(_07334_),
    .B1(net4093),
    .B2(\soc_inst.cpu_core.csr_file.mtval[11] ),
    .A2(net4098),
    .A1(\soc_inst.cpu_core.csr_file.mcause[11] ));
 sg13g2_a22oi_1 _12631_ (.Y(_07335_),
    .B1(_06695_),
    .B2(\soc_inst.cpu_core.csr_file.mie[11] ),
    .A2(net4193),
    .A1(\soc_inst.cpu_core.csr_file.mepc[11] ));
 sg13g2_a221oi_1 _12632_ (.B2(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .C1(net4245),
    .B1(net4235),
    .A1(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .Y(_07336_),
    .A2(net4238));
 sg13g2_nand4_1 _12633_ (.B(_07334_),
    .C(_07335_),
    .A(_07333_),
    .Y(_07337_),
    .D(_07336_));
 sg13g2_a21oi_1 _12634_ (.A1(_05420_),
    .A2(net4243),
    .Y(_07338_),
    .B1(net4626));
 sg13g2_a22oi_1 _12635_ (.Y(_07339_),
    .B1(_07337_),
    .B2(_07338_),
    .A2(_07330_),
    .A1(net4628));
 sg13g2_nor2_1 _12636_ (.A(net1806),
    .B(net4636),
    .Y(_07340_));
 sg13g2_a21oi_1 _12637_ (.A1(net4636),
    .A2(net3922),
    .Y(_00481_),
    .B1(_07340_));
 sg13g2_nand2_1 _12638_ (.Y(_07341_),
    .A(\soc_inst.core_mem_rdata[12] ),
    .B(net4177));
 sg13g2_nand2_1 _12639_ (.Y(_07342_),
    .A(net4228),
    .B(_07341_));
 sg13g2_a21oi_1 _12640_ (.A1(_05423_),
    .A2(net4243),
    .Y(_07343_),
    .B1(net4628));
 sg13g2_a221oi_1 _12641_ (.B2(\soc_inst.cpu_core.csr_file.mtval[12] ),
    .C1(_06721_),
    .B1(_06820_),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[12] ),
    .Y(_07344_),
    .A2(net4184));
 sg13g2_nand2_1 _12642_ (.Y(_07345_),
    .A(\soc_inst.cpu_core.csr_file.mscratch[12] ),
    .B(_06723_));
 sg13g2_o21ai_1 _12643_ (.B1(_07345_),
    .Y(_07346_),
    .A1(_00294_),
    .A2(_06672_));
 sg13g2_a221oi_1 _12644_ (.B2(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .C1(_07346_),
    .B1(net4236),
    .A1(\soc_inst.cpu_core.csr_file.mepc[12] ),
    .Y(_07347_),
    .A2(net4190));
 sg13g2_a22oi_1 _12645_ (.Y(_07348_),
    .B1(_06797_),
    .B2(\soc_inst.cpu_core.csr_file.mcause[12] ),
    .A2(net4239),
    .A1(\soc_inst.cpu_core.csr_file.mtime[44] ));
 sg13g2_nand3_1 _12646_ (.B(_07347_),
    .C(_07348_),
    .A(_07344_),
    .Y(_07349_));
 sg13g2_a22oi_1 _12647_ (.Y(_07350_),
    .B1(_07343_),
    .B2(_07349_),
    .A2(_07342_),
    .A1(net4628));
 sg13g2_nor2_1 _12648_ (.A(net1232),
    .B(net4640),
    .Y(_07351_));
 sg13g2_a21oi_1 _12649_ (.A1(net4640),
    .A2(net3833),
    .Y(_00482_),
    .B1(_07351_));
 sg13g2_nand2_1 _12650_ (.Y(_07352_),
    .A(\soc_inst.core_mem_rdata[13] ),
    .B(net4177));
 sg13g2_nand2_2 _12651_ (.Y(_07353_),
    .A(net4228),
    .B(_07352_));
 sg13g2_a21oi_1 _12652_ (.A1(_05422_),
    .A2(net4241),
    .Y(_07354_),
    .B1(net4630));
 sg13g2_a22oi_1 _12653_ (.Y(_07355_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[13] ),
    .A2(net4256),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[13] ));
 sg13g2_a22oi_1 _12654_ (.Y(_07356_),
    .B1(net4186),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[13] ),
    .A2(net4192),
    .A1(\soc_inst.cpu_core.csr_file.mepc[13] ));
 sg13g2_a221oi_1 _12655_ (.B2(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .C1(net4244),
    .B1(net4235),
    .A1(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .Y(_07357_),
    .A2(net4238));
 sg13g2_inv_2 _12656_ (.Y(_07358_),
    .A(_07357_));
 sg13g2_a221oi_1 _12657_ (.B2(\soc_inst.cpu_core.csr_file.mtval[13] ),
    .C1(_07358_),
    .B1(net4090),
    .A1(\soc_inst.cpu_core.csr_file.mcause[13] ),
    .Y(_07359_),
    .A2(net4096));
 sg13g2_nand3_1 _12658_ (.B(_07356_),
    .C(_07359_),
    .A(_07355_),
    .Y(_07360_));
 sg13g2_a22oi_1 _12659_ (.Y(_07361_),
    .B1(_07354_),
    .B2(_07360_),
    .A2(_07353_),
    .A1(net4624));
 sg13g2_nor2_1 _12660_ (.A(net889),
    .B(net4632),
    .Y(_07362_));
 sg13g2_a21oi_1 _12661_ (.A1(net4632),
    .A2(net3919),
    .Y(_00483_),
    .B1(_07362_));
 sg13g2_nand2_1 _12662_ (.Y(_07363_),
    .A(\soc_inst.core_mem_rdata[14] ),
    .B(_07295_));
 sg13g2_nand2_1 _12663_ (.Y(_07364_),
    .A(_07294_),
    .B(_07363_));
 sg13g2_a21oi_1 _12664_ (.A1(_05425_),
    .A2(net4246),
    .Y(_07365_),
    .B1(net4629));
 sg13g2_a22oi_1 _12665_ (.Y(_07366_),
    .B1(net4183),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[14] ),
    .A2(net4193),
    .A1(\soc_inst.cpu_core.csr_file.mepc[14] ));
 sg13g2_a22oi_1 _12666_ (.Y(_07367_),
    .B1(net4187),
    .B2(\soc_inst.cpu_core.csr_file.mtvec[14] ),
    .A2(net4257),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[14] ));
 sg13g2_a221oi_1 _12667_ (.B2(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .C1(net4244),
    .B1(net4235),
    .A1(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .Y(_07368_),
    .A2(net4238));
 sg13g2_inv_1 _12668_ (.Y(_07369_),
    .A(_07368_));
 sg13g2_a221oi_1 _12669_ (.B2(\soc_inst.cpu_core.csr_file.mtval[14] ),
    .C1(_07369_),
    .B1(net4093),
    .A1(\soc_inst.cpu_core.csr_file.mcause[14] ),
    .Y(_07370_),
    .A2(net4098));
 sg13g2_nand3_1 _12670_ (.B(_07367_),
    .C(_07370_),
    .A(_07366_),
    .Y(_07371_));
 sg13g2_a22oi_1 _12671_ (.Y(_07372_),
    .B1(_07365_),
    .B2(_07371_),
    .A2(_07364_),
    .A1(net4629));
 sg13g2_nor2_1 _12672_ (.A(net1225),
    .B(net4639),
    .Y(_07373_));
 sg13g2_a21oi_1 _12673_ (.A1(net4639),
    .A2(net3917),
    .Y(_00484_),
    .B1(_07373_));
 sg13g2_nand2_1 _12674_ (.Y(_07374_),
    .A(\soc_inst.core_mem_rdata[15] ),
    .B(_07295_));
 sg13g2_nand2_2 _12675_ (.Y(_07375_),
    .A(net4228),
    .B(_07374_));
 sg13g2_a21oi_1 _12676_ (.A1(_05424_),
    .A2(net4242),
    .Y(_07376_),
    .B1(net4627));
 sg13g2_a22oi_1 _12677_ (.Y(_07377_),
    .B1(net4189),
    .B2(\soc_inst.cpu_core.csr_file.mepc[15] ),
    .A2(net4251),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[15] ));
 sg13g2_a22oi_1 _12678_ (.Y(_07378_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[15] ),
    .A2(net4184),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[15] ));
 sg13g2_a221oi_1 _12679_ (.B2(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .C1(net4244),
    .B1(net4235),
    .A1(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .Y(_07379_),
    .A2(net4238));
 sg13g2_inv_2 _12680_ (.Y(_07380_),
    .A(_07379_));
 sg13g2_a221oi_1 _12681_ (.B2(\soc_inst.cpu_core.csr_file.mtval[15] ),
    .C1(_07380_),
    .B1(net4092),
    .A1(\soc_inst.cpu_core.csr_file.mcause[15] ),
    .Y(_07381_),
    .A2(net4097));
 sg13g2_nand3_1 _12682_ (.B(_07378_),
    .C(_07381_),
    .A(_07377_),
    .Y(_07382_));
 sg13g2_a22oi_1 _12683_ (.Y(_07383_),
    .B1(_07376_),
    .B2(_07382_),
    .A2(_07375_),
    .A1(net4630));
 sg13g2_nor2_1 _12684_ (.A(net1398),
    .B(net4634),
    .Y(_07384_));
 sg13g2_a21oi_1 _12685_ (.A1(net4634),
    .A2(net3916),
    .Y(_00485_),
    .B1(_07384_));
 sg13g2_nor2_1 _12686_ (.A(net4869),
    .B(_06750_),
    .Y(_07385_));
 sg13g2_nand2_1 _12687_ (.Y(_07386_),
    .A(\soc_inst.core_mem_rdata[15] ),
    .B(net4227));
 sg13g2_nand2_1 _12688_ (.Y(_07387_),
    .A(net4228),
    .B(_07386_));
 sg13g2_nor2_1 _12689_ (.A(net4868),
    .B(_06748_),
    .Y(_07388_));
 sg13g2_nand2b_1 _12690_ (.Y(_07389_),
    .B(net4753),
    .A_N(_06748_));
 sg13g2_a21o_2 _12691_ (.A2(net4619),
    .A1(\soc_inst.core_mem_rdata[16] ),
    .B1(net4085),
    .X(_07390_));
 sg13g2_a21oi_1 _12692_ (.A1(_05426_),
    .A2(net4240),
    .Y(_07391_),
    .B1(net4624));
 sg13g2_a22oi_1 _12693_ (.Y(_07392_),
    .B1(net4190),
    .B2(\soc_inst.cpu_core.csr_file.mepc[16] ),
    .A2(net4252),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[16] ));
 sg13g2_a21oi_1 _12694_ (.A1(\soc_inst.cpu_core.csr_file.mscratch[16] ),
    .A2(net4181),
    .Y(_07393_),
    .B1(net4240));
 sg13g2_a22oi_1 _12695_ (.Y(_07394_),
    .B1(net4232),
    .B2(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .A2(net4185),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[16] ));
 sg13g2_a22oi_1 _12696_ (.Y(_07395_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[16] ),
    .A2(net4097),
    .A1(\soc_inst.cpu_core.csr_file.mcause[16] ));
 sg13g2_nand4_1 _12697_ (.B(_07393_),
    .C(_07394_),
    .A(_07392_),
    .Y(_07396_),
    .D(_07395_));
 sg13g2_a22oi_1 _12698_ (.Y(_07397_),
    .B1(_07391_),
    .B2(_07396_),
    .A2(_07390_),
    .A1(net4624));
 sg13g2_nor2_1 _12699_ (.A(net876),
    .B(net4632),
    .Y(_07398_));
 sg13g2_a21oi_1 _12700_ (.A1(net4632),
    .A2(net3911),
    .Y(_00486_),
    .B1(_07398_));
 sg13g2_a21oi_2 _12701_ (.B1(net4085),
    .Y(_07399_),
    .A2(net4619),
    .A1(\soc_inst.core_mem_rdata[17] ));
 sg13g2_nand2_1 _12702_ (.Y(_07400_),
    .A(\soc_inst.cpu_core.csr_file.mstatus[17] ),
    .B(net4252));
 sg13g2_a22oi_1 _12703_ (.Y(_07401_),
    .B1(net4181),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[17] ),
    .A2(net4185),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[17] ));
 sg13g2_a221oi_1 _12704_ (.B2(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .C1(net4240),
    .B1(net4232),
    .A1(\soc_inst.cpu_core.csr_file.mepc[17] ),
    .Y(_07402_),
    .A2(net4190));
 sg13g2_a22oi_1 _12705_ (.Y(_07403_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[17] ),
    .A2(net4097),
    .A1(\soc_inst.cpu_core.csr_file.mcause[17] ));
 sg13g2_nand4_1 _12706_ (.B(_07401_),
    .C(_07402_),
    .A(_07400_),
    .Y(_07404_),
    .D(_07403_));
 sg13g2_o21ai_1 _12707_ (.B1(_07404_),
    .Y(_07405_),
    .A1(\soc_inst.core_mem_addr[17] ),
    .A2(net4247));
 sg13g2_mux2_1 _12708_ (.A0(_07399_),
    .A1(_07405_),
    .S(_07216_),
    .X(_07406_));
 sg13g2_nor2_1 _12709_ (.A(net1853),
    .B(net4633),
    .Y(_07407_));
 sg13g2_a21oi_1 _12710_ (.A1(net4633),
    .A2(net3831),
    .Y(_00487_),
    .B1(_07407_));
 sg13g2_a21o_2 _12711_ (.A2(net4619),
    .A1(\soc_inst.core_mem_rdata[18] ),
    .B1(net4085),
    .X(_07408_));
 sg13g2_a21oi_1 _12712_ (.A1(_05428_),
    .A2(net4240),
    .Y(_07409_),
    .B1(net4624));
 sg13g2_a22oi_1 _12713_ (.Y(_07410_),
    .B1(net4189),
    .B2(\soc_inst.cpu_core.csr_file.mepc[18] ),
    .A2(net4249),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[18] ));
 sg13g2_a21oi_1 _12714_ (.A1(\soc_inst.cpu_core.csr_file.mtval[18] ),
    .A2(_06820_),
    .Y(_07411_),
    .B1(_06721_));
 sg13g2_a22oi_1 _12715_ (.Y(_07412_),
    .B1(_06723_),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[18] ),
    .A2(net4184),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[18] ));
 sg13g2_a22oi_1 _12716_ (.Y(_07413_),
    .B1(_06797_),
    .B2(\soc_inst.cpu_core.csr_file.mcause[18] ),
    .A2(net4235),
    .A1(\soc_inst.cpu_core.csr_file.mtime[18] ));
 sg13g2_nand4_1 _12717_ (.B(_07411_),
    .C(_07412_),
    .A(_07410_),
    .Y(_07414_),
    .D(_07413_));
 sg13g2_a22oi_1 _12718_ (.Y(_07415_),
    .B1(_07409_),
    .B2(_07414_),
    .A2(_07408_),
    .A1(net4624));
 sg13g2_nor2_1 _12719_ (.A(net1506),
    .B(net4631),
    .Y(_07416_));
 sg13g2_a21oi_1 _12720_ (.A1(net4631),
    .A2(net3909),
    .Y(_00488_),
    .B1(_07416_));
 sg13g2_a21o_2 _12721_ (.A2(net4619),
    .A1(\soc_inst.core_mem_rdata[19] ),
    .B1(net4085),
    .X(_07417_));
 sg13g2_a21oi_1 _12722_ (.A1(_05427_),
    .A2(net4240),
    .Y(_07418_),
    .B1(net4624));
 sg13g2_a22oi_1 _12723_ (.Y(_07419_),
    .B1(net4189),
    .B2(\soc_inst.cpu_core.csr_file.mepc[19] ),
    .A2(net4249),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[19] ));
 sg13g2_a22oi_1 _12724_ (.Y(_07420_),
    .B1(_06820_),
    .B2(\soc_inst.cpu_core.csr_file.mtval[19] ),
    .A2(_06797_),
    .A1(\soc_inst.cpu_core.csr_file.mcause[19] ));
 sg13g2_a22oi_1 _12725_ (.Y(_07421_),
    .B1(_06723_),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[19] ),
    .A2(net4184),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[19] ));
 sg13g2_a21oi_1 _12726_ (.A1(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .A2(net4236),
    .Y(_07422_),
    .B1(_06721_));
 sg13g2_nand4_1 _12727_ (.B(_07420_),
    .C(_07421_),
    .A(_07419_),
    .Y(_07423_),
    .D(_07422_));
 sg13g2_a22oi_1 _12728_ (.Y(_07424_),
    .B1(_07418_),
    .B2(_07423_),
    .A2(_07417_),
    .A1(net4624));
 sg13g2_nor2_1 _12729_ (.A(net1971),
    .B(net4633),
    .Y(_07425_));
 sg13g2_a21oi_1 _12730_ (.A1(net4633),
    .A2(net3906),
    .Y(_00489_),
    .B1(_07425_));
 sg13g2_a21o_2 _12731_ (.A2(net4619),
    .A1(\soc_inst.core_mem_rdata[20] ),
    .B1(net4085),
    .X(_07426_));
 sg13g2_a21oi_1 _12732_ (.A1(_05430_),
    .A2(net4241),
    .Y(_07427_),
    .B1(net4625));
 sg13g2_a22oi_1 _12733_ (.Y(_07428_),
    .B1(net4097),
    .B2(\soc_inst.cpu_core.csr_file.mcause[20] ),
    .A2(net4190),
    .A1(\soc_inst.cpu_core.csr_file.mepc[20] ));
 sg13g2_a21oi_1 _12734_ (.A1(\soc_inst.cpu_core.csr_file.mstatus[20] ),
    .A2(net4250),
    .Y(_07429_),
    .B1(net4240));
 sg13g2_a22oi_1 _12735_ (.Y(_07430_),
    .B1(net4232),
    .B2(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .A2(net4181),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[20] ));
 sg13g2_a22oi_1 _12736_ (.Y(_07431_),
    .B1(net4091),
    .B2(\soc_inst.cpu_core.csr_file.mtval[20] ),
    .A2(net4184),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[20] ));
 sg13g2_nand4_1 _12737_ (.B(_07429_),
    .C(_07430_),
    .A(_07428_),
    .Y(_07432_),
    .D(_07431_));
 sg13g2_a22oi_1 _12738_ (.Y(_07433_),
    .B1(_07427_),
    .B2(_07432_),
    .A2(_07426_),
    .A1(net4624));
 sg13g2_nor2_1 _12739_ (.A(net1599),
    .B(net4631),
    .Y(_07434_));
 sg13g2_a21oi_1 _12740_ (.A1(net4631),
    .A2(net3904),
    .Y(_00490_),
    .B1(_07434_));
 sg13g2_a21o_2 _12741_ (.A2(net4619),
    .A1(\soc_inst.core_mem_rdata[21] ),
    .B1(net4085),
    .X(_07435_));
 sg13g2_a21oi_1 _12742_ (.A1(_05429_),
    .A2(net4241),
    .Y(_07436_),
    .B1(net4625));
 sg13g2_a22oi_1 _12743_ (.Y(_07437_),
    .B1(net4232),
    .B2(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .A2(net4250),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[21] ));
 sg13g2_a21oi_1 _12744_ (.A1(\soc_inst.cpu_core.csr_file.mtvec[21] ),
    .A2(net4184),
    .Y(_07438_),
    .B1(net4241));
 sg13g2_a22oi_1 _12745_ (.Y(_07439_),
    .B1(net4091),
    .B2(\soc_inst.cpu_core.csr_file.mtval[21] ),
    .A2(net4100),
    .A1(\soc_inst.cpu_core.csr_file.mcause[21] ));
 sg13g2_a22oi_1 _12746_ (.Y(_07440_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[21] ),
    .A2(net4189),
    .A1(\soc_inst.cpu_core.csr_file.mepc[21] ));
 sg13g2_nand4_1 _12747_ (.B(_07438_),
    .C(_07439_),
    .A(_07437_),
    .Y(_07441_),
    .D(_07440_));
 sg13g2_a22oi_1 _12748_ (.Y(_07442_),
    .B1(_07436_),
    .B2(_07441_),
    .A2(_07435_),
    .A1(net4625));
 sg13g2_nor2_1 _12749_ (.A(net1099),
    .B(net4633),
    .Y(_07443_));
 sg13g2_a21oi_1 _12750_ (.A1(net4633),
    .A2(net3902),
    .Y(_00491_),
    .B1(_07443_));
 sg13g2_a21o_2 _12751_ (.A2(net4619),
    .A1(\soc_inst.core_mem_rdata[22] ),
    .B1(net4086),
    .X(_07444_));
 sg13g2_a21oi_1 _12752_ (.A1(_05432_),
    .A2(net4241),
    .Y(_07445_),
    .B1(net4625));
 sg13g2_a21oi_1 _12753_ (.A1(\soc_inst.cpu_core.csr_file.mtval[22] ),
    .A2(_06820_),
    .Y(_07446_),
    .B1(_06721_));
 sg13g2_a22oi_1 _12754_ (.Y(_07447_),
    .B1(_06723_),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[22] ),
    .A2(net4184),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[22] ));
 sg13g2_a22oi_1 _12755_ (.Y(_07448_),
    .B1(net4189),
    .B2(\soc_inst.cpu_core.csr_file.mepc[22] ),
    .A2(net4250),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[22] ));
 sg13g2_a22oi_1 _12756_ (.Y(_07449_),
    .B1(_06797_),
    .B2(\soc_inst.cpu_core.csr_file.mcause[22] ),
    .A2(net4235),
    .A1(\soc_inst.cpu_core.csr_file.mtime[22] ));
 sg13g2_nand4_1 _12757_ (.B(_07447_),
    .C(_07448_),
    .A(_07446_),
    .Y(_07450_),
    .D(_07449_));
 sg13g2_a22oi_1 _12758_ (.Y(_07451_),
    .B1(_07445_),
    .B2(_07450_),
    .A2(_07444_),
    .A1(net4625));
 sg13g2_nor2_1 _12759_ (.A(net1650),
    .B(net4633),
    .Y(_07452_));
 sg13g2_a21oi_1 _12760_ (.A1(net4633),
    .A2(net3900),
    .Y(_00492_),
    .B1(_07452_));
 sg13g2_a21o_2 _12761_ (.A2(net4620),
    .A1(\soc_inst.core_mem_rdata[23] ),
    .B1(net4086),
    .X(_07453_));
 sg13g2_a21oi_1 _12762_ (.A1(_05431_),
    .A2(net4241),
    .Y(_07454_),
    .B1(net4625));
 sg13g2_a22oi_1 _12763_ (.Y(_07455_),
    .B1(net4180),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[23] ),
    .A2(net4184),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[23] ));
 sg13g2_a21oi_2 _12764_ (.B1(net4244),
    .Y(_07456_),
    .A2(net4232),
    .A1(\soc_inst.cpu_core.csr_file.mtime[23] ));
 sg13g2_a22oi_1 _12765_ (.Y(_07457_),
    .B1(net4091),
    .B2(\soc_inst.cpu_core.csr_file.mtval[23] ),
    .A2(net4249),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[23] ));
 sg13g2_a22oi_1 _12766_ (.Y(_07458_),
    .B1(net4100),
    .B2(\soc_inst.cpu_core.csr_file.mcause[23] ),
    .A2(net4189),
    .A1(\soc_inst.cpu_core.csr_file.mepc[23] ));
 sg13g2_nand4_1 _12767_ (.B(_07456_),
    .C(_07457_),
    .A(_07455_),
    .Y(_07459_),
    .D(_07458_));
 sg13g2_a22oi_1 _12768_ (.Y(_07460_),
    .B1(_07454_),
    .B2(_07459_),
    .A2(_07453_),
    .A1(net4625));
 sg13g2_nor2_1 _12769_ (.A(net1685),
    .B(net4631),
    .Y(_07461_));
 sg13g2_a21oi_1 _12770_ (.A1(net4631),
    .A2(net3897),
    .Y(_00493_),
    .B1(_07461_));
 sg13g2_a21oi_2 _12771_ (.B1(net4087),
    .Y(_07462_),
    .A2(net4621),
    .A1(\soc_inst.core_mem_rdata[24] ));
 sg13g2_a22oi_1 _12772_ (.Y(_07463_),
    .B1(net4094),
    .B2(\soc_inst.cpu_core.csr_file.mtval[24] ),
    .A2(net4097),
    .A1(\soc_inst.cpu_core.csr_file.mcause[24] ));
 sg13g2_a21oi_1 _12773_ (.A1(\soc_inst.cpu_core.csr_file.mscratch[24] ),
    .A2(net4182),
    .Y(_07464_),
    .B1(net4244));
 sg13g2_a22oi_1 _12774_ (.Y(_07465_),
    .B1(_06716_),
    .B2(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .A2(net4254),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[24] ));
 sg13g2_nand3_1 _12775_ (.B(_07464_),
    .C(_07465_),
    .A(_07463_),
    .Y(_07466_));
 sg13g2_o21ai_1 _12776_ (.B1(_07466_),
    .Y(_07467_),
    .A1(\soc_inst.core_mem_addr[24] ),
    .A2(net4247));
 sg13g2_mux2_1 _12777_ (.A0(_07462_),
    .A1(_07467_),
    .S(_07216_),
    .X(_07468_));
 sg13g2_nor2_1 _12778_ (.A(net1820),
    .B(net4638),
    .Y(_07469_));
 sg13g2_a21oi_1 _12779_ (.A1(net4638),
    .A2(net3830),
    .Y(_00494_),
    .B1(_07469_));
 sg13g2_a21oi_2 _12780_ (.B1(net4087),
    .Y(_07470_),
    .A2(net4621),
    .A1(\soc_inst.core_mem_rdata[25] ));
 sg13g2_a22oi_1 _12781_ (.Y(_07471_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[25] ),
    .A2(net4097),
    .A1(\soc_inst.cpu_core.csr_file.mcause[25] ));
 sg13g2_nand2_1 _12782_ (.Y(_07472_),
    .A(\soc_inst.cpu_core.csr_file.mstatus[25] ),
    .B(net4253));
 sg13g2_a22oi_1 _12783_ (.Y(_07473_),
    .B1(net4232),
    .B2(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .A2(net4182),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[25] ));
 sg13g2_nand4_1 _12784_ (.B(_07471_),
    .C(_07472_),
    .A(net4247),
    .Y(_07474_),
    .D(_07473_));
 sg13g2_o21ai_1 _12785_ (.B1(_07474_),
    .Y(_07475_),
    .A1(\soc_inst.core_mem_addr[25] ),
    .A2(net4247));
 sg13g2_mux2_1 _12786_ (.A0(_07470_),
    .A1(_07475_),
    .S(_07216_),
    .X(_07476_));
 sg13g2_nor2_1 _12787_ (.A(net881),
    .B(net4638),
    .Y(_07477_));
 sg13g2_a21oi_1 _12788_ (.A1(net4638),
    .A2(net3827),
    .Y(_00495_),
    .B1(_07477_));
 sg13g2_a21oi_2 _12789_ (.B1(net4087),
    .Y(_07478_),
    .A2(net4621),
    .A1(\soc_inst.core_mem_rdata[26] ));
 sg13g2_a21oi_1 _12790_ (.A1(\soc_inst.cpu_core.csr_file.mcause[26] ),
    .A2(net4099),
    .Y(_07479_),
    .B1(net4244));
 sg13g2_a22oi_1 _12791_ (.Y(_07480_),
    .B1(_06716_),
    .B2(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .A2(net4258),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[26] ));
 sg13g2_a22oi_1 _12792_ (.Y(_07481_),
    .B1(net4094),
    .B2(\soc_inst.cpu_core.csr_file.mtval[26] ),
    .A2(net4181),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[26] ));
 sg13g2_nand3_1 _12793_ (.B(_07480_),
    .C(_07481_),
    .A(_07479_),
    .Y(_07482_));
 sg13g2_o21ai_1 _12794_ (.B1(_07482_),
    .Y(_07483_),
    .A1(\soc_inst.core_mem_addr[26] ),
    .A2(net4247));
 sg13g2_mux2_1 _12795_ (.A0(_07478_),
    .A1(_07483_),
    .S(_07216_),
    .X(_07484_));
 sg13g2_nor2_1 _12796_ (.A(net1280),
    .B(net4637),
    .Y(_07485_));
 sg13g2_a21oi_1 _12797_ (.A1(net4637),
    .A2(net3824),
    .Y(_00496_),
    .B1(_07485_));
 sg13g2_a21o_2 _12798_ (.A2(net4620),
    .A1(\soc_inst.core_mem_rdata[27] ),
    .B1(net4086),
    .X(_07486_));
 sg13g2_a21oi_2 _12799_ (.B1(net4626),
    .Y(_07487_),
    .A2(net4243),
    .A1(_05433_));
 sg13g2_a22oi_1 _12800_ (.Y(_07488_),
    .B1(_06820_),
    .B2(\soc_inst.cpu_core.csr_file.mtval[27] ),
    .A2(_06797_),
    .A1(\soc_inst.cpu_core.csr_file.mcause[27] ));
 sg13g2_a21oi_1 _12801_ (.A1(\soc_inst.cpu_core.csr_file.mscratch[27] ),
    .A2(_06723_),
    .Y(_07489_),
    .B1(_06721_));
 sg13g2_a22oi_1 _12802_ (.Y(_07490_),
    .B1(net4236),
    .B2(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .A2(net4252),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[27] ));
 sg13g2_nand3_1 _12803_ (.B(_07489_),
    .C(_07490_),
    .A(_07488_),
    .Y(_07491_));
 sg13g2_a22oi_1 _12804_ (.Y(_07492_),
    .B1(_07487_),
    .B2(_07491_),
    .A2(_07486_),
    .A1(net4625));
 sg13g2_nor2_1 _12805_ (.A(net1475),
    .B(net4634),
    .Y(_07493_));
 sg13g2_a21oi_1 _12806_ (.A1(net4634),
    .A2(net3895),
    .Y(_00497_),
    .B1(_07493_));
 sg13g2_a21oi_2 _12807_ (.B1(net4085),
    .Y(_07494_),
    .A2(net4620),
    .A1(\soc_inst.core_mem_rdata[28] ));
 sg13g2_a22oi_1 _12808_ (.Y(_07495_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[28] ),
    .A2(net4099),
    .A1(\soc_inst.cpu_core.csr_file.mcause[28] ));
 sg13g2_nand2_1 _12809_ (.Y(_07496_),
    .A(\soc_inst.cpu_core.csr_file.mstatus[28] ),
    .B(net4252));
 sg13g2_a22oi_1 _12810_ (.Y(_07497_),
    .B1(_06716_),
    .B2(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .A2(net4182),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[28] ));
 sg13g2_nand4_1 _12811_ (.B(_07495_),
    .C(_07496_),
    .A(net4248),
    .Y(_07498_),
    .D(_07497_));
 sg13g2_o21ai_1 _12812_ (.B1(_07498_),
    .Y(_07499_),
    .A1(\soc_inst.core_mem_addr[28] ),
    .A2(net4247));
 sg13g2_mux2_1 _12813_ (.A0(_07494_),
    .A1(_07499_),
    .S(_07216_),
    .X(_07500_));
 sg13g2_nor2_1 _12814_ (.A(net795),
    .B(net4631),
    .Y(_07501_));
 sg13g2_a21oi_1 _12815_ (.A1(net4631),
    .A2(net3821),
    .Y(_00498_),
    .B1(_07501_));
 sg13g2_a21oi_2 _12816_ (.B1(net4085),
    .Y(_07502_),
    .A2(net4619),
    .A1(\soc_inst.core_mem_rdata[29] ));
 sg13g2_a22oi_1 _12817_ (.Y(_07503_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[29] ),
    .A2(net4097),
    .A1(\soc_inst.cpu_core.csr_file.mcause[29] ));
 sg13g2_nand2_1 _12818_ (.Y(_07504_),
    .A(\soc_inst.cpu_core.csr_file.mstatus[29] ),
    .B(net4252));
 sg13g2_a22oi_1 _12819_ (.Y(_07505_),
    .B1(net4232),
    .B2(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .A2(net4181),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[29] ));
 sg13g2_nand4_1 _12820_ (.B(_07503_),
    .C(_07504_),
    .A(net4248),
    .Y(_07506_),
    .D(_07505_));
 sg13g2_o21ai_1 _12821_ (.B1(_07506_),
    .Y(_07507_),
    .A1(\soc_inst.core_mem_addr[29] ),
    .A2(net4247));
 sg13g2_mux2_1 _12822_ (.A0(_07502_),
    .A1(_07507_),
    .S(_07216_),
    .X(_07508_));
 sg13g2_nor2_1 _12823_ (.A(net1038),
    .B(net4634),
    .Y(_07509_));
 sg13g2_a21oi_1 _12824_ (.A1(net4634),
    .A2(net3820),
    .Y(_00499_),
    .B1(_07509_));
 sg13g2_a21o_1 _12825_ (.A2(net4621),
    .A1(\soc_inst.core_mem_rdata[30] ),
    .B1(net4087),
    .X(_07510_));
 sg13g2_a21oi_1 _12826_ (.A1(_05434_),
    .A2(net4242),
    .Y(_07511_),
    .B1(net4627));
 sg13g2_a22oi_1 _12827_ (.Y(_07512_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[30] ),
    .A2(net4097),
    .A1(\soc_inst.cpu_core.csr_file.mcause[30] ));
 sg13g2_a22oi_1 _12828_ (.Y(_07513_),
    .B1(net4181),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[30] ),
    .A2(net4254),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[30] ));
 sg13g2_nand2_1 _12829_ (.Y(_07514_),
    .A(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .B(net4236));
 sg13g2_nand4_1 _12830_ (.B(_07512_),
    .C(_07513_),
    .A(_07240_),
    .Y(_07515_),
    .D(_07514_));
 sg13g2_a22oi_1 _12831_ (.Y(_07516_),
    .B1(_07511_),
    .B2(_07515_),
    .A2(_07510_),
    .A1(net4629));
 sg13g2_nor2_1 _12832_ (.A(net1113),
    .B(net4638),
    .Y(_07517_));
 sg13g2_a21oi_1 _12833_ (.A1(net4638),
    .A2(net3893),
    .Y(_00500_),
    .B1(_07517_));
 sg13g2_a21oi_2 _12834_ (.B1(net4086),
    .Y(_07518_),
    .A2(net4620),
    .A1(\soc_inst.core_mem_rdata[31] ));
 sg13g2_a22oi_1 _12835_ (.Y(_07519_),
    .B1(net4092),
    .B2(\soc_inst.cpu_core.csr_file.mtval[31] ),
    .A2(net4099),
    .A1(\soc_inst.cpu_core.csr_file.mcause[31] ));
 sg13g2_nand2_1 _12836_ (.Y(_07520_),
    .A(\soc_inst.cpu_core.csr_file.mstatus[31] ),
    .B(net4254));
 sg13g2_a22oi_1 _12837_ (.Y(_07521_),
    .B1(net4232),
    .B2(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .A2(net4181),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[31] ));
 sg13g2_nand4_1 _12838_ (.B(_07519_),
    .C(_07520_),
    .A(net4248),
    .Y(_07522_),
    .D(_07521_));
 sg13g2_o21ai_1 _12839_ (.B1(_07522_),
    .Y(_07523_),
    .A1(\soc_inst.core_mem_addr[31] ),
    .A2(net4247));
 sg13g2_mux2_1 _12840_ (.A0(_07518_),
    .A1(_07523_),
    .S(_07216_),
    .X(_07524_));
 sg13g2_nor2_1 _12841_ (.A(net797),
    .B(net4632),
    .Y(_07525_));
 sg13g2_a21oi_1 _12842_ (.A1(net4632),
    .A2(net3818),
    .Y(_00501_),
    .B1(_07525_));
 sg13g2_nor2_1 _12843_ (.A(_07120_),
    .B(_07130_),
    .Y(_07526_));
 sg13g2_mux2_1 _12844_ (.A0(net1999),
    .A1(net5049),
    .S(_07526_),
    .X(_00502_));
 sg13g2_nor2_2 _12845_ (.A(_06592_),
    .B(_07130_),
    .Y(_07527_));
 sg13g2_mux2_1 _12846_ (.A0(net1944),
    .A1(net5049),
    .S(_07527_),
    .X(_00503_));
 sg13g2_mux2_1 _12847_ (.A0(net1753),
    .A1(net5045),
    .S(_07527_),
    .X(_00504_));
 sg13g2_mux2_1 _12848_ (.A0(net2592),
    .A1(net5043),
    .S(_07527_),
    .X(_00505_));
 sg13g2_mux2_1 _12849_ (.A0(net1827),
    .A1(net5040),
    .S(_07527_),
    .X(_00506_));
 sg13g2_mux2_1 _12850_ (.A0(net1909),
    .A1(net5037),
    .S(_07527_),
    .X(_00507_));
 sg13g2_mux2_1 _12851_ (.A0(net1854),
    .A1(net5034),
    .S(_07527_),
    .X(_00508_));
 sg13g2_mux2_1 _12852_ (.A0(net1591),
    .A1(net5031),
    .S(_07527_),
    .X(_00509_));
 sg13g2_nor2_2 _12853_ (.A(_06298_),
    .B(_07130_),
    .Y(_07528_));
 sg13g2_mux2_1 _12854_ (.A0(net2150),
    .A1(net5049),
    .S(_07528_),
    .X(_00510_));
 sg13g2_mux2_1 _12855_ (.A0(net2178),
    .A1(net5045),
    .S(_07528_),
    .X(_00511_));
 sg13g2_mux2_1 _12856_ (.A0(net2101),
    .A1(net5043),
    .S(_07528_),
    .X(_00512_));
 sg13g2_mux2_1 _12857_ (.A0(net2409),
    .A1(net5039),
    .S(_07528_),
    .X(_00513_));
 sg13g2_mux2_1 _12858_ (.A0(net1969),
    .A1(net5037),
    .S(_07528_),
    .X(_00514_));
 sg13g2_mux2_1 _12859_ (.A0(net2169),
    .A1(net5034),
    .S(_07528_),
    .X(_00515_));
 sg13g2_mux2_1 _12860_ (.A0(net2211),
    .A1(net5031),
    .S(_07528_),
    .X(_00516_));
 sg13g2_a21oi_2 _12861_ (.B1(_05907_),
    .Y(_07529_),
    .A2(_05948_),
    .A1(_05866_));
 sg13g2_nand2b_2 _12862_ (.Y(_07530_),
    .B(_00276_),
    .A_N(\soc_inst.mem_ctrl.access_state[4] ));
 sg13g2_nand2_1 _12863_ (.Y(_07531_),
    .A(_07529_),
    .B(_07530_));
 sg13g2_nor2_2 _12864_ (.A(\soc_inst.mem_ctrl.access_state[4] ),
    .B(_05869_),
    .Y(_07532_));
 sg13g2_nand2b_2 _12865_ (.Y(_07533_),
    .B(_05870_),
    .A_N(net2748));
 sg13g2_nor3_1 _12866_ (.A(net4711),
    .B(net3767),
    .C(_07533_),
    .Y(_07534_));
 sg13g2_a21o_1 _12867_ (.A2(net3767),
    .A1(net2759),
    .B1(_07534_),
    .X(_00517_));
 sg13g2_nor3_1 _12868_ (.A(_06750_),
    .B(net3767),
    .C(_07533_),
    .Y(_07535_));
 sg13g2_a21o_1 _12869_ (.A2(net3767),
    .A1(net2741),
    .B1(_07535_),
    .X(_00518_));
 sg13g2_nor3_1 _12870_ (.A(net4616),
    .B(net3767),
    .C(_07533_),
    .Y(_07536_));
 sg13g2_a21o_1 _12871_ (.A2(net3767),
    .A1(net2723),
    .B1(_07536_),
    .X(_00519_));
 sg13g2_a221oi_1 _12872_ (.B2(net4773),
    .C1(_05908_),
    .B1(_05946_),
    .A1(\soc_inst.mem_ctrl.access_state[3] ),
    .Y(_07537_),
    .A2(_05470_));
 sg13g2_nand2_1 _12873_ (.Y(_07538_),
    .A(_07529_),
    .B(_07537_));
 sg13g2_nor2_1 _12874_ (.A(_00276_),
    .B(_05869_),
    .Y(_07539_));
 sg13g2_nand2_1 _12875_ (.Y(_07540_),
    .A(_05467_),
    .B(_05469_));
 sg13g2_nor2_1 _12876_ (.A(net4773),
    .B(_07530_),
    .Y(_07541_));
 sg13g2_nor2_1 _12877_ (.A(_07530_),
    .B(_07540_),
    .Y(_07542_));
 sg13g2_nor3_1 _12878_ (.A(net4779),
    .B(_07530_),
    .C(_07540_),
    .Y(_07543_));
 sg13g2_nor4_1 _12879_ (.A(_06014_),
    .B(_07538_),
    .C(_07539_),
    .D(_07543_),
    .Y(_07544_));
 sg13g2_nor2_1 _12880_ (.A(_06015_),
    .B(_06026_),
    .Y(_07545_));
 sg13g2_a21oi_1 _12881_ (.A1(_07544_),
    .A2(_07545_),
    .Y(_07546_),
    .B1(net403));
 sg13g2_a21oi_1 _12882_ (.A1(_05466_),
    .A2(_07544_),
    .Y(_00520_),
    .B1(net404));
 sg13g2_nor2_1 _12883_ (.A(_06675_),
    .B(_07533_),
    .Y(_07547_));
 sg13g2_a21oi_1 _12884_ (.A1(\soc_inst.core_mem_wdata[24] ),
    .A2(net4175),
    .Y(_07548_),
    .B1(net3773));
 sg13g2_a21oi_1 _12885_ (.A1(_05841_),
    .A2(net3773),
    .Y(_00521_),
    .B1(_07548_));
 sg13g2_nand2_1 _12886_ (.Y(_07549_),
    .A(\soc_inst.core_mem_wdata[25] ),
    .B(net4175));
 sg13g2_nand2_1 _12887_ (.Y(_07550_),
    .A(net465),
    .B(net3773));
 sg13g2_o21ai_1 _12888_ (.B1(_07550_),
    .Y(_00522_),
    .A1(net3773),
    .A2(_07549_));
 sg13g2_nand2_1 _12889_ (.Y(_07551_),
    .A(\soc_inst.core_mem_wdata[26] ),
    .B(net4175));
 sg13g2_nand2_1 _12890_ (.Y(_07552_),
    .A(net389),
    .B(net3774));
 sg13g2_o21ai_1 _12891_ (.B1(_07552_),
    .Y(_00523_),
    .A1(net3775),
    .A2(_07551_));
 sg13g2_nand2_1 _12892_ (.Y(_07553_),
    .A(net480),
    .B(net4175));
 sg13g2_nand2_1 _12893_ (.Y(_07554_),
    .A(net588),
    .B(net3774));
 sg13g2_o21ai_1 _12894_ (.B1(_07554_),
    .Y(_00524_),
    .A1(net3775),
    .A2(_07553_));
 sg13g2_nand2_1 _12895_ (.Y(_07555_),
    .A(\soc_inst.core_mem_wdata[28] ),
    .B(net4175));
 sg13g2_nand2_1 _12896_ (.Y(_07556_),
    .A(net530),
    .B(net3773));
 sg13g2_o21ai_1 _12897_ (.B1(_07556_),
    .Y(_00525_),
    .A1(net3773),
    .A2(_07555_));
 sg13g2_nand2_1 _12898_ (.Y(_07557_),
    .A(\soc_inst.core_mem_wdata[29] ),
    .B(net4176));
 sg13g2_nand2_1 _12899_ (.Y(_07558_),
    .A(net427),
    .B(net3770));
 sg13g2_o21ai_1 _12900_ (.B1(_07558_),
    .Y(_00526_),
    .A1(net3770),
    .A2(_07557_));
 sg13g2_nand2_1 _12901_ (.Y(_07559_),
    .A(net383),
    .B(net4176));
 sg13g2_nand2_1 _12902_ (.Y(_07560_),
    .A(net429),
    .B(net3770));
 sg13g2_o21ai_1 _12903_ (.B1(_07560_),
    .Y(_00527_),
    .A1(net3770),
    .A2(_07559_));
 sg13g2_nand2_1 _12904_ (.Y(_07561_),
    .A(\soc_inst.core_mem_wdata[31] ),
    .B(net4174));
 sg13g2_nand2_1 _12905_ (.Y(_07562_),
    .A(net412),
    .B(net3770));
 sg13g2_o21ai_1 _12906_ (.B1(_07562_),
    .Y(_00528_),
    .A1(net3770),
    .A2(_07561_));
 sg13g2_nand2_1 _12907_ (.Y(_07563_),
    .A(\soc_inst.core_mem_wdata[16] ),
    .B(net4174));
 sg13g2_nand2_1 _12908_ (.Y(_07564_),
    .A(net671),
    .B(net3771));
 sg13g2_o21ai_1 _12909_ (.B1(_07564_),
    .Y(_00529_),
    .A1(net3771),
    .A2(_07563_));
 sg13g2_nand2_1 _12910_ (.Y(_07565_),
    .A(\soc_inst.core_mem_wdata[17] ),
    .B(net4175));
 sg13g2_nand2_1 _12911_ (.Y(_07566_),
    .A(net565),
    .B(net3775));
 sg13g2_o21ai_1 _12912_ (.B1(_07566_),
    .Y(_00530_),
    .A1(net3775),
    .A2(_07565_));
 sg13g2_nand2_1 _12913_ (.Y(_07567_),
    .A(\soc_inst.core_mem_wdata[18] ),
    .B(net4174));
 sg13g2_nand2_1 _12914_ (.Y(_07568_),
    .A(net778),
    .B(net3771));
 sg13g2_o21ai_1 _12915_ (.B1(_07568_),
    .Y(_00531_),
    .A1(net3771),
    .A2(_07567_));
 sg13g2_nand2_1 _12916_ (.Y(_07569_),
    .A(\soc_inst.core_mem_wdata[19] ),
    .B(net4174));
 sg13g2_nand2_1 _12917_ (.Y(_07570_),
    .A(net360),
    .B(net3771));
 sg13g2_o21ai_1 _12918_ (.B1(_07570_),
    .Y(_00532_),
    .A1(net3772),
    .A2(_07569_));
 sg13g2_nand2_1 _12919_ (.Y(_07571_),
    .A(\soc_inst.core_mem_wdata[20] ),
    .B(net4174));
 sg13g2_nand2_1 _12920_ (.Y(_07572_),
    .A(net580),
    .B(net3771));
 sg13g2_o21ai_1 _12921_ (.B1(_07572_),
    .Y(_00533_),
    .A1(net3772),
    .A2(_07571_));
 sg13g2_nand2_1 _12922_ (.Y(_07573_),
    .A(\soc_inst.core_mem_wdata[21] ),
    .B(net4174));
 sg13g2_nand2_1 _12923_ (.Y(_07574_),
    .A(net557),
    .B(net3771));
 sg13g2_o21ai_1 _12924_ (.B1(_07574_),
    .Y(_00534_),
    .A1(net3771),
    .A2(_07573_));
 sg13g2_nand2_1 _12925_ (.Y(_07575_),
    .A(\soc_inst.core_mem_wdata[22] ),
    .B(net4174));
 sg13g2_nand2_1 _12926_ (.Y(_07576_),
    .A(net534),
    .B(net3772));
 sg13g2_o21ai_1 _12927_ (.B1(_07576_),
    .Y(_00535_),
    .A1(net3772),
    .A2(_07575_));
 sg13g2_nand2_1 _12928_ (.Y(_07577_),
    .A(\soc_inst.core_mem_wdata[23] ),
    .B(net4174));
 sg13g2_nand2_1 _12929_ (.Y(_07578_),
    .A(net488),
    .B(net3772));
 sg13g2_o21ai_1 _12930_ (.B1(_07578_),
    .Y(_00536_),
    .A1(net3772),
    .A2(_07577_));
 sg13g2_nor2_2 _12931_ (.A(_06676_),
    .B(_07533_),
    .Y(_07579_));
 sg13g2_a21oi_1 _12932_ (.A1(net5027),
    .A2(_07579_),
    .Y(_07580_),
    .B1(net3773));
 sg13g2_a21oi_1 _12933_ (.A1(_05850_),
    .A2(net3774),
    .Y(_00537_),
    .B1(_07580_));
 sg13g2_a21oi_1 _12934_ (.A1(net5025),
    .A2(_07579_),
    .Y(_07581_),
    .B1(net3770));
 sg13g2_a21oi_1 _12935_ (.A1(_05852_),
    .A2(net3770),
    .Y(_00538_),
    .B1(_07581_));
 sg13g2_a21oi_1 _12936_ (.A1(\soc_inst.core_mem_wdata[10] ),
    .A2(_07579_),
    .Y(_07582_),
    .B1(net3774));
 sg13g2_a21oi_1 _12937_ (.A1(_05853_),
    .A2(net3774),
    .Y(_00539_),
    .B1(_07582_));
 sg13g2_a21oi_1 _12938_ (.A1(\soc_inst.core_mem_wdata[11] ),
    .A2(_07579_),
    .Y(_07583_),
    .B1(net3773));
 sg13g2_a21oi_1 _12939_ (.A1(_05855_),
    .A2(net3778),
    .Y(_00540_),
    .B1(_07583_));
 sg13g2_a21oi_1 _12940_ (.A1(net5021),
    .A2(_07579_),
    .Y(_07584_),
    .B1(net3777));
 sg13g2_a21oi_1 _12941_ (.A1(_05857_),
    .A2(net3777),
    .Y(_00541_),
    .B1(_07584_));
 sg13g2_a21oi_1 _12942_ (.A1(\soc_inst.core_mem_wdata[13] ),
    .A2(_07579_),
    .Y(_07585_),
    .B1(net3774));
 sg13g2_a21oi_1 _12943_ (.A1(_05858_),
    .A2(net3774),
    .Y(_00542_),
    .B1(_07585_));
 sg13g2_a21oi_1 _12944_ (.A1(\soc_inst.core_mem_wdata[14] ),
    .A2(_07579_),
    .Y(_07586_),
    .B1(net3777));
 sg13g2_a21oi_1 _12945_ (.A1(_05859_),
    .A2(net3777),
    .Y(_00543_),
    .B1(_07586_));
 sg13g2_a21oi_1 _12946_ (.A1(net5018),
    .A2(_07579_),
    .Y(_07587_),
    .B1(net3777));
 sg13g2_a21oi_1 _12947_ (.A1(_05861_),
    .A2(net3777),
    .Y(_00544_),
    .B1(_07587_));
 sg13g2_nand2_1 _12948_ (.Y(_07588_),
    .A(net5050),
    .B(_07532_));
 sg13g2_nand2_1 _12949_ (.Y(_07589_),
    .A(net296),
    .B(net3768));
 sg13g2_o21ai_1 _12950_ (.B1(_07589_),
    .Y(_00545_),
    .A1(net3768),
    .A2(_07588_));
 sg13g2_nand2_1 _12951_ (.Y(_07590_),
    .A(\soc_inst.core_mem_wdata[1] ),
    .B(_07532_));
 sg13g2_nand2_1 _12952_ (.Y(_07591_),
    .A(net327),
    .B(net3768));
 sg13g2_o21ai_1 _12953_ (.B1(_07591_),
    .Y(_00546_),
    .A1(net3769),
    .A2(_07590_));
 sg13g2_nand2_1 _12954_ (.Y(_07592_),
    .A(\soc_inst.core_mem_wdata[2] ),
    .B(_07532_));
 sg13g2_nand2_1 _12955_ (.Y(_07593_),
    .A(net313),
    .B(net3777));
 sg13g2_o21ai_1 _12956_ (.B1(_07593_),
    .Y(_00547_),
    .A1(net3768),
    .A2(_07592_));
 sg13g2_nand2_1 _12957_ (.Y(_07594_),
    .A(\soc_inst.core_mem_wdata[3] ),
    .B(_07532_));
 sg13g2_nand2_1 _12958_ (.Y(_07595_),
    .A(net213),
    .B(net3769));
 sg13g2_o21ai_1 _12959_ (.B1(_07595_),
    .Y(_00548_),
    .A1(net3768),
    .A2(_07594_));
 sg13g2_nand2_1 _12960_ (.Y(_07596_),
    .A(\soc_inst.core_mem_wdata[4] ),
    .B(_07532_));
 sg13g2_nand2_1 _12961_ (.Y(_07597_),
    .A(net264),
    .B(net3768));
 sg13g2_o21ai_1 _12962_ (.B1(_07597_),
    .Y(_00549_),
    .A1(net3769),
    .A2(_07596_));
 sg13g2_nand2_1 _12963_ (.Y(_07598_),
    .A(\soc_inst.core_mem_wdata[5] ),
    .B(_07532_));
 sg13g2_nand2_1 _12964_ (.Y(_07599_),
    .A(net226),
    .B(net3768));
 sg13g2_o21ai_1 _12965_ (.B1(_07599_),
    .Y(_00550_),
    .A1(net3768),
    .A2(_07598_));
 sg13g2_nand2_1 _12966_ (.Y(_07600_),
    .A(\soc_inst.core_mem_wdata[6] ),
    .B(_07532_));
 sg13g2_nand2_1 _12967_ (.Y(_07601_),
    .A(net277),
    .B(net3769));
 sg13g2_o21ai_1 _12968_ (.B1(_07601_),
    .Y(_00551_),
    .A1(net3769),
    .A2(_07600_));
 sg13g2_nand2_1 _12969_ (.Y(_07602_),
    .A(net5030),
    .B(_07532_));
 sg13g2_nand2_1 _12970_ (.Y(_07603_),
    .A(net354),
    .B(net3767));
 sg13g2_o21ai_1 _12971_ (.B1(_07603_),
    .Y(_00552_),
    .A1(net3767),
    .A2(_07602_));
 sg13g2_nand2_1 _12972_ (.Y(_07604_),
    .A(net4753),
    .B(_06738_));
 sg13g2_o21ai_1 _12973_ (.B1(net4616),
    .Y(_07605_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .A2(net4609));
 sg13g2_o21ai_1 _12974_ (.B1(_06750_),
    .Y(_07606_),
    .A1(net4755),
    .A2(net4869));
 sg13g2_nand3_1 _12975_ (.B(net4248),
    .C(_07606_),
    .A(net4256),
    .Y(_07607_));
 sg13g2_o21ai_1 _12976_ (.B1(net470),
    .Y(_07608_),
    .A1(_07605_),
    .A2(net4173));
 sg13g2_nor2b_1 _12977_ (.A(net4870),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .Y(_07609_));
 sg13g2_nor2_2 _12978_ (.A(net4868),
    .B(net4231),
    .Y(_07610_));
 sg13g2_nand2_1 _12979_ (.Y(_07611_),
    .A(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .B(net4169));
 sg13g2_o21ai_1 _12980_ (.B1(_07608_),
    .Y(_00553_),
    .A1(net4173),
    .A2(_07611_));
 sg13g2_o21ai_1 _12981_ (.B1(net4616),
    .Y(_07612_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .A2(net4610));
 sg13g2_o21ai_1 _12982_ (.B1(net446),
    .Y(_07613_),
    .A1(net4173),
    .A2(_07612_));
 sg13g2_nor2b_1 _12983_ (.A(net4870),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .Y(_07614_));
 sg13g2_nand2_1 _12984_ (.Y(_07615_),
    .A(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .B(net4169));
 sg13g2_o21ai_1 _12985_ (.B1(_07613_),
    .Y(_00554_),
    .A1(net4173),
    .A2(_07615_));
 sg13g2_o21ai_1 _12986_ (.B1(net4616),
    .Y(_07616_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .A2(net4610));
 sg13g2_o21ai_1 _12987_ (.B1(net434),
    .Y(_07617_),
    .A1(net4173),
    .A2(_07616_));
 sg13g2_nor2b_1 _12988_ (.A(net4869),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .Y(_07618_));
 sg13g2_nand2_1 _12989_ (.Y(_07619_),
    .A(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .B(net4169));
 sg13g2_o21ai_1 _12990_ (.B1(_07617_),
    .Y(_00555_),
    .A1(net4173),
    .A2(_07619_));
 sg13g2_o21ai_1 _12991_ (.B1(net4616),
    .Y(_07620_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .A2(net4610));
 sg13g2_o21ai_1 _12992_ (.B1(net478),
    .Y(_07621_),
    .A1(net4173),
    .A2(_07620_));
 sg13g2_nor2b_1 _12993_ (.A(net4869),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .Y(_07622_));
 sg13g2_nand2_1 _12994_ (.Y(_07623_),
    .A(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .B(net4169));
 sg13g2_o21ai_1 _12995_ (.B1(_07621_),
    .Y(_00556_),
    .A1(net4173),
    .A2(_07623_));
 sg13g2_o21ai_1 _12996_ (.B1(net4616),
    .Y(_07624_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .A2(net4610));
 sg13g2_o21ai_1 _12997_ (.B1(net462),
    .Y(_07625_),
    .A1(_07607_),
    .A2(_07624_));
 sg13g2_nor2b_1 _12998_ (.A(net4869),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .Y(_07626_));
 sg13g2_nand2_1 _12999_ (.Y(_07627_),
    .A(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .B(net4170));
 sg13g2_o21ai_1 _13000_ (.B1(net463),
    .Y(_00557_),
    .A1(_07607_),
    .A2(_07627_));
 sg13g2_a21oi_1 _13001_ (.A1(_06670_),
    .A2(net4177),
    .Y(_07628_),
    .B1(_06696_));
 sg13g2_nor2b_1 _13002_ (.A(_06732_),
    .B_N(_07628_),
    .Y(_07629_));
 sg13g2_nor2_1 _13003_ (.A(net1559),
    .B(net3764),
    .Y(_07630_));
 sg13g2_nand2b_1 _13004_ (.Y(_07631_),
    .B(_06754_),
    .A_N(net1559));
 sg13g2_nor2_1 _13005_ (.A(net4872),
    .B(_06754_),
    .Y(_07632_));
 sg13g2_a21oi_1 _13006_ (.A1(_06757_),
    .A2(_07631_),
    .Y(_07633_),
    .B1(_07632_));
 sg13g2_a21oi_1 _13007_ (.A1(net3764),
    .A2(_07633_),
    .Y(_00558_),
    .B1(_07630_));
 sg13g2_nor2_1 _13008_ (.A(net752),
    .B(net3765),
    .Y(_07634_));
 sg13g2_nand2_1 _13009_ (.Y(_07635_),
    .A(_05613_),
    .B(_06766_));
 sg13g2_nor2_1 _13010_ (.A(net4872),
    .B(_06766_),
    .Y(_07636_));
 sg13g2_a21oi_1 _13011_ (.A1(_06769_),
    .A2(_07635_),
    .Y(_07637_),
    .B1(_07636_));
 sg13g2_a21oi_1 _13012_ (.A1(net3765),
    .A2(_07637_),
    .Y(_00559_),
    .B1(_07634_));
 sg13g2_nor2_1 _13013_ (.A(net1605),
    .B(net3764),
    .Y(_07638_));
 sg13g2_nand2b_1 _13014_ (.Y(_07639_),
    .B(_06774_),
    .A_N(net1605));
 sg13g2_nor2_1 _13015_ (.A(net4871),
    .B(_06774_),
    .Y(_07640_));
 sg13g2_a21oi_1 _13016_ (.A1(_06777_),
    .A2(_07639_),
    .Y(_07641_),
    .B1(_07640_));
 sg13g2_a21oi_1 _13017_ (.A1(net3764),
    .A2(_07641_),
    .Y(_00560_),
    .B1(_07638_));
 sg13g2_a21oi_1 _13018_ (.A1(_06741_),
    .A2(net3764),
    .Y(_07642_),
    .B1(net499));
 sg13g2_a21oi_1 _13019_ (.A1(_06743_),
    .A2(net3764),
    .Y(_00561_),
    .B1(_07642_));
 sg13g2_nor2_1 _13020_ (.A(net1533),
    .B(net3764),
    .Y(_07643_));
 sg13g2_nand2b_1 _13021_ (.Y(_07644_),
    .B(_06787_),
    .A_N(net1533));
 sg13g2_nor2_1 _13022_ (.A(net4872),
    .B(_06787_),
    .Y(_07645_));
 sg13g2_a21oi_1 _13023_ (.A1(_06790_),
    .A2(_07644_),
    .Y(_07646_),
    .B1(_07645_));
 sg13g2_a21oi_1 _13024_ (.A1(net3764),
    .A2(_07646_),
    .Y(_00562_),
    .B1(_07643_));
 sg13g2_o21ai_1 _13025_ (.B1(net4274),
    .Y(_07647_),
    .A1(_07140_),
    .A2(_07154_));
 sg13g2_nand2_1 _13026_ (.Y(_07648_),
    .A(_06974_),
    .B(_07164_));
 sg13g2_o21ai_1 _13027_ (.B1(net4275),
    .Y(_07649_),
    .A1(_07172_),
    .A2(_07648_));
 sg13g2_nor2b_1 _13028_ (.A(_06966_),
    .B_N(_07647_),
    .Y(_07650_));
 sg13g2_and2_1 _13029_ (.A(_07649_),
    .B(_07650_),
    .X(_07651_));
 sg13g2_o21ai_1 _13030_ (.B1(_07651_),
    .Y(_07652_),
    .A1(\soc_inst.i2c_inst.stop_pending ),
    .A2(_06963_));
 sg13g2_nand2b_1 _13031_ (.Y(_07653_),
    .B(\soc_inst.i2c_inst.bit_cnt[3] ),
    .A_N(\soc_inst.i2c_inst.bit_cnt[2] ));
 sg13g2_nor4_1 _13032_ (.A(\soc_inst.i2c_inst.bit_cnt[0] ),
    .B(\soc_inst.i2c_inst.bit_cnt[1] ),
    .C(_06975_),
    .D(_07653_),
    .Y(_07654_));
 sg13g2_o21ai_1 _13033_ (.B1(_06927_),
    .Y(_07655_),
    .A1(net824),
    .A2(\soc_inst.i2c_inst.restart_pending ));
 sg13g2_nor3_1 _13034_ (.A(_06022_),
    .B(_07170_),
    .C(_07654_),
    .Y(_07656_));
 sg13g2_nand2_1 _13035_ (.Y(_07657_),
    .A(_07655_),
    .B(_07656_));
 sg13g2_mux2_1 _13036_ (.A0(_07657_),
    .A1(net2175),
    .S(_07652_),
    .X(_00563_));
 sg13g2_nand2b_1 _13037_ (.Y(_07658_),
    .B(_06927_),
    .A_N(net824));
 sg13g2_a221oi_1 _13038_ (.B2(_06416_),
    .C1(_07154_),
    .B1(_07155_),
    .A1(_05471_),
    .Y(_07659_),
    .A2(_06439_));
 sg13g2_o21ai_1 _13039_ (.B1(_07659_),
    .Y(_07660_),
    .A1(_05864_),
    .A2(_07658_));
 sg13g2_nor2_1 _13040_ (.A(_07652_),
    .B(_07660_),
    .Y(_07661_));
 sg13g2_a21oi_1 _13041_ (.A1(_05471_),
    .A2(_07652_),
    .Y(_00564_),
    .B1(_07661_));
 sg13g2_nand4_1 _13042_ (.B(_06975_),
    .C(_07164_),
    .A(_06442_),
    .Y(_07662_),
    .D(_07658_));
 sg13g2_mux2_1 _13043_ (.A0(_07662_),
    .A1(net5118),
    .S(_07652_),
    .X(_00565_));
 sg13g2_a22oi_1 _13044_ (.Y(_07663_),
    .B1(_07155_),
    .B2(_06416_),
    .A2(_06927_),
    .A1(net824));
 sg13g2_nand2_1 _13045_ (.Y(_07664_),
    .A(_07156_),
    .B(_07663_));
 sg13g2_mux2_1 _13046_ (.A0(_07664_),
    .A1(net5116),
    .S(_07652_),
    .X(_00566_));
 sg13g2_nor2_1 _13047_ (.A(_06014_),
    .B(_06032_),
    .Y(_07665_));
 sg13g2_a21oi_1 _13048_ (.A1(net4772),
    .A2(_05946_),
    .Y(_07666_),
    .B1(_07541_));
 sg13g2_and3_1 _13049_ (.X(_07667_),
    .A(_07529_),
    .B(_07665_),
    .C(_07666_));
 sg13g2_o21ai_1 _13050_ (.B1(_05467_),
    .Y(_07668_),
    .A1(\soc_inst.mem_ctrl.access_state[4] ),
    .A2(_05870_));
 sg13g2_nor2_1 _13051_ (.A(net4773),
    .B(_07533_),
    .Y(_07669_));
 sg13g2_a22oi_1 _13052_ (.Y(_07670_),
    .B1(net4163),
    .B2(\soc_inst.core_mem_addr[0] ),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[0] ));
 sg13g2_nor2_1 _13053_ (.A(net1907),
    .B(net3710),
    .Y(_07671_));
 sg13g2_a21oi_1 _13054_ (.A1(net3710),
    .A2(_07670_),
    .Y(_00567_),
    .B1(_07671_));
 sg13g2_a22oi_1 _13055_ (.Y(_07672_),
    .B1(net4165),
    .B2(\soc_inst.core_mem_addr[1] ),
    .A2(net4224),
    .A1(net2533));
 sg13g2_nor2_1 _13056_ (.A(net2699),
    .B(net3707),
    .Y(_07673_));
 sg13g2_a21oi_1 _13057_ (.A1(net3707),
    .A2(_07672_),
    .Y(_00568_),
    .B1(_07673_));
 sg13g2_a22oi_1 _13058_ (.Y(_07674_),
    .B1(net4163),
    .B2(net4799),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[2] ));
 sg13g2_nor2_1 _13059_ (.A(net2690),
    .B(net3708),
    .Y(_07675_));
 sg13g2_a21oi_1 _13060_ (.A1(net3708),
    .A2(_07674_),
    .Y(_00569_),
    .B1(_07675_));
 sg13g2_a22oi_1 _13061_ (.Y(_07676_),
    .B1(net4163),
    .B2(net4796),
    .A2(net4222),
    .A1(net2496));
 sg13g2_nor2_1 _13062_ (.A(net2572),
    .B(net3708),
    .Y(_07677_));
 sg13g2_a21oi_1 _13063_ (.A1(net3708),
    .A2(_07676_),
    .Y(_00570_),
    .B1(_07677_));
 sg13g2_a22oi_1 _13064_ (.Y(_07678_),
    .B1(net4163),
    .B2(\soc_inst.pwm_inst.channel_idx [0]),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[4] ));
 sg13g2_nor2_1 _13065_ (.A(net2503),
    .B(net3709),
    .Y(_07679_));
 sg13g2_a21oi_1 _13066_ (.A1(net3708),
    .A2(_07678_),
    .Y(_00571_),
    .B1(_07679_));
 sg13g2_a22oi_1 _13067_ (.Y(_07680_),
    .B1(net4163),
    .B2(net2017),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[5] ));
 sg13g2_nor2_1 _13068_ (.A(net2335),
    .B(net3709),
    .Y(_07681_));
 sg13g2_a21oi_1 _13069_ (.A1(net3708),
    .A2(_07680_),
    .Y(_00572_),
    .B1(_07681_));
 sg13g2_a22oi_1 _13070_ (.Y(_07682_),
    .B1(net4164),
    .B2(net1902),
    .A2(net4223),
    .A1(\soc_inst.core_instr_addr[6] ));
 sg13g2_nor2_1 _13071_ (.A(net2561),
    .B(net3709),
    .Y(_07683_));
 sg13g2_a21oi_1 _13072_ (.A1(net3709),
    .A2(_07682_),
    .Y(_00573_),
    .B1(_07683_));
 sg13g2_a22oi_1 _13073_ (.Y(_07684_),
    .B1(net4164),
    .B2(net1798),
    .A2(net4223),
    .A1(\soc_inst.core_instr_addr[7] ));
 sg13g2_nor2_1 _13074_ (.A(net2511),
    .B(net3708),
    .Y(_07685_));
 sg13g2_a21oi_1 _13075_ (.A1(net3708),
    .A2(_07684_),
    .Y(_00574_),
    .B1(_07685_));
 sg13g2_a22oi_1 _13076_ (.Y(_07686_),
    .B1(net4165),
    .B2(\soc_inst.core_mem_addr[8] ),
    .A2(net4224),
    .A1(\soc_inst.core_instr_addr[8] ));
 sg13g2_nor2_1 _13077_ (.A(net2494),
    .B(net3707),
    .Y(_07687_));
 sg13g2_a21oi_1 _13078_ (.A1(net3707),
    .A2(_07686_),
    .Y(_00575_),
    .B1(_07687_));
 sg13g2_a22oi_1 _13079_ (.Y(_07688_),
    .B1(net4166),
    .B2(net2371),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[9] ));
 sg13g2_nor2_1 _13080_ (.A(net2387),
    .B(net3705),
    .Y(_07689_));
 sg13g2_a21oi_1 _13081_ (.A1(net3704),
    .A2(_07688_),
    .Y(_00576_),
    .B1(_07689_));
 sg13g2_a22oi_1 _13082_ (.Y(_07690_),
    .B1(net4166),
    .B2(net2195),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[10] ));
 sg13g2_nor2_1 _13083_ (.A(net2326),
    .B(net3705),
    .Y(_07691_));
 sg13g2_a21oi_1 _13084_ (.A1(net3704),
    .A2(_07690_),
    .Y(_00577_),
    .B1(_07691_));
 sg13g2_a22oi_1 _13085_ (.Y(_07692_),
    .B1(net4166),
    .B2(net1807),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[11] ));
 sg13g2_nor2_1 _13086_ (.A(net2574),
    .B(net3705),
    .Y(_07693_));
 sg13g2_a21oi_1 _13087_ (.A1(net3704),
    .A2(_07692_),
    .Y(_00578_),
    .B1(_07693_));
 sg13g2_a22oi_1 _13088_ (.Y(_07694_),
    .B1(net4163),
    .B2(net4787),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[12] ));
 sg13g2_nor2_1 _13089_ (.A(net2570),
    .B(net3709),
    .Y(_07695_));
 sg13g2_a21oi_1 _13090_ (.A1(net3709),
    .A2(_07694_),
    .Y(_00579_),
    .B1(_07695_));
 sg13g2_a22oi_1 _13091_ (.Y(_07696_),
    .B1(net4163),
    .B2(\soc_inst.core_mem_addr[13] ),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[13] ));
 sg13g2_nor2_1 _13092_ (.A(net2526),
    .B(net3710),
    .Y(_07697_));
 sg13g2_a21oi_1 _13093_ (.A1(net3710),
    .A2(_07696_),
    .Y(_00580_),
    .B1(_07697_));
 sg13g2_a22oi_1 _13094_ (.Y(_07698_),
    .B1(net4163),
    .B2(\soc_inst.core_mem_addr[14] ),
    .A2(net4222),
    .A1(\soc_inst.core_instr_addr[14] ));
 sg13g2_nor2_1 _13095_ (.A(net2421),
    .B(net3711),
    .Y(_07699_));
 sg13g2_a21oi_1 _13096_ (.A1(net3710),
    .A2(_07698_),
    .Y(_00581_),
    .B1(_07699_));
 sg13g2_a22oi_1 _13097_ (.Y(_07700_),
    .B1(net4164),
    .B2(\soc_inst.core_mem_addr[15] ),
    .A2(net4223),
    .A1(\soc_inst.core_instr_addr[15] ));
 sg13g2_nor2_1 _13098_ (.A(net2507),
    .B(net3710),
    .Y(_07701_));
 sg13g2_a21oi_1 _13099_ (.A1(net3709),
    .A2(_07700_),
    .Y(_00582_),
    .B1(_07701_));
 sg13g2_a22oi_1 _13100_ (.Y(_07702_),
    .B1(net4165),
    .B2(net2515),
    .A2(net4224),
    .A1(\soc_inst.core_instr_addr[16] ));
 sg13g2_nor2_1 _13101_ (.A(net2685),
    .B(net3707),
    .Y(_07703_));
 sg13g2_a21oi_1 _13102_ (.A1(net3707),
    .A2(_07702_),
    .Y(_00583_),
    .B1(_07703_));
 sg13g2_a22oi_1 _13103_ (.Y(_07704_),
    .B1(net4165),
    .B2(\soc_inst.core_mem_addr[17] ),
    .A2(net4224),
    .A1(\soc_inst.core_instr_addr[17] ));
 sg13g2_nor2_1 _13104_ (.A(net2458),
    .B(net3707),
    .Y(_07705_));
 sg13g2_a21oi_1 _13105_ (.A1(net3706),
    .A2(_07704_),
    .Y(_00584_),
    .B1(_07705_));
 sg13g2_a22oi_1 _13106_ (.Y(_07706_),
    .B1(net4165),
    .B2(\soc_inst.core_mem_addr[18] ),
    .A2(net4224),
    .A1(\soc_inst.core_instr_addr[18] ));
 sg13g2_nor2_1 _13107_ (.A(net2624),
    .B(net3707),
    .Y(_07707_));
 sg13g2_a21oi_1 _13108_ (.A1(net3711),
    .A2(_07706_),
    .Y(_00585_),
    .B1(_07707_));
 sg13g2_a22oi_1 _13109_ (.Y(_07708_),
    .B1(net4165),
    .B2(\soc_inst.core_mem_addr[19] ),
    .A2(net4224),
    .A1(\soc_inst.core_instr_addr[19] ));
 sg13g2_nor2_1 _13110_ (.A(net2522),
    .B(net3706),
    .Y(_07709_));
 sg13g2_a21oi_1 _13111_ (.A1(net3706),
    .A2(_07708_),
    .Y(_00586_),
    .B1(_07709_));
 sg13g2_a22oi_1 _13112_ (.Y(_07710_),
    .B1(net4166),
    .B2(\soc_inst.core_mem_addr[20] ),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[20] ));
 sg13g2_nor2_1 _13113_ (.A(net2513),
    .B(net3706),
    .Y(_07711_));
 sg13g2_a21oi_1 _13114_ (.A1(net3705),
    .A2(_07710_),
    .Y(_00587_),
    .B1(_07711_));
 sg13g2_a22oi_1 _13115_ (.Y(_07712_),
    .B1(net4166),
    .B2(\soc_inst.core_mem_addr[21] ),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[21] ));
 sg13g2_nor2_1 _13116_ (.A(net2486),
    .B(net3705),
    .Y(_07713_));
 sg13g2_a21oi_1 _13117_ (.A1(net3704),
    .A2(_07712_),
    .Y(_00588_),
    .B1(_07713_));
 sg13g2_a22oi_1 _13118_ (.Y(_07714_),
    .B1(net4166),
    .B2(\soc_inst.core_mem_addr[22] ),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[22] ));
 sg13g2_nor2_1 _13119_ (.A(net1777),
    .B(net3704),
    .Y(_07715_));
 sg13g2_a21oi_1 _13120_ (.A1(net3704),
    .A2(_07714_),
    .Y(_00589_),
    .B1(_07715_));
 sg13g2_a22oi_1 _13121_ (.Y(_07716_),
    .B1(net4166),
    .B2(\soc_inst.core_mem_addr[23] ),
    .A2(net4225),
    .A1(\soc_inst.core_instr_addr[23] ));
 sg13g2_nor2_1 _13122_ (.A(net2427),
    .B(net3704),
    .Y(_07717_));
 sg13g2_a21oi_1 _13123_ (.A1(net3704),
    .A2(_07716_),
    .Y(_00590_),
    .B1(_07717_));
 sg13g2_nand4_1 _13124_ (.B(_07537_),
    .C(_07540_),
    .A(_05906_),
    .Y(_07718_),
    .D(_07665_));
 sg13g2_nand2b_1 _13125_ (.Y(_07719_),
    .B(net4770),
    .A_N(net241));
 sg13g2_o21ai_1 _13126_ (.B1(_07719_),
    .Y(_07720_),
    .A1(net4770),
    .A2(net2879));
 sg13g2_nand2_1 _13127_ (.Y(_07721_),
    .A(net5114),
    .B(net3703));
 sg13g2_o21ai_1 _13128_ (.B1(_07721_),
    .Y(_00591_),
    .A1(net3703),
    .A2(_07720_));
 sg13g2_nand2b_1 _13129_ (.Y(_07722_),
    .B(net4772),
    .A_N(net211));
 sg13g2_o21ai_1 _13130_ (.B1(_07722_),
    .Y(_07723_),
    .A1(net4772),
    .A2(\soc_inst.mem_ctrl.spi_data_out[25] ));
 sg13g2_nand2_1 _13131_ (.Y(_07724_),
    .A(net543),
    .B(net3703));
 sg13g2_o21ai_1 _13132_ (.B1(_07724_),
    .Y(_00592_),
    .A1(net3703),
    .A2(_07723_));
 sg13g2_nand2_1 _13133_ (.Y(_07725_),
    .A(net4768),
    .B(net202));
 sg13g2_o21ai_1 _13134_ (.B1(_07725_),
    .Y(_07726_),
    .A1(net4767),
    .A2(_05583_));
 sg13g2_mux2_1 _13135_ (.A0(_07726_),
    .A1(net5112),
    .S(net3698),
    .X(_00593_));
 sg13g2_nand2b_1 _13136_ (.Y(_07727_),
    .B(net4767),
    .A_N(net108));
 sg13g2_o21ai_1 _13137_ (.B1(_07727_),
    .Y(_07728_),
    .A1(net4767),
    .A2(\soc_inst.mem_ctrl.spi_data_out[27] ));
 sg13g2_nand2_1 _13138_ (.Y(_07729_),
    .A(net5110),
    .B(net3698));
 sg13g2_o21ai_1 _13139_ (.B1(_07729_),
    .Y(_00594_),
    .A1(net3698),
    .A2(_07728_));
 sg13g2_nand2b_1 _13140_ (.Y(_07730_),
    .B(net4767),
    .A_N(net106));
 sg13g2_o21ai_1 _13141_ (.B1(_07730_),
    .Y(_07731_),
    .A1(net4767),
    .A2(net2615));
 sg13g2_nand2_1 _13142_ (.Y(_07732_),
    .A(net5109),
    .B(net3698));
 sg13g2_o21ai_1 _13143_ (.B1(_07732_),
    .Y(_00595_),
    .A1(net3698),
    .A2(_07731_));
 sg13g2_nand2b_1 _13144_ (.Y(_07733_),
    .B(net4768),
    .A_N(net124));
 sg13g2_o21ai_1 _13145_ (.B1(_07733_),
    .Y(_07734_),
    .A1(net4768),
    .A2(\soc_inst.mem_ctrl.spi_data_out[29] ));
 sg13g2_nand2_1 _13146_ (.Y(_07735_),
    .A(net5107),
    .B(net3699));
 sg13g2_o21ai_1 _13147_ (.B1(_07735_),
    .Y(_00596_),
    .A1(net3699),
    .A2(_07734_));
 sg13g2_nand2b_1 _13148_ (.Y(_07736_),
    .B(net4768),
    .A_N(net182));
 sg13g2_o21ai_1 _13149_ (.B1(_07736_),
    .Y(_07737_),
    .A1(net4768),
    .A2(net2000));
 sg13g2_nand2_1 _13150_ (.Y(_07738_),
    .A(net5105),
    .B(net3700));
 sg13g2_o21ai_1 _13151_ (.B1(_07738_),
    .Y(_00597_),
    .A1(net3699),
    .A2(_07737_));
 sg13g2_nand2_1 _13152_ (.Y(_07739_),
    .A(net4768),
    .B(net282));
 sg13g2_o21ai_1 _13153_ (.B1(_07739_),
    .Y(_07740_),
    .A1(net4767),
    .A2(_05584_));
 sg13g2_mux2_1 _13154_ (.A0(_07740_),
    .A1(net5103),
    .S(net3698),
    .X(_00598_));
 sg13g2_nand2b_1 _13155_ (.Y(_07741_),
    .B(net4771),
    .A_N(net139));
 sg13g2_o21ai_1 _13156_ (.B1(_07741_),
    .Y(_07742_),
    .A1(net4771),
    .A2(net2677));
 sg13g2_nand2_1 _13157_ (.Y(_07743_),
    .A(net5101),
    .B(net3701));
 sg13g2_o21ai_1 _13158_ (.B1(_07743_),
    .Y(_00599_),
    .A1(net3702),
    .A2(_07742_));
 sg13g2_nand2b_1 _13159_ (.Y(_07744_),
    .B(net4769),
    .A_N(net332));
 sg13g2_o21ai_1 _13160_ (.B1(_07744_),
    .Y(_07745_),
    .A1(net4769),
    .A2(\soc_inst.mem_ctrl.spi_data_out[17] ));
 sg13g2_nand2_1 _13161_ (.Y(_07746_),
    .A(net947),
    .B(net3701));
 sg13g2_o21ai_1 _13162_ (.B1(_07746_),
    .Y(_00600_),
    .A1(net3701),
    .A2(_07745_));
 sg13g2_mux2_1 _13163_ (.A0(net2647),
    .A1(net179),
    .S(net4766),
    .X(_07747_));
 sg13g2_nor2_1 _13164_ (.A(net3698),
    .B(_07747_),
    .Y(_07748_));
 sg13g2_a21oi_1 _13165_ (.A1(_05649_),
    .A2(net3698),
    .Y(_00601_),
    .B1(_07748_));
 sg13g2_nand2b_1 _13166_ (.Y(_07749_),
    .B(net4771),
    .A_N(net200));
 sg13g2_o21ai_1 _13167_ (.B1(_07749_),
    .Y(_07750_),
    .A1(net4769),
    .A2(net2881));
 sg13g2_nand2_1 _13168_ (.Y(_07751_),
    .A(net5094),
    .B(net3701));
 sg13g2_o21ai_1 _13169_ (.B1(_07751_),
    .Y(_00602_),
    .A1(net3702),
    .A2(_07750_));
 sg13g2_mux2_1 _13170_ (.A0(net2848),
    .A1(net228),
    .S(net4769),
    .X(_07752_));
 sg13g2_nor2_1 _13171_ (.A(net3700),
    .B(_07752_),
    .Y(_07753_));
 sg13g2_a21oi_1 _13172_ (.A1(_05650_),
    .A2(net3700),
    .Y(_00603_),
    .B1(_07753_));
 sg13g2_nand2b_1 _13173_ (.Y(_07754_),
    .B(net4771),
    .A_N(net234));
 sg13g2_o21ai_1 _13174_ (.B1(_07754_),
    .Y(_07755_),
    .A1(net4769),
    .A2(net2564));
 sg13g2_nand2_1 _13175_ (.Y(_07756_),
    .A(net5088),
    .B(net3701));
 sg13g2_o21ai_1 _13176_ (.B1(_07756_),
    .Y(_00604_),
    .A1(net3701),
    .A2(_07755_));
 sg13g2_nand2b_1 _13177_ (.Y(_07757_),
    .B(net4771),
    .A_N(net287));
 sg13g2_o21ai_1 _13178_ (.B1(_07757_),
    .Y(_07758_),
    .A1(net4769),
    .A2(net2565));
 sg13g2_nand2_1 _13179_ (.Y(_07759_),
    .A(net5085),
    .B(net3701));
 sg13g2_o21ai_1 _13180_ (.B1(_07759_),
    .Y(_00605_),
    .A1(net3701),
    .A2(_07758_));
 sg13g2_mux2_1 _13181_ (.A0(net2666),
    .A1(net255),
    .S(net4767),
    .X(_07760_));
 sg13g2_nor2_1 _13182_ (.A(net3699),
    .B(_07760_),
    .Y(_07761_));
 sg13g2_a21oi_1 _13183_ (.A1(_05648_),
    .A2(net3699),
    .Y(_00606_),
    .B1(_07761_));
 sg13g2_nand2b_1 _13184_ (.Y(_07762_),
    .B(net4765),
    .A_N(\soc_inst.mem_ctrl.next_instr_data[16] ));
 sg13g2_o21ai_1 _13185_ (.B1(_07762_),
    .Y(_07763_),
    .A1(net4763),
    .A2(\soc_inst.mem_ctrl.spi_data_out[8] ));
 sg13g2_nand2_1 _13186_ (.Y(_07764_),
    .A(net198),
    .B(net3696));
 sg13g2_o21ai_1 _13187_ (.B1(_07764_),
    .Y(_00607_),
    .A1(net3696),
    .A2(_07763_));
 sg13g2_nand2b_1 _13188_ (.Y(_07765_),
    .B(net4764),
    .A_N(net161));
 sg13g2_o21ai_1 _13189_ (.B1(_07765_),
    .Y(_07766_),
    .A1(net4764),
    .A2(\soc_inst.mem_ctrl.spi_data_out[9] ));
 sg13g2_nand2_1 _13190_ (.Y(_07767_),
    .A(net391),
    .B(net3695));
 sg13g2_o21ai_1 _13191_ (.B1(_07767_),
    .Y(_00608_),
    .A1(net3695),
    .A2(_07766_));
 sg13g2_nand2b_1 _13192_ (.Y(_07768_),
    .B(net4765),
    .A_N(net115));
 sg13g2_o21ai_1 _13193_ (.B1(_07768_),
    .Y(_07769_),
    .A1(net4765),
    .A2(\soc_inst.mem_ctrl.spi_data_out[10] ));
 sg13g2_nand2_1 _13194_ (.Y(_07770_),
    .A(net362),
    .B(net3696));
 sg13g2_o21ai_1 _13195_ (.B1(_07770_),
    .Y(_00609_),
    .A1(net3697),
    .A2(_07769_));
 sg13g2_nand2b_1 _13196_ (.Y(_07771_),
    .B(net4765),
    .A_N(net126));
 sg13g2_o21ai_1 _13197_ (.B1(_07771_),
    .Y(_07772_),
    .A1(net4765),
    .A2(\soc_inst.mem_ctrl.spi_data_out[11] ));
 sg13g2_nand2_1 _13198_ (.Y(_07773_),
    .A(net395),
    .B(net3696));
 sg13g2_o21ai_1 _13199_ (.B1(_07773_),
    .Y(_00610_),
    .A1(net3696),
    .A2(_07772_));
 sg13g2_nand2b_1 _13200_ (.Y(_07774_),
    .B(net4763),
    .A_N(net262));
 sg13g2_o21ai_1 _13201_ (.B1(_07774_),
    .Y(_07775_),
    .A1(net4764),
    .A2(\soc_inst.mem_ctrl.spi_data_out[12] ));
 sg13g2_nand2_1 _13202_ (.Y(_07776_),
    .A(net370),
    .B(net3695));
 sg13g2_o21ai_1 _13203_ (.B1(_07776_),
    .Y(_00611_),
    .A1(net3697),
    .A2(_07775_));
 sg13g2_nand2b_1 _13204_ (.Y(_07777_),
    .B(net4766),
    .A_N(net122));
 sg13g2_o21ai_1 _13205_ (.B1(_07777_),
    .Y(_07778_),
    .A1(net4764),
    .A2(\soc_inst.mem_ctrl.spi_data_out[13] ));
 sg13g2_nand2_1 _13206_ (.Y(_07779_),
    .A(net309),
    .B(net3694));
 sg13g2_o21ai_1 _13207_ (.B1(_07779_),
    .Y(_00612_),
    .A1(net3694),
    .A2(_07778_));
 sg13g2_mux2_1 _13208_ (.A0(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .A1(net251),
    .S(net4763),
    .X(_07780_));
 sg13g2_nor2_1 _13209_ (.A(net3694),
    .B(_07780_),
    .Y(_07781_));
 sg13g2_a21oi_1 _13210_ (.A1(_05733_),
    .A2(net3694),
    .Y(_00613_),
    .B1(_07781_));
 sg13g2_nand2b_1 _13211_ (.Y(_07782_),
    .B(net4763),
    .A_N(net184));
 sg13g2_o21ai_1 _13212_ (.B1(_07782_),
    .Y(_07783_),
    .A1(net4764),
    .A2(\soc_inst.mem_ctrl.spi_data_out[15] ));
 sg13g2_nand2_1 _13213_ (.Y(_07784_),
    .A(net191),
    .B(net3694));
 sg13g2_o21ai_1 _13214_ (.B1(_07784_),
    .Y(_00614_),
    .A1(net3694),
    .A2(_07783_));
 sg13g2_nand2b_1 _13215_ (.Y(_07785_),
    .B(net4765),
    .A_N(net146));
 sg13g2_o21ai_1 _13216_ (.B1(_07785_),
    .Y(_07786_),
    .A1(net4765),
    .A2(\soc_inst.mem_ctrl.spi_data_out[0] ));
 sg13g2_nand2_1 _13217_ (.Y(_07787_),
    .A(net266),
    .B(net3696));
 sg13g2_o21ai_1 _13218_ (.B1(_07787_),
    .Y(_00615_),
    .A1(net3696),
    .A2(_07786_));
 sg13g2_nand2_1 _13219_ (.Y(_07788_),
    .A(net4770),
    .B(net298));
 sg13g2_o21ai_1 _13220_ (.B1(_07788_),
    .Y(_07789_),
    .A1(net4770),
    .A2(_05585_));
 sg13g2_mux2_1 _13221_ (.A0(_07789_),
    .A1(net2096),
    .S(net3703),
    .X(_00616_));
 sg13g2_nand2b_1 _13222_ (.Y(_07790_),
    .B(net4767),
    .A_N(net230));
 sg13g2_o21ai_1 _13223_ (.B1(_07790_),
    .Y(_07791_),
    .A1(net4765),
    .A2(\soc_inst.mem_ctrl.spi_data_out[2] ));
 sg13g2_nand2_1 _13224_ (.Y(_07792_),
    .A(net275),
    .B(net3697));
 sg13g2_o21ai_1 _13225_ (.B1(_07792_),
    .Y(_00617_),
    .A1(net3696),
    .A2(_07791_));
 sg13g2_nand2_1 _13226_ (.Y(_07793_),
    .A(net4770),
    .B(net222));
 sg13g2_o21ai_1 _13227_ (.B1(_07793_),
    .Y(_07794_),
    .A1(net4770),
    .A2(_05586_));
 sg13g2_mux2_1 _13228_ (.A0(_07794_),
    .A1(net1441),
    .S(net3703),
    .X(_00618_));
 sg13g2_nand2b_1 _13229_ (.Y(_07795_),
    .B(net4763),
    .A_N(net247));
 sg13g2_o21ai_1 _13230_ (.B1(_07795_),
    .Y(_07796_),
    .A1(net4763),
    .A2(\soc_inst.mem_ctrl.spi_data_out[4] ));
 sg13g2_nand2_1 _13231_ (.Y(_07797_),
    .A(net452),
    .B(net3695));
 sg13g2_o21ai_1 _13232_ (.B1(_07797_),
    .Y(_00619_),
    .A1(net3695),
    .A2(_07796_));
 sg13g2_nand2_1 _13233_ (.Y(_07798_),
    .A(net4770),
    .B(net253));
 sg13g2_o21ai_1 _13234_ (.B1(_07798_),
    .Y(_07799_),
    .A1(net4770),
    .A2(_05587_));
 sg13g2_mux2_1 _13235_ (.A0(_07799_),
    .A1(net1136),
    .S(net3702),
    .X(_00620_));
 sg13g2_nand2b_1 _13236_ (.Y(_07800_),
    .B(net4764),
    .A_N(net189));
 sg13g2_o21ai_1 _13237_ (.B1(_07800_),
    .Y(_07801_),
    .A1(net4764),
    .A2(\soc_inst.mem_ctrl.spi_data_out[6] ));
 sg13g2_nand2_1 _13238_ (.Y(_07802_),
    .A(net321),
    .B(net3694));
 sg13g2_o21ai_1 _13239_ (.B1(_07802_),
    .Y(_00621_),
    .A1(net3694),
    .A2(_07801_));
 sg13g2_nand2b_1 _13240_ (.Y(_07803_),
    .B(net4763),
    .A_N(net249));
 sg13g2_o21ai_1 _13241_ (.B1(_07803_),
    .Y(_07804_),
    .A1(net4763),
    .A2(\soc_inst.mem_ctrl.spi_data_out[7] ));
 sg13g2_nand2_1 _13242_ (.Y(_07805_),
    .A(net319),
    .B(net3695));
 sg13g2_o21ai_1 _13243_ (.B1(_07805_),
    .Y(_00622_),
    .A1(net3695),
    .A2(_07804_));
 sg13g2_nor2_1 _13244_ (.A(_05871_),
    .B(_06018_),
    .Y(_07806_));
 sg13g2_o21ai_1 _13245_ (.B1(_06030_),
    .Y(_07807_),
    .A1(net4015),
    .A2(_07806_));
 sg13g2_nand2_1 _13246_ (.Y(_07808_),
    .A(_05417_),
    .B(\soc_inst.mem_ctrl.access_state[3] ));
 sg13g2_a21oi_1 _13247_ (.A1(_05906_),
    .A2(_07808_),
    .Y(_07809_),
    .B1(_07807_));
 sg13g2_a21o_2 _13248_ (.A2(_07808_),
    .A1(_05906_),
    .B1(_07807_),
    .X(_07810_));
 sg13g2_a21oi_1 _13249_ (.A1(net4757),
    .A2(net4868),
    .Y(_07811_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[24] ));
 sg13g2_a21oi_1 _13250_ (.A1(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .A2(net4704),
    .Y(_07812_),
    .B1(_06676_));
 sg13g2_o21ai_1 _13251_ (.B1(_07812_),
    .Y(_07813_),
    .A1(net4704),
    .A2(_07811_));
 sg13g2_o21ai_1 _13252_ (.B1(_07813_),
    .Y(_07814_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .A2(net4711));
 sg13g2_a22oi_1 _13253_ (.Y(_07815_),
    .B1(net4261),
    .B2(\soc_inst.gpio_inst.int_pend_reg[0] ),
    .A2(net4206),
    .A1(\soc_inst.gpio_inst.int_en_reg[0] ));
 sg13g2_nand2_1 _13254_ (.Y(_07816_),
    .A(\soc_inst.gpio_bidir_out [0]),
    .B(net4260));
 sg13g2_nand2_1 _13255_ (.Y(_07817_),
    .A(net13),
    .B(net4179));
 sg13g2_nand4_1 _13256_ (.B(_07815_),
    .C(_07816_),
    .A(_07120_),
    .Y(_07818_),
    .D(_07817_));
 sg13g2_o21ai_1 _13257_ (.B1(_07818_),
    .Y(_07819_),
    .A1(\soc_inst.gpio_bidir_oe [0]),
    .A2(_07120_));
 sg13g2_and2_1 _13258_ (.A(net4800),
    .B(_05897_),
    .X(_07820_));
 sg13g2_nand2_1 _13259_ (.Y(_07821_),
    .A(net4801),
    .B(_05897_));
 sg13g2_nor2_1 _13260_ (.A(_07819_),
    .B(_07821_),
    .Y(_07822_));
 sg13g2_nor2_2 _13261_ (.A(net4651),
    .B(_06523_),
    .Y(_07823_));
 sg13g2_or2_1 _13262_ (.X(_07824_),
    .B(_06523_),
    .A(net4651));
 sg13g2_or2_1 _13263_ (.X(_07825_),
    .B(\soc_inst.spi_inst.len_sel[0] ),
    .A(net5125));
 sg13g2_a22oi_1 _13264_ (.Y(_07826_),
    .B1(_06939_),
    .B2(_05544_),
    .A2(net5125),
    .A1(_05545_));
 sg13g2_o21ai_1 _13265_ (.B1(_07826_),
    .Y(_07827_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .A2(net4697));
 sg13g2_o21ai_1 _13266_ (.B1(_07120_),
    .Y(_07828_),
    .A1(_07824_),
    .A2(_07827_));
 sg13g2_a221oi_1 _13267_ (.B2(\soc_inst.spi_inst.busy ),
    .C1(_07828_),
    .B1(net4178),
    .A1(_05409_),
    .Y(_07829_),
    .A2(net4261));
 sg13g2_nor2_1 _13268_ (.A(\soc_inst.spi_ena ),
    .B(_07120_),
    .Y(_07830_));
 sg13g2_nor2_1 _13269_ (.A(_00295_),
    .B(net4269),
    .Y(_07831_));
 sg13g2_nor2_1 _13270_ (.A(_00277_),
    .B(net4654),
    .Y(_07832_));
 sg13g2_nor3_1 _13271_ (.A(net4715),
    .B(_07831_),
    .C(_07832_),
    .Y(_07833_));
 sg13g2_a221oi_1 _13272_ (.B2(_05516_),
    .C1(_07833_),
    .B1(net4264),
    .A1(_00169_),
    .Y(_07834_),
    .A2(_06411_));
 sg13g2_nand3_1 _13273_ (.B(_05423_),
    .C(_05883_),
    .A(net4801),
    .Y(_07835_));
 sg13g2_nand2_1 _13274_ (.Y(_07836_),
    .A(net4793),
    .B(\soc_inst.pwm_inst.channel_counter[1][0] ));
 sg13g2_o21ai_1 _13275_ (.B1(_07836_),
    .Y(_07837_),
    .A1(net4793),
    .A2(_05582_));
 sg13g2_mux2_1 _13276_ (.A0(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .A1(\soc_inst.pwm_inst.channel_duty[1][0] ),
    .S(net4794),
    .X(_07838_));
 sg13g2_nor2_1 _13277_ (.A(_00230_),
    .B(net4793),
    .Y(_07839_));
 sg13g2_o21ai_1 _13278_ (.B1(net4797),
    .Y(_07840_),
    .A1(_00246_),
    .A2(net4738));
 sg13g2_o21ai_1 _13279_ (.B1(net4714),
    .Y(_07841_),
    .A1(_07839_),
    .A2(_07840_));
 sg13g2_a22oi_1 _13280_ (.Y(_07842_),
    .B1(_07838_),
    .B2(net4273),
    .A2(_07837_),
    .A1(net4277));
 sg13g2_nand2_1 _13281_ (.Y(_07843_),
    .A(net4789),
    .B(\soc_inst.pwm_ena[1] ));
 sg13g2_a21oi_1 _13282_ (.A1(net4740),
    .A2(\soc_inst.pwm_ena[0] ),
    .Y(_07844_),
    .B1(net4652));
 sg13g2_a22oi_1 _13283_ (.Y(_07845_),
    .B1(_07843_),
    .B2(_07844_),
    .A2(_07842_),
    .A1(_07841_));
 sg13g2_nand4_1 _13284_ (.B(net4787),
    .C(_05883_),
    .A(net4801),
    .Y(_07846_),
    .D(_06287_));
 sg13g2_and4_1 _13285_ (.A(net4800),
    .B(net4787),
    .C(_05896_),
    .D(_06287_),
    .X(_07847_));
 sg13g2_a21oi_1 _13286_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ),
    .A2(net4206),
    .Y(_07848_),
    .B1(net4259));
 sg13g2_a22oi_1 _13287_ (.Y(_07849_),
    .B1(_07823_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .A2(net4178),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ));
 sg13g2_nor2_2 _13288_ (.A(net2738),
    .B(net2809),
    .Y(_07850_));
 sg13g2_a21oi_1 _13289_ (.A1(_00222_),
    .A2(net4795),
    .Y(_07851_),
    .B1(net4655));
 sg13g2_a21o_1 _13290_ (.A2(net4272),
    .A1(\soc_inst.i2c_inst.data_reg[0] ),
    .B1(_07851_),
    .X(_07852_));
 sg13g2_o21ai_1 _13291_ (.B1(_07852_),
    .Y(_07853_),
    .A1(\soc_inst.i2c_inst.status_reg[0] ),
    .A2(net4643));
 sg13g2_nand2_2 _13292_ (.Y(_07854_),
    .A(net4800),
    .B(_05899_));
 sg13g2_nor3_1 _13293_ (.A(_07829_),
    .B(_07830_),
    .C(_07854_),
    .Y(_07855_));
 sg13g2_nand2_2 _13294_ (.Y(_07856_),
    .A(net4800),
    .B(_05901_));
 sg13g2_a221oi_1 _13295_ (.B2(net4259),
    .C1(_07856_),
    .B1(_07850_),
    .A1(_07848_),
    .Y(_07857_),
    .A2(_07849_));
 sg13g2_nor3_1 _13296_ (.A(_07822_),
    .B(_07855_),
    .C(_07857_),
    .Y(_07858_));
 sg13g2_nand2_2 _13297_ (.Y(_07859_),
    .A(net4800),
    .B(_05902_));
 sg13g2_o21ai_1 _13298_ (.B1(net4018),
    .Y(_07860_),
    .A1(_07853_),
    .A2(_07859_));
 sg13g2_nor3_2 _13299_ (.A(net4787),
    .B(_05876_),
    .C(_05895_),
    .Y(_07861_));
 sg13g2_and2_1 _13300_ (.A(net4800),
    .B(_07861_),
    .X(_07862_));
 sg13g2_a221oi_1 _13301_ (.B2(_07834_),
    .C1(_07860_),
    .B1(_07862_),
    .A1(_07845_),
    .Y(_07863_),
    .A2(net4044));
 sg13g2_a22oi_1 _13302_ (.Y(_07864_),
    .B1(_07858_),
    .B2(_07863_),
    .A2(_07814_),
    .A1(_05905_));
 sg13g2_mux2_1 _13303_ (.A0(net2502),
    .A1(_07864_),
    .S(net3815),
    .X(_00623_));
 sg13g2_o21ai_1 _13304_ (.B1(net4652),
    .Y(_07865_),
    .A1(_00296_),
    .A2(net4269));
 sg13g2_a221oi_1 _13305_ (.B2(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .C1(_07865_),
    .B1(net4264),
    .A1(_05402_),
    .Y(_07866_),
    .A2(_06295_));
 sg13g2_nand2_1 _13306_ (.Y(_07867_),
    .A(_00223_),
    .B(net4795));
 sg13g2_a22oi_1 _13307_ (.Y(_07868_),
    .B1(_07867_),
    .B2(net4657),
    .A2(net4272),
    .A1(\soc_inst.i2c_inst.data_reg[1] ));
 sg13g2_nor2_1 _13308_ (.A(\soc_inst.i2c_inst.status_reg[1] ),
    .B(net4644),
    .Y(_07869_));
 sg13g2_nand2_1 _13309_ (.Y(_07870_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .B(net4206));
 sg13g2_a22oi_1 _13310_ (.Y(_07871_),
    .B1(_07823_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .A2(net4178),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ));
 sg13g2_nand2b_1 _13311_ (.Y(_07872_),
    .B(net5125),
    .A_N(\soc_inst.spi_inst.rx_shift_reg[25] ));
 sg13g2_o21ai_1 _13312_ (.B1(_07872_),
    .Y(_07873_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .A2(net4702));
 sg13g2_nor2_1 _13313_ (.A(_07824_),
    .B(_07873_),
    .Y(_07874_));
 sg13g2_o21ai_1 _13314_ (.B1(_07874_),
    .Y(_07875_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .A2(_07825_));
 sg13g2_a21oi_1 _13315_ (.A1(\soc_inst.gpio_inst.int_en_reg[1] ),
    .A2(net4206),
    .Y(_07876_),
    .B1(net4260));
 sg13g2_a22oi_1 _13316_ (.Y(_07877_),
    .B1(net4179),
    .B2(net3),
    .A2(net4261),
    .A1(\soc_inst.gpio_inst.int_pend_reg[1] ));
 sg13g2_nand2b_1 _13317_ (.Y(_07878_),
    .B(net4704),
    .A_N(\soc_inst.mem_ctrl.spi_data_out[9] ));
 sg13g2_o21ai_1 _13318_ (.B1(_07878_),
    .Y(_07879_),
    .A1(net4757),
    .A2(\soc_inst.mem_ctrl.spi_data_out[25] ));
 sg13g2_a21oi_2 _13319_ (.B1(_07879_),
    .Y(_07880_),
    .A2(_06673_),
    .A1(_05585_));
 sg13g2_mux2_1 _13320_ (.A0(_05589_),
    .A1(_05590_),
    .S(net4794),
    .X(_07881_));
 sg13g2_a21oi_1 _13321_ (.A1(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .A2(net4277),
    .Y(_07882_),
    .B1(net4792));
 sg13g2_o21ai_1 _13322_ (.B1(_07882_),
    .Y(_07883_),
    .A1(_00231_),
    .A2(net4642));
 sg13g2_nor2_1 _13323_ (.A(_05574_),
    .B(_06296_),
    .Y(_07884_));
 sg13g2_o21ai_1 _13324_ (.B1(net4792),
    .Y(_07885_),
    .A1(_00247_),
    .A2(net4642));
 sg13g2_o21ai_1 _13325_ (.B1(_07883_),
    .Y(_07886_),
    .A1(_07884_),
    .A2(_07885_));
 sg13g2_o21ai_1 _13326_ (.B1(_07886_),
    .Y(_07887_),
    .A1(net4270),
    .A2(_07881_));
 sg13g2_a21oi_1 _13327_ (.A1(_05408_),
    .A2(net4261),
    .Y(_07888_),
    .B1(net4178));
 sg13g2_a221oi_1 _13328_ (.B2(_07877_),
    .C1(_07821_),
    .B1(_07876_),
    .A1(_05588_),
    .Y(_07889_),
    .A2(net4260));
 sg13g2_a21oi_2 _13329_ (.B1(_07856_),
    .Y(_07890_),
    .A2(_07871_),
    .A1(_07870_));
 sg13g2_a221oi_1 _13330_ (.B2(_07888_),
    .C1(_07854_),
    .B1(_07875_),
    .A1(_05591_),
    .Y(_07891_),
    .A2(net4178));
 sg13g2_o21ai_1 _13331_ (.B1(net4043),
    .Y(_07892_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .A2(net4651));
 sg13g2_nor3_1 _13332_ (.A(_07859_),
    .B(_07868_),
    .C(_07869_),
    .Y(_07893_));
 sg13g2_a21oi_1 _13333_ (.A1(net4044),
    .A2(_07887_),
    .Y(_07894_),
    .B1(_07893_));
 sg13g2_o21ai_1 _13334_ (.B1(_07894_),
    .Y(_07895_),
    .A1(_07866_),
    .A2(_07892_));
 sg13g2_nor4_2 _13335_ (.A(_07889_),
    .B(_07890_),
    .C(_07891_),
    .Y(_07896_),
    .D(_07895_));
 sg13g2_a21oi_1 _13336_ (.A1(_05905_),
    .A2(_07880_),
    .Y(_07897_),
    .B1(net3808));
 sg13g2_a22oi_1 _13337_ (.Y(_00624_),
    .B1(_07896_),
    .B2(_07897_),
    .A2(net3808),
    .A1(_05611_));
 sg13g2_nand2_1 _13338_ (.Y(_07898_),
    .A(net289),
    .B(net3809));
 sg13g2_a22oi_1 _13339_ (.Y(_07899_),
    .B1(net4704),
    .B2(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .A2(_06673_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[2] ));
 sg13g2_o21ai_1 _13340_ (.B1(_07899_),
    .Y(_07900_),
    .A1(net4757),
    .A2(_05583_));
 sg13g2_nand2_1 _13341_ (.Y(_07901_),
    .A(_00224_),
    .B(net4795));
 sg13g2_a22oi_1 _13342_ (.Y(_07902_),
    .B1(_07901_),
    .B2(net4657),
    .A2(net4272),
    .A1(\soc_inst.i2c_inst.data_reg[2] ));
 sg13g2_nor2_1 _13343_ (.A(\soc_inst.i2c_inst.status_reg[2] ),
    .B(net4644),
    .Y(_07903_));
 sg13g2_o21ai_1 _13344_ (.B1(net4651),
    .Y(_07904_),
    .A1(_07902_),
    .A2(_07903_));
 sg13g2_or2_1 _13345_ (.X(_07905_),
    .B(net4697),
    .A(\soc_inst.spi_inst.rx_shift_reg[2] ));
 sg13g2_o21ai_1 _13346_ (.B1(_07905_),
    .Y(_07906_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .A2(net4702));
 sg13g2_a21oi_1 _13347_ (.A1(_05546_),
    .A2(net5126),
    .Y(_07907_),
    .B1(_07906_));
 sg13g2_and3_1 _13348_ (.X(_07908_),
    .A(net4800),
    .B(_06299_),
    .C(_07823_));
 sg13g2_a21oi_1 _13349_ (.A1(net4),
    .A2(net4179),
    .Y(_07909_),
    .B1(net4260));
 sg13g2_a22oi_1 _13350_ (.Y(_07910_),
    .B1(net4261),
    .B2(\soc_inst.gpio_inst.int_pend_reg[2] ),
    .A2(net4206),
    .A1(\soc_inst.gpio_inst.int_en_reg[2] ));
 sg13g2_a221oi_1 _13351_ (.B2(_05396_),
    .C1(net4714),
    .B1(net4273),
    .A1(_05401_),
    .Y(_07911_),
    .A2(_06295_));
 sg13g2_a221oi_1 _13352_ (.B2(_05515_),
    .C1(_07911_),
    .B1(net4264),
    .A1(_05508_),
    .Y(_07912_),
    .A2(_06411_));
 sg13g2_nor2_1 _13353_ (.A(_00327_),
    .B(_07824_),
    .Y(_07913_));
 sg13g2_mux2_1 _13354_ (.A0(_00232_),
    .A1(_00248_),
    .S(net4792),
    .X(_07914_));
 sg13g2_nor2_1 _13355_ (.A(net4792),
    .B(\soc_inst.pwm_inst.channel_duty[0][2] ),
    .Y(_07915_));
 sg13g2_a21oi_1 _13356_ (.A1(net4793),
    .A2(_05593_),
    .Y(_07916_),
    .B1(_07915_));
 sg13g2_nor2_1 _13357_ (.A(net4792),
    .B(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .Y(_07917_));
 sg13g2_a21oi_1 _13358_ (.A1(net4792),
    .A2(_05573_),
    .Y(_07918_),
    .B1(_07917_));
 sg13g2_a221oi_1 _13359_ (.B2(net4277),
    .C1(net4264),
    .B1(_07918_),
    .A1(net4271),
    .Y(_07919_),
    .A2(_07916_));
 sg13g2_a21oi_1 _13360_ (.A1(_06521_),
    .A2(_07914_),
    .Y(_07920_),
    .B1(_07919_));
 sg13g2_o21ai_1 _13361_ (.B1(_07904_),
    .Y(_07921_),
    .A1(net5128),
    .A2(net4651));
 sg13g2_nor2_1 _13362_ (.A(_07859_),
    .B(_07921_),
    .Y(_07922_));
 sg13g2_o21ai_1 _13363_ (.B1(_07820_),
    .Y(_07923_),
    .A1(\soc_inst.gpio_inst.gpio_out[1] ),
    .A2(_06592_));
 sg13g2_a21oi_2 _13364_ (.B1(_07923_),
    .Y(_07924_),
    .A2(_07910_),
    .A1(_07909_));
 sg13g2_a221oi_1 _13365_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ),
    .C1(_07913_),
    .B1(net4178),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_rx_break_reg ),
    .Y(_07925_),
    .A2(net4206));
 sg13g2_nor2_1 _13366_ (.A(_07856_),
    .B(_07925_),
    .Y(_07926_));
 sg13g2_nor3_1 _13367_ (.A(_07922_),
    .B(_07924_),
    .C(_07926_),
    .Y(_07927_));
 sg13g2_a22oi_1 _13368_ (.Y(_07928_),
    .B1(_07920_),
    .B2(net4044),
    .A2(_07912_),
    .A1(net4043));
 sg13g2_nor2_2 _13369_ (.A(_07824_),
    .B(_07854_),
    .Y(_07929_));
 sg13g2_nor2_2 _13370_ (.A(_06525_),
    .B(_07854_),
    .Y(_07930_));
 sg13g2_a22oi_1 _13371_ (.Y(_07931_),
    .B1(_07930_),
    .B2(_05407_),
    .A2(net3978),
    .A1(_07907_));
 sg13g2_nand4_1 _13372_ (.B(_07927_),
    .C(_07928_),
    .A(net4018),
    .Y(_07932_),
    .D(_07931_));
 sg13g2_o21ai_1 _13373_ (.B1(_07932_),
    .Y(_07933_),
    .A1(net4016),
    .A2(_07900_));
 sg13g2_o21ai_1 _13374_ (.B1(_07898_),
    .Y(_00625_),
    .A1(net3809),
    .A2(_07933_));
 sg13g2_nand2_1 _13375_ (.Y(_07934_),
    .A(net294),
    .B(net3809));
 sg13g2_a22oi_1 _13376_ (.Y(_07935_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .B2(net4704),
    .A2(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .A1(net4873));
 sg13g2_o21ai_1 _13377_ (.B1(_07935_),
    .Y(_07936_),
    .A1(_05586_),
    .A2(net4711));
 sg13g2_o21ai_1 _13378_ (.B1(net3816),
    .Y(_07937_),
    .A1(net4015),
    .A2(_07936_));
 sg13g2_a21oi_1 _13379_ (.A1(_05400_),
    .A2(net4657),
    .Y(_07938_),
    .B1(net4714));
 sg13g2_o21ai_1 _13380_ (.B1(_07938_),
    .Y(_07939_),
    .A1(_00298_),
    .A2(net4269));
 sg13g2_o21ai_1 _13381_ (.B1(_07939_),
    .Y(_07940_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .A2(net4643));
 sg13g2_a21oi_1 _13382_ (.A1(_05507_),
    .A2(_06411_),
    .Y(_07941_),
    .B1(_07940_));
 sg13g2_a22oi_1 _13383_ (.Y(_07942_),
    .B1(net4261),
    .B2(\soc_inst.gpio_inst.int_pend_reg[3] ),
    .A2(net4207),
    .A1(\soc_inst.gpio_inst.int_en_reg[3] ));
 sg13g2_a21oi_1 _13384_ (.A1(net5),
    .A2(net4179),
    .Y(_07943_),
    .B1(net4260));
 sg13g2_or2_1 _13385_ (.X(_07944_),
    .B(net4792),
    .A(_00233_));
 sg13g2_o21ai_1 _13386_ (.B1(_07944_),
    .Y(_07945_),
    .A1(_00249_),
    .A2(net4738));
 sg13g2_a221oi_1 _13387_ (.B2(\soc_inst.pwm_inst.channel_duty[1][3] ),
    .C1(net4738),
    .B1(net4271),
    .A1(\soc_inst.pwm_inst.channel_counter[1][3] ),
    .Y(_07946_),
    .A2(net4277));
 sg13g2_a221oi_1 _13388_ (.B2(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .C1(net4792),
    .B1(net4271),
    .A1(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .Y(_07947_),
    .A2(net4277));
 sg13g2_nor3_1 _13389_ (.A(net4262),
    .B(_07946_),
    .C(_07947_),
    .Y(_07948_));
 sg13g2_a21o_1 _13390_ (.A2(_07945_),
    .A1(net4264),
    .B1(_07948_),
    .X(_07949_));
 sg13g2_nand2_1 _13391_ (.Y(_07950_),
    .A(_00225_),
    .B(net4796));
 sg13g2_a22oi_1 _13392_ (.Y(_07951_),
    .B1(_07950_),
    .B2(net4657),
    .A2(net4273),
    .A1(\soc_inst.i2c_inst.data_reg[3] ));
 sg13g2_nor2_1 _13393_ (.A(\soc_inst.i2c_inst.status_reg[3] ),
    .B(net4644),
    .Y(_07952_));
 sg13g2_o21ai_1 _13394_ (.B1(net4652),
    .Y(_07953_),
    .A1(_07951_),
    .A2(_07952_));
 sg13g2_or2_1 _13395_ (.X(_07954_),
    .B(net4697),
    .A(\soc_inst.spi_inst.rx_shift_reg[3] ));
 sg13g2_o21ai_1 _13396_ (.B1(_07954_),
    .Y(_07955_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .A2(net4701));
 sg13g2_a21oi_1 _13397_ (.A1(_05547_),
    .A2(net5125),
    .Y(_07956_),
    .B1(_07955_));
 sg13g2_o21ai_1 _13398_ (.B1(_07953_),
    .Y(_07957_),
    .A1(\soc_inst.i2c_inst.ack_enable ),
    .A2(net4652));
 sg13g2_a22oi_1 _13399_ (.Y(_07958_),
    .B1(_07949_),
    .B2(net4044),
    .A2(_07941_),
    .A1(net4043));
 sg13g2_o21ai_1 _13400_ (.B1(_07958_),
    .Y(_07959_),
    .A1(_07859_),
    .A2(_07957_));
 sg13g2_o21ai_1 _13401_ (.B1(_07820_),
    .Y(_07960_),
    .A1(\soc_inst.gpio_inst.gpio_out[2] ),
    .A2(_06592_));
 sg13g2_a21oi_1 _13402_ (.A1(_07942_),
    .A2(_07943_),
    .Y(_07961_),
    .B1(_07960_));
 sg13g2_nor3_2 _13403_ (.A(_06289_),
    .B(net4269),
    .C(_07856_),
    .Y(_07962_));
 sg13g2_a22oi_1 _13404_ (.Y(_07963_),
    .B1(_07962_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ),
    .A2(_07930_),
    .A1(_05406_));
 sg13g2_nor2_2 _13405_ (.A(_07824_),
    .B(_07856_),
    .Y(_07964_));
 sg13g2_a22oi_1 _13406_ (.Y(_07965_),
    .B1(_07964_),
    .B2(_05389_),
    .A2(_07956_),
    .A1(net3978));
 sg13g2_nand2_1 _13407_ (.Y(_07966_),
    .A(_07963_),
    .B(_07965_));
 sg13g2_nor4_2 _13408_ (.A(_05905_),
    .B(_07959_),
    .C(_07961_),
    .Y(_07967_),
    .D(_07966_));
 sg13g2_o21ai_1 _13409_ (.B1(_07934_),
    .Y(_00626_),
    .A1(_07937_),
    .A2(_07967_));
 sg13g2_and2_1 _13410_ (.A(net4873),
    .B(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .X(_07968_));
 sg13g2_a221oi_1 _13411_ (.B2(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .C1(_07968_),
    .B1(net4704),
    .A1(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .Y(_07969_),
    .A2(_06673_));
 sg13g2_or2_1 _13412_ (.X(_07970_),
    .B(net4697),
    .A(\soc_inst.spi_inst.rx_shift_reg[4] ));
 sg13g2_o21ai_1 _13413_ (.B1(_07970_),
    .Y(_07971_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .A2(net4701));
 sg13g2_a21oi_1 _13414_ (.A1(_05548_),
    .A2(\soc_inst.spi_inst.len_sel[1] ),
    .Y(_07972_),
    .B1(_07971_));
 sg13g2_a22oi_1 _13415_ (.Y(_07973_),
    .B1(net4261),
    .B2(\soc_inst.gpio_inst.int_pend_reg[4] ),
    .A2(net4207),
    .A1(\soc_inst.gpio_inst.int_en_reg[4] ));
 sg13g2_a21oi_1 _13416_ (.A1(net6),
    .A2(net4179),
    .Y(_07974_),
    .B1(net4260));
 sg13g2_a22oi_1 _13417_ (.Y(_07975_),
    .B1(net4272),
    .B2(\soc_inst.pwm_inst.channel_duty[0][4] ),
    .A2(net4656),
    .A1(\soc_inst.pwm_inst.channel_counter[0][4] ));
 sg13g2_or2_1 _13418_ (.X(_07976_),
    .B(_07975_),
    .A(net4790));
 sg13g2_nand2_1 _13419_ (.Y(_07977_),
    .A(\soc_inst.pwm_inst.channel_counter[1][4] ),
    .B(net4656));
 sg13g2_o21ai_1 _13420_ (.B1(_07977_),
    .Y(_07978_),
    .A1(_05595_),
    .A2(net4270));
 sg13g2_a21oi_1 _13421_ (.A1(net4790),
    .A2(_07978_),
    .Y(_07979_),
    .B1(net4262));
 sg13g2_mux2_1 _13422_ (.A0(_00234_),
    .A1(_00250_),
    .S(net4790),
    .X(_07980_));
 sg13g2_nor2_1 _13423_ (.A(_00226_),
    .B(_06296_),
    .Y(_07981_));
 sg13g2_a221oi_1 _13424_ (.B2(\soc_inst.i2c_inst.data_reg[4] ),
    .C1(_07981_),
    .B1(net4273),
    .A1(\soc_inst.i2c_inst.ctrl_reg[4] ),
    .Y(_07982_),
    .A2(_06411_));
 sg13g2_nor2_1 _13425_ (.A(_00299_),
    .B(net4269),
    .Y(_07983_));
 sg13g2_nor2_1 _13426_ (.A(_00281_),
    .B(net4655),
    .Y(_07984_));
 sg13g2_nor3_1 _13427_ (.A(net4714),
    .B(_07983_),
    .C(_07984_),
    .Y(_07985_));
 sg13g2_nor2_1 _13428_ (.A(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .B(net4643),
    .Y(_07986_));
 sg13g2_nor2_1 _13429_ (.A(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .B(net4651),
    .Y(_07987_));
 sg13g2_nor3_1 _13430_ (.A(_07985_),
    .B(_07986_),
    .C(_07987_),
    .Y(_07988_));
 sg13g2_a22oi_1 _13431_ (.Y(_07989_),
    .B1(_07980_),
    .B2(net4262),
    .A2(_07979_),
    .A1(_07976_));
 sg13g2_nor3_1 _13432_ (.A(_00221_),
    .B(_06525_),
    .C(_07854_),
    .Y(_07990_));
 sg13g2_a221oi_1 _13433_ (.B2(net4044),
    .C1(_07990_),
    .B1(_07989_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .Y(_07991_),
    .A2(_07964_));
 sg13g2_a22oi_1 _13434_ (.Y(_07992_),
    .B1(_07973_),
    .B2(_07974_),
    .A2(net4260),
    .A1(_05594_));
 sg13g2_nor2_1 _13435_ (.A(_07859_),
    .B(_07982_),
    .Y(_07993_));
 sg13g2_a21oi_1 _13436_ (.A1(net3978),
    .A2(_07972_),
    .Y(_07994_),
    .B1(_07993_));
 sg13g2_a22oi_1 _13437_ (.Y(_07995_),
    .B1(_07988_),
    .B2(net4043),
    .A2(_07962_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ));
 sg13g2_nand3_1 _13438_ (.B(_07994_),
    .C(_07995_),
    .A(net4018),
    .Y(_07996_));
 sg13g2_a21oi_2 _13439_ (.B1(_07996_),
    .Y(_07997_),
    .A2(_07992_),
    .A1(_07820_));
 sg13g2_a221oi_1 _13440_ (.B2(_07997_),
    .C1(net3808),
    .B1(_07991_),
    .A1(_05905_),
    .Y(_07998_),
    .A2(_07969_));
 sg13g2_a21o_1 _13441_ (.A2(net3808),
    .A1(net1884),
    .B1(_07998_),
    .X(_00627_));
 sg13g2_nand2_1 _13442_ (.Y(_07999_),
    .A(net300),
    .B(net3809));
 sg13g2_nand2b_1 _13443_ (.Y(_08000_),
    .B(net4704),
    .A_N(\soc_inst.mem_ctrl.spi_data_out[13] ));
 sg13g2_o21ai_1 _13444_ (.B1(_08000_),
    .Y(_08001_),
    .A1(net4757),
    .A2(\soc_inst.mem_ctrl.spi_data_out[29] ));
 sg13g2_a21oi_1 _13445_ (.A1(_05587_),
    .A2(_06673_),
    .Y(_08002_),
    .B1(_08001_));
 sg13g2_nor2_1 _13446_ (.A(_00300_),
    .B(net4269),
    .Y(_08003_));
 sg13g2_nor2_1 _13447_ (.A(_00282_),
    .B(net4655),
    .Y(_08004_));
 sg13g2_nor3_1 _13448_ (.A(net4714),
    .B(_08003_),
    .C(_08004_),
    .Y(_08005_));
 sg13g2_nor2_1 _13449_ (.A(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .B(net4651),
    .Y(_08006_));
 sg13g2_nor2_1 _13450_ (.A(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .B(net4643),
    .Y(_08007_));
 sg13g2_nor3_1 _13451_ (.A(_08005_),
    .B(_08006_),
    .C(_08007_),
    .Y(_08008_));
 sg13g2_mux2_1 _13452_ (.A0(\soc_inst.i2c_inst.data_reg[5] ),
    .A1(\soc_inst.i2c_inst.prescale_reg[5] ),
    .S(net4798),
    .X(_08009_));
 sg13g2_or2_1 _13453_ (.X(_08010_),
    .B(net4697),
    .A(\soc_inst.spi_inst.rx_shift_reg[5] ));
 sg13g2_o21ai_1 _13454_ (.B1(_08010_),
    .Y(_08011_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .A2(net4701));
 sg13g2_a21oi_1 _13455_ (.A1(_05549_),
    .A2(\soc_inst.spi_inst.len_sel[1] ),
    .Y(_08012_),
    .B1(_08011_));
 sg13g2_nor2_1 _13456_ (.A(net4790),
    .B(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .Y(_08013_));
 sg13g2_a21oi_1 _13457_ (.A1(net4790),
    .A2(_05597_),
    .Y(_08014_),
    .B1(_08013_));
 sg13g2_mux2_1 _13458_ (.A0(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .A1(\soc_inst.pwm_inst.channel_counter[1][5] ),
    .S(net4791),
    .X(_08015_));
 sg13g2_a221oi_1 _13459_ (.B2(net4277),
    .C1(net4262),
    .B1(_08015_),
    .A1(net4271),
    .Y(_08016_),
    .A2(_08014_));
 sg13g2_mux2_1 _13460_ (.A0(_00235_),
    .A1(_00251_),
    .S(net4790),
    .X(_08017_));
 sg13g2_a21oi_2 _13461_ (.B1(_08016_),
    .Y(_08018_),
    .A2(_08017_),
    .A1(net4262));
 sg13g2_a21oi_1 _13462_ (.A1(net7),
    .A2(net4178),
    .Y(_08019_),
    .B1(net4259));
 sg13g2_a22oi_1 _13463_ (.Y(_08020_),
    .B1(net4261),
    .B2(\soc_inst.gpio_inst.int_pend_reg[5] ),
    .A2(net4207),
    .A1(\soc_inst.gpio_inst.int_en_reg[5] ));
 sg13g2_a22oi_1 _13464_ (.Y(_08021_),
    .B1(_07964_),
    .B2(_05388_),
    .A2(_07930_),
    .A1(\soc_inst.spi_inst.clock_divider[5] ));
 sg13g2_a22oi_1 _13465_ (.Y(_08022_),
    .B1(_08008_),
    .B2(net4043),
    .A2(_07962_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ));
 sg13g2_a22oi_1 _13466_ (.Y(_08023_),
    .B1(_08019_),
    .B2(_08020_),
    .A2(net4259),
    .A1(_05596_));
 sg13g2_a22oi_1 _13467_ (.Y(_08024_),
    .B1(_08018_),
    .B2(net4044),
    .A2(_08012_),
    .A1(net3978));
 sg13g2_nand4_1 _13468_ (.B(_05902_),
    .C(_06293_),
    .A(net4800),
    .Y(_08025_),
    .D(_08009_));
 sg13g2_nand3_1 _13469_ (.B(_08024_),
    .C(_08025_),
    .A(net4018),
    .Y(_08026_));
 sg13g2_a21oi_1 _13470_ (.A1(_07820_),
    .A2(_08023_),
    .Y(_08027_),
    .B1(_08026_));
 sg13g2_nand3_1 _13471_ (.B(_08022_),
    .C(_08027_),
    .A(_08021_),
    .Y(_08028_));
 sg13g2_o21ai_1 _13472_ (.B1(_08028_),
    .Y(_08029_),
    .A1(net4016),
    .A2(_08002_));
 sg13g2_o21ai_1 _13473_ (.B1(_07999_),
    .Y(_00628_),
    .A1(net3809),
    .A2(_08029_));
 sg13g2_and2_1 _13474_ (.A(net4873),
    .B(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .X(_08030_));
 sg13g2_a221oi_1 _13475_ (.B2(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .C1(_08030_),
    .B1(net4705),
    .A1(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .Y(_08031_),
    .A2(_06673_));
 sg13g2_a21oi_1 _13476_ (.A1(_05905_),
    .A2(_08031_),
    .Y(_08032_),
    .B1(_07810_));
 sg13g2_nor2_1 _13477_ (.A(_00301_),
    .B(net4268),
    .Y(_08033_));
 sg13g2_nor2_1 _13478_ (.A(_00283_),
    .B(net4655),
    .Y(_08034_));
 sg13g2_nor3_1 _13479_ (.A(net4715),
    .B(_08033_),
    .C(_08034_),
    .Y(_08035_));
 sg13g2_nor2_1 _13480_ (.A(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .B(net4643),
    .Y(_08036_));
 sg13g2_nor2_1 _13481_ (.A(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .B(net4653),
    .Y(_08037_));
 sg13g2_nor3_1 _13482_ (.A(_08035_),
    .B(_08036_),
    .C(_08037_),
    .Y(_08038_));
 sg13g2_or2_1 _13483_ (.X(_08039_),
    .B(net4697),
    .A(\soc_inst.spi_inst.rx_shift_reg[6] ));
 sg13g2_o21ai_1 _13484_ (.B1(_08039_),
    .Y(_08040_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .A2(net4702));
 sg13g2_a21oi_1 _13485_ (.A1(_05550_),
    .A2(net5125),
    .Y(_08041_),
    .B1(_08040_));
 sg13g2_nor2b_1 _13486_ (.A(net4798),
    .B_N(\soc_inst.i2c_inst.data_reg[6] ),
    .Y(_08042_));
 sg13g2_a21oi_1 _13487_ (.A1(\soc_inst.i2c_inst.prescale_reg[6] ),
    .A2(net4798),
    .Y(_08043_),
    .B1(_08042_));
 sg13g2_a22oi_1 _13488_ (.Y(_08044_),
    .B1(net4272),
    .B2(\soc_inst.pwm_inst.channel_duty[1][6] ),
    .A2(net4656),
    .A1(\soc_inst.pwm_inst.channel_counter[1][6] ));
 sg13g2_a22oi_1 _13489_ (.Y(_08045_),
    .B1(net4271),
    .B2(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .A2(net4656),
    .A1(\soc_inst.pwm_inst.channel_counter[0][6] ));
 sg13g2_a21oi_1 _13490_ (.A1(net8),
    .A2(net4179),
    .Y(_08046_),
    .B1(net4259));
 sg13g2_a22oi_1 _13491_ (.Y(_08047_),
    .B1(_06524_),
    .B2(\soc_inst.gpio_inst.int_pend_reg[6] ),
    .A2(net4207),
    .A1(\soc_inst.gpio_inst.int_en_reg[6] ));
 sg13g2_mux4_1 _13492_ (.S0(net4738),
    .A0(_00252_),
    .A1(_00236_),
    .A2(_08044_),
    .A3(_08045_),
    .S1(net4642),
    .X(_08048_));
 sg13g2_nor3_1 _13493_ (.A(_06294_),
    .B(_07859_),
    .C(_08043_),
    .Y(_08049_));
 sg13g2_a221oi_1 _13494_ (.B2(net4043),
    .C1(_08049_),
    .B1(_08038_),
    .A1(net4759),
    .Y(_08050_),
    .A2(_07964_));
 sg13g2_a22oi_1 _13495_ (.Y(_08051_),
    .B1(_08046_),
    .B2(_08047_),
    .A2(net4259),
    .A1(_05598_));
 sg13g2_a22oi_1 _13496_ (.Y(_08052_),
    .B1(_08051_),
    .B2(_07820_),
    .A2(_08041_),
    .A1(net3978));
 sg13g2_nor2b_1 _13497_ (.A(_08048_),
    .B_N(_07847_),
    .Y(_08053_));
 sg13g2_a221oi_1 _13498_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ),
    .C1(_08053_),
    .B1(_07962_),
    .A1(\soc_inst.spi_inst.clock_divider[6] ),
    .Y(_08054_),
    .A2(_07930_));
 sg13g2_nand4_1 _13499_ (.B(_08050_),
    .C(_08052_),
    .A(net4018),
    .Y(_08055_),
    .D(_08054_));
 sg13g2_a22oi_1 _13500_ (.Y(_08056_),
    .B1(_08032_),
    .B2(_08055_),
    .A2(net3808),
    .A1(net1465));
 sg13g2_inv_1 _13501_ (.Y(_00629_),
    .A(_08056_));
 sg13g2_nand2_1 _13502_ (.Y(_08057_),
    .A(net762),
    .B(net3809));
 sg13g2_a22oi_1 _13503_ (.Y(_08058_),
    .B1(net4704),
    .B2(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .A2(_06673_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[7] ));
 sg13g2_o21ai_1 _13504_ (.B1(_08058_),
    .Y(_08059_),
    .A1(net4757),
    .A2(_05584_));
 sg13g2_or2_1 _13505_ (.X(_08060_),
    .B(net4697),
    .A(\soc_inst.spi_inst.rx_shift_reg[7] ));
 sg13g2_o21ai_1 _13506_ (.B1(_08060_),
    .Y(_08061_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .A2(net4702));
 sg13g2_a21oi_1 _13507_ (.A1(\soc_inst.spi_inst.len_sel[1] ),
    .A2(_05603_),
    .Y(_08062_),
    .B1(_08061_));
 sg13g2_nand2_1 _13508_ (.Y(_08063_),
    .A(net4790),
    .B(\soc_inst.pwm_inst.channel_duty[1][7] ));
 sg13g2_o21ai_1 _13509_ (.B1(_08063_),
    .Y(_08064_),
    .A1(net4790),
    .A2(_05601_));
 sg13g2_mux2_1 _13510_ (.A0(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .A1(\soc_inst.pwm_inst.channel_counter[1][7] ),
    .S(net4791),
    .X(_08065_));
 sg13g2_a221oi_1 _13511_ (.B2(net4656),
    .C1(net4262),
    .B1(_08065_),
    .A1(net4272),
    .Y(_08066_),
    .A2(_08064_));
 sg13g2_mux2_1 _13512_ (.A0(_00237_),
    .A1(_00253_),
    .S(net4791),
    .X(_08067_));
 sg13g2_a21oi_2 _13513_ (.B1(_08066_),
    .Y(_08068_),
    .A2(_08067_),
    .A1(net4262));
 sg13g2_nand2_1 _13514_ (.Y(_08069_),
    .A(_00227_),
    .B(net4798));
 sg13g2_o21ai_1 _13515_ (.B1(_08069_),
    .Y(_08070_),
    .A1(net4798),
    .A2(\soc_inst.i2c_inst.data_reg[7] ));
 sg13g2_a21o_1 _13516_ (.A2(net4795),
    .A1(_00284_),
    .B1(net4655),
    .X(_08071_));
 sg13g2_o21ai_1 _13517_ (.B1(_08071_),
    .Y(_08072_),
    .A1(_00302_),
    .A2(net4268));
 sg13g2_nand2b_1 _13518_ (.Y(_08073_),
    .B(net4715),
    .A_N(\soc_inst.cpu_core.csr_file.mtime[39] ));
 sg13g2_a22oi_1 _13519_ (.Y(_08074_),
    .B1(_08072_),
    .B2(_08073_),
    .A2(_06411_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[7] ));
 sg13g2_inv_1 _13520_ (.Y(_08075_),
    .A(_08074_));
 sg13g2_nor3_1 _13521_ (.A(_06294_),
    .B(_07859_),
    .C(_08070_),
    .Y(_08076_));
 sg13g2_a221oi_1 _13522_ (.B2(net4043),
    .C1(_08076_),
    .B1(_08075_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .Y(_08077_),
    .A2(_07964_));
 sg13g2_a22oi_1 _13523_ (.Y(_08078_),
    .B1(_08068_),
    .B2(_07847_),
    .A2(_07962_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ));
 sg13g2_a22oi_1 _13524_ (.Y(_08079_),
    .B1(_08062_),
    .B2(_07929_),
    .A2(_07930_),
    .A1(\soc_inst.spi_inst.clock_divider[7] ));
 sg13g2_nand4_1 _13525_ (.B(_08077_),
    .C(_08078_),
    .A(net4018),
    .Y(_08080_),
    .D(_08079_));
 sg13g2_o21ai_1 _13526_ (.B1(_08080_),
    .Y(_08081_),
    .A1(net4016),
    .A2(_08059_));
 sg13g2_o21ai_1 _13527_ (.B1(_08057_),
    .Y(_00630_),
    .A1(net3809),
    .A2(_08081_));
 sg13g2_nor2_1 _13528_ (.A(_00303_),
    .B(net4266),
    .Y(_08082_));
 sg13g2_nor2_1 _13529_ (.A(_00285_),
    .B(net4654),
    .Y(_08083_));
 sg13g2_nor3_1 _13530_ (.A(net4713),
    .B(_08082_),
    .C(_08083_),
    .Y(_08084_));
 sg13g2_nor2_1 _13531_ (.A(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .B(net4641),
    .Y(_08085_));
 sg13g2_nor2_1 _13532_ (.A(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .B(net4647),
    .Y(_08086_));
 sg13g2_nor3_1 _13533_ (.A(_08084_),
    .B(_08085_),
    .C(_08086_),
    .Y(_08087_));
 sg13g2_nand2_1 _13534_ (.Y(_08088_),
    .A(net4738),
    .B(_05604_));
 sg13g2_o21ai_1 _13535_ (.B1(_08088_),
    .Y(_08089_),
    .A1(net4738),
    .A2(\soc_inst.pwm_inst.channel_duty[1][8] ));
 sg13g2_a21oi_1 _13536_ (.A1(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .A2(net4277),
    .Y(_08090_),
    .B1(net4791));
 sg13g2_o21ai_1 _13537_ (.B1(_08090_),
    .Y(_08091_),
    .A1(_00238_),
    .A2(net4642));
 sg13g2_nor2_1 _13538_ (.A(_05571_),
    .B(_06296_),
    .Y(_08092_));
 sg13g2_o21ai_1 _13539_ (.B1(net4791),
    .Y(_08093_),
    .A1(_00254_),
    .A2(net4642));
 sg13g2_o21ai_1 _13540_ (.B1(_08091_),
    .Y(_08094_),
    .A1(_08092_),
    .A2(_08093_));
 sg13g2_o21ai_1 _13541_ (.B1(_08094_),
    .Y(_08095_),
    .A1(net4270),
    .A2(_08089_));
 sg13g2_and2_1 _13542_ (.A(net5125),
    .B(_07908_),
    .X(_08096_));
 sg13g2_a221oi_1 _13543_ (.B2(net4705),
    .C1(net4016),
    .B1(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .A1(net4875),
    .Y(_08097_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[16] ));
 sg13g2_a22oi_1 _13544_ (.Y(_08098_),
    .B1(_08095_),
    .B2(net4044),
    .A2(_08087_),
    .A1(net4043));
 sg13g2_a22oi_1 _13545_ (.Y(_08099_),
    .B1(_07964_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .A2(_07930_),
    .A1(\soc_inst.spi_inst.cpha ));
 sg13g2_a22oi_1 _13546_ (.Y(_08100_),
    .B1(_06939_),
    .B2(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .A2(net5125),
    .A1(\soc_inst.spi_inst.rx_shift_reg[16] ));
 sg13g2_nand2b_1 _13547_ (.Y(_08101_),
    .B(net3978),
    .A_N(_08100_));
 sg13g2_and4_1 _13548_ (.A(net4018),
    .B(_08098_),
    .C(_08099_),
    .D(_08101_),
    .X(_08102_));
 sg13g2_nor3_1 _13549_ (.A(net3806),
    .B(_08097_),
    .C(_08102_),
    .Y(_08103_));
 sg13g2_a21o_1 _13550_ (.A2(net3806),
    .A1(net591),
    .B1(_08103_),
    .X(_00631_));
 sg13g2_a221oi_1 _13551_ (.B2(net4705),
    .C1(net4015),
    .B1(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .A1(net4873),
    .Y(_08104_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[17] ));
 sg13g2_nor2_1 _13552_ (.A(_00304_),
    .B(net4266),
    .Y(_08105_));
 sg13g2_nor2_1 _13553_ (.A(_00286_),
    .B(net4654),
    .Y(_08106_));
 sg13g2_nor3_1 _13554_ (.A(net4713),
    .B(_08105_),
    .C(_08106_),
    .Y(_08107_));
 sg13g2_a221oi_1 _13555_ (.B2(_05514_),
    .C1(_08107_),
    .B1(net4264),
    .A1(_05511_),
    .Y(_08108_),
    .A2(_06411_));
 sg13g2_a22oi_1 _13556_ (.Y(_08109_),
    .B1(net4271),
    .B2(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .A2(net4656),
    .A1(\soc_inst.pwm_inst.channel_counter[0][9] ));
 sg13g2_nor2_1 _13557_ (.A(net4788),
    .B(_08109_),
    .Y(_08110_));
 sg13g2_a22oi_1 _13558_ (.Y(_08111_),
    .B1(net4271),
    .B2(\soc_inst.pwm_inst.channel_duty[1][9] ),
    .A2(net4656),
    .A1(\soc_inst.pwm_inst.channel_counter[1][9] ));
 sg13g2_o21ai_1 _13559_ (.B1(net4641),
    .Y(_08112_),
    .A1(net4738),
    .A2(_08111_));
 sg13g2_nor2_1 _13560_ (.A(_08110_),
    .B(_08112_),
    .Y(_08113_));
 sg13g2_mux2_1 _13561_ (.A0(_00239_),
    .A1(_00255_),
    .S(net4788),
    .X(_08114_));
 sg13g2_a21oi_2 _13562_ (.B1(_08113_),
    .Y(_08115_),
    .A2(_08114_),
    .A1(net4263));
 sg13g2_a22oi_1 _13563_ (.Y(_08116_),
    .B1(_08115_),
    .B2(_07847_),
    .A2(_07964_),
    .A1(_05387_));
 sg13g2_and2_1 _13564_ (.A(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .B(_06939_),
    .X(_08117_));
 sg13g2_a22oi_1 _13565_ (.Y(_08118_),
    .B1(_08117_),
    .B2(net3978),
    .A2(_08108_),
    .A1(_07862_));
 sg13g2_and2_1 _13566_ (.A(net5126),
    .B(_07929_),
    .X(_08119_));
 sg13g2_a22oi_1 _13567_ (.Y(_08120_),
    .B1(_08119_),
    .B2(\soc_inst.spi_inst.rx_shift_reg[17] ),
    .A2(_07930_),
    .A1(\soc_inst.spi_inst.cpol ));
 sg13g2_and4_1 _13568_ (.A(_05904_),
    .B(_08116_),
    .C(_08118_),
    .D(_08120_),
    .X(_08121_));
 sg13g2_nor3_1 _13569_ (.A(net3807),
    .B(_08104_),
    .C(_08121_),
    .Y(_08122_));
 sg13g2_a21o_1 _13570_ (.A2(net3806),
    .A1(net594),
    .B1(_08122_),
    .X(_00632_));
 sg13g2_mux2_1 _13571_ (.A0(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[18] ),
    .S(_06940_),
    .X(_08123_));
 sg13g2_and2_1 _13572_ (.A(net4697),
    .B(_07908_),
    .X(_08124_));
 sg13g2_a21oi_1 _13573_ (.A1(_05399_),
    .A2(net4656),
    .Y(_08125_),
    .B1(net4714));
 sg13g2_o21ai_1 _13574_ (.B1(_08125_),
    .Y(_08126_),
    .A1(_00305_),
    .A2(net4266));
 sg13g2_o21ai_1 _13575_ (.B1(_08126_),
    .Y(_08127_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .A2(net4641));
 sg13g2_a21oi_1 _13576_ (.A1(_05510_),
    .A2(_06411_),
    .Y(_08128_),
    .B1(_08127_));
 sg13g2_mux2_1 _13577_ (.A0(_00240_),
    .A1(_00256_),
    .S(net4788),
    .X(_08129_));
 sg13g2_nor2_1 _13578_ (.A(net4788),
    .B(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .Y(_08130_));
 sg13g2_a21oi_1 _13579_ (.A1(net4788),
    .A2(_05606_),
    .Y(_08131_),
    .B1(_08130_));
 sg13g2_mux2_1 _13580_ (.A0(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .A1(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .S(net4788),
    .X(_08132_));
 sg13g2_a221oi_1 _13581_ (.B2(net4277),
    .C1(net4263),
    .B1(_08132_),
    .A1(net4271),
    .Y(_08133_),
    .A2(_08131_));
 sg13g2_a21oi_2 _13582_ (.B1(_08133_),
    .Y(_08134_),
    .A2(_08129_),
    .A1(net4263));
 sg13g2_a22oi_1 _13583_ (.Y(_08135_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .B2(net4705),
    .A2(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .A1(net4873));
 sg13g2_nand3_1 _13584_ (.B(net3978),
    .C(_08123_),
    .A(_07825_),
    .Y(_08136_));
 sg13g2_a221oi_1 _13585_ (.B2(net4044),
    .C1(_05905_),
    .B1(_08134_),
    .A1(_07862_),
    .Y(_08137_),
    .A2(_08128_));
 sg13g2_a221oi_1 _13586_ (.B2(_08137_),
    .C1(net3808),
    .B1(_08136_),
    .A1(_05905_),
    .Y(_08138_),
    .A2(_08135_));
 sg13g2_a21o_1 _13587_ (.A2(net3808),
    .A1(net989),
    .B1(_08138_),
    .X(_00633_));
 sg13g2_mux2_1 _13588_ (.A0(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[19] ),
    .S(net4701),
    .X(_08139_));
 sg13g2_mux4_1 _13589_ (.S0(net4789),
    .A0(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .A1(\soc_inst.pwm_inst.channel_duty[1][11] ),
    .A2(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .A3(\soc_inst.pwm_inst.channel_counter[1][11] ),
    .S1(net4797),
    .X(_08140_));
 sg13g2_or2_1 _13590_ (.X(_08141_),
    .B(net4788),
    .A(_00241_));
 sg13g2_o21ai_1 _13591_ (.B1(_08141_),
    .Y(_08142_),
    .A1(_00257_),
    .A2(net4739));
 sg13g2_a22oi_1 _13592_ (.Y(_08143_),
    .B1(_08142_),
    .B2(net4263),
    .A2(_08140_),
    .A1(_06293_));
 sg13g2_nor2_1 _13593_ (.A(_00306_),
    .B(net4266),
    .Y(_08144_));
 sg13g2_nor2_1 _13594_ (.A(_00288_),
    .B(net4654),
    .Y(_08145_));
 sg13g2_nor3_1 _13595_ (.A(net4713),
    .B(_08144_),
    .C(_08145_),
    .Y(_08146_));
 sg13g2_nor2_1 _13596_ (.A(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .B(net4647),
    .Y(_08147_));
 sg13g2_nor2_1 _13597_ (.A(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .B(net4641),
    .Y(_08148_));
 sg13g2_nor4_1 _13598_ (.A(net4045),
    .B(_08146_),
    .C(_08147_),
    .D(_08148_),
    .Y(_08149_));
 sg13g2_nor2_1 _13599_ (.A(net4066),
    .B(_08149_),
    .Y(_08150_));
 sg13g2_o21ai_1 _13600_ (.B1(_08150_),
    .Y(_08151_),
    .A1(_07846_),
    .A2(_08143_));
 sg13g2_a21oi_1 _13601_ (.A1(_08124_),
    .A2(_08139_),
    .Y(_08152_),
    .B1(_08151_));
 sg13g2_a221oi_1 _13602_ (.B2(net4705),
    .C1(net4016),
    .B1(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .A1(net4875),
    .Y(_08153_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[19] ));
 sg13g2_nor3_1 _13603_ (.A(net3807),
    .B(_08152_),
    .C(_08153_),
    .Y(_08154_));
 sg13g2_a21o_1 _13604_ (.A2(net3807),
    .A1(net607),
    .B1(_08154_),
    .X(_00634_));
 sg13g2_mux2_1 _13605_ (.A0(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[20] ),
    .S(net4701),
    .X(_08155_));
 sg13g2_mux4_1 _13606_ (.S0(net4788),
    .A0(\soc_inst.pwm_inst.channel_duty[0][12] ),
    .A1(\soc_inst.pwm_inst.channel_duty[1][12] ),
    .A2(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .A3(\soc_inst.pwm_inst.channel_counter[1][12] ),
    .S1(net4797),
    .X(_08156_));
 sg13g2_or2_1 _13607_ (.X(_08157_),
    .B(net4789),
    .A(_00242_));
 sg13g2_o21ai_1 _13608_ (.B1(_08157_),
    .Y(_08158_),
    .A1(_00258_),
    .A2(net4739));
 sg13g2_a22oi_1 _13609_ (.Y(_08159_),
    .B1(_08158_),
    .B2(net4263),
    .A2(_08156_),
    .A1(_06293_));
 sg13g2_nor2_1 _13610_ (.A(_00307_),
    .B(net4266),
    .Y(_08160_));
 sg13g2_nor2_1 _13611_ (.A(_00289_),
    .B(net4654),
    .Y(_08161_));
 sg13g2_nor3_1 _13612_ (.A(net4713),
    .B(_08160_),
    .C(_08161_),
    .Y(_08162_));
 sg13g2_nor2_1 _13613_ (.A(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .B(net4647),
    .Y(_08163_));
 sg13g2_nor2_1 _13614_ (.A(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .B(net4641),
    .Y(_08164_));
 sg13g2_nor4_1 _13615_ (.A(net4046),
    .B(_08162_),
    .C(_08163_),
    .D(_08164_),
    .Y(_08165_));
 sg13g2_nor2_1 _13616_ (.A(net4066),
    .B(_08165_),
    .Y(_08166_));
 sg13g2_o21ai_1 _13617_ (.B1(_08166_),
    .Y(_08167_),
    .A1(_07846_),
    .A2(_08159_));
 sg13g2_a21oi_1 _13618_ (.A1(_08124_),
    .A2(_08155_),
    .Y(_08168_),
    .B1(_08167_));
 sg13g2_a221oi_1 _13619_ (.B2(net4705),
    .C1(net4016),
    .B1(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .A1(net4875),
    .Y(_08169_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[20] ));
 sg13g2_nor3_1 _13620_ (.A(net3806),
    .B(_08168_),
    .C(_08169_),
    .Y(_08170_));
 sg13g2_a21o_1 _13621_ (.A2(net3807),
    .A1(net593),
    .B1(_08170_),
    .X(_00635_));
 sg13g2_mux2_1 _13622_ (.A0(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[21] ),
    .S(net4701),
    .X(_08171_));
 sg13g2_mux4_1 _13623_ (.S0(net4789),
    .A0(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .A1(\soc_inst.pwm_inst.channel_duty[1][13] ),
    .A2(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .A3(\soc_inst.pwm_inst.channel_counter[1][13] ),
    .S1(net4797),
    .X(_08172_));
 sg13g2_or2_1 _13624_ (.X(_08173_),
    .B(net4789),
    .A(_00243_));
 sg13g2_o21ai_1 _13625_ (.B1(_08173_),
    .Y(_08174_),
    .A1(_00259_),
    .A2(net4738));
 sg13g2_a22oi_1 _13626_ (.Y(_08175_),
    .B1(_08174_),
    .B2(net4263),
    .A2(_08172_),
    .A1(_06293_));
 sg13g2_nor2_1 _13627_ (.A(_00308_),
    .B(net4266),
    .Y(_08176_));
 sg13g2_nor2_1 _13628_ (.A(_00290_),
    .B(net4654),
    .Y(_08177_));
 sg13g2_nor3_1 _13629_ (.A(net4713),
    .B(_08176_),
    .C(_08177_),
    .Y(_08178_));
 sg13g2_nor2_1 _13630_ (.A(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .B(net4647),
    .Y(_08179_));
 sg13g2_nor2_1 _13631_ (.A(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .B(net4641),
    .Y(_08180_));
 sg13g2_nor4_1 _13632_ (.A(net4046),
    .B(_08178_),
    .C(_08179_),
    .D(_08180_),
    .Y(_08181_));
 sg13g2_nor2_1 _13633_ (.A(_05886_),
    .B(_08181_),
    .Y(_08182_));
 sg13g2_o21ai_1 _13634_ (.B1(_08182_),
    .Y(_08183_),
    .A1(_07846_),
    .A2(_08175_));
 sg13g2_a21oi_1 _13635_ (.A1(_08124_),
    .A2(_08171_),
    .Y(_08184_),
    .B1(_08183_));
 sg13g2_a221oi_1 _13636_ (.B2(net4705),
    .C1(net4017),
    .B1(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .A1(\soc_inst.core_mem_flag[1] ),
    .Y(_08185_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[21] ));
 sg13g2_nor3_1 _13637_ (.A(net3806),
    .B(_08184_),
    .C(_08185_),
    .Y(_08186_));
 sg13g2_a21o_1 _13638_ (.A2(net3806),
    .A1(net674),
    .B1(_08186_),
    .X(_00636_));
 sg13g2_mux2_1 _13639_ (.A0(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[22] ),
    .S(net4701),
    .X(_08187_));
 sg13g2_mux4_1 _13640_ (.S0(net4793),
    .A0(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .A1(\soc_inst.pwm_inst.channel_duty[1][14] ),
    .A2(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .A3(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .S1(net4797),
    .X(_08188_));
 sg13g2_or2_1 _13641_ (.X(_08189_),
    .B(net4793),
    .A(_00244_));
 sg13g2_o21ai_1 _13642_ (.B1(_08189_),
    .Y(_08190_),
    .A1(_00260_),
    .A2(net4739));
 sg13g2_a22oi_1 _13643_ (.Y(_08191_),
    .B1(_08190_),
    .B2(net4262),
    .A2(_08188_),
    .A1(_06293_));
 sg13g2_nor2_1 _13644_ (.A(_00309_),
    .B(net4266),
    .Y(_08192_));
 sg13g2_nor2_1 _13645_ (.A(_00291_),
    .B(net4654),
    .Y(_08193_));
 sg13g2_nor3_1 _13646_ (.A(net4713),
    .B(_08192_),
    .C(_08193_),
    .Y(_08194_));
 sg13g2_nor2_1 _13647_ (.A(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .B(net4647),
    .Y(_08195_));
 sg13g2_nor2_1 _13648_ (.A(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .B(net4641),
    .Y(_08196_));
 sg13g2_nor4_1 _13649_ (.A(net4046),
    .B(_08194_),
    .C(_08195_),
    .D(_08196_),
    .Y(_08197_));
 sg13g2_nor2_1 _13650_ (.A(net4066),
    .B(_08197_),
    .Y(_08198_));
 sg13g2_o21ai_1 _13651_ (.B1(_08198_),
    .Y(_08199_),
    .A1(_07846_),
    .A2(_08191_));
 sg13g2_a21oi_1 _13652_ (.A1(_08124_),
    .A2(_08187_),
    .Y(_08200_),
    .B1(_08199_));
 sg13g2_a221oi_1 _13653_ (.B2(net4706),
    .C1(net4016),
    .B1(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .A1(net4875),
    .Y(_08201_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[22] ));
 sg13g2_nor3_1 _13654_ (.A(net3806),
    .B(_08200_),
    .C(_08201_),
    .Y(_08202_));
 sg13g2_a21o_1 _13655_ (.A2(net3807),
    .A1(net651),
    .B1(_08202_),
    .X(_00637_));
 sg13g2_mux2_1 _13656_ (.A0(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[23] ),
    .S(net4701),
    .X(_08203_));
 sg13g2_mux4_1 _13657_ (.S0(net4789),
    .A0(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .A1(\soc_inst.pwm_inst.channel_duty[1][15] ),
    .A2(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .A3(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .S1(net4797),
    .X(_08204_));
 sg13g2_or2_1 _13658_ (.X(_08205_),
    .B(net4793),
    .A(_00245_));
 sg13g2_o21ai_1 _13659_ (.B1(_08205_),
    .Y(_08206_),
    .A1(_00261_),
    .A2(net4739));
 sg13g2_a22oi_1 _13660_ (.Y(_08207_),
    .B1(_08206_),
    .B2(net4263),
    .A2(_08204_),
    .A1(_06293_));
 sg13g2_nor2_1 _13661_ (.A(_00310_),
    .B(net4266),
    .Y(_08208_));
 sg13g2_nor2_1 _13662_ (.A(_00292_),
    .B(net4654),
    .Y(_08209_));
 sg13g2_nor3_1 _13663_ (.A(net4713),
    .B(_08208_),
    .C(_08209_),
    .Y(_08210_));
 sg13g2_nor2_1 _13664_ (.A(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .B(net4647),
    .Y(_08211_));
 sg13g2_nor2_1 _13665_ (.A(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .B(net4641),
    .Y(_08212_));
 sg13g2_nor4_1 _13666_ (.A(net4046),
    .B(_08210_),
    .C(_08211_),
    .D(_08212_),
    .Y(_08213_));
 sg13g2_nor2_1 _13667_ (.A(net4066),
    .B(_08213_),
    .Y(_08214_));
 sg13g2_o21ai_1 _13668_ (.B1(_08214_),
    .Y(_08215_),
    .A1(_07846_),
    .A2(_08207_));
 sg13g2_a21oi_1 _13669_ (.A1(_08124_),
    .A2(_08203_),
    .Y(_08216_),
    .B1(_08215_));
 sg13g2_a221oi_1 _13670_ (.B2(net4706),
    .C1(net4016),
    .B1(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .A1(net4875),
    .Y(_08217_),
    .A2(\soc_inst.mem_ctrl.spi_data_out[23] ));
 sg13g2_nor3_1 _13671_ (.A(net3806),
    .B(_08216_),
    .C(_08217_),
    .Y(_08218_));
 sg13g2_a21o_1 _13672_ (.A2(net3807),
    .A1(net1571),
    .B1(_08218_),
    .X(_00638_));
 sg13g2_nand3_1 _13673_ (.B(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .C(_05905_),
    .A(net4875),
    .Y(_08219_));
 sg13g2_o21ai_1 _13674_ (.B1(net4646),
    .Y(_08220_),
    .A1(_00311_),
    .A2(net4265));
 sg13g2_o21ai_1 _13675_ (.B1(_08220_),
    .Y(_08221_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .A2(net4646));
 sg13g2_o21ai_1 _13676_ (.B1(_08219_),
    .Y(_08222_),
    .A1(net4047),
    .A2(_08221_));
 sg13g2_a21oi_1 _13677_ (.A1(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .A2(net4041),
    .Y(_08223_),
    .B1(_08222_));
 sg13g2_nor2_1 _13678_ (.A(net1436),
    .B(net3812),
    .Y(_08224_));
 sg13g2_a21oi_1 _13679_ (.A1(net3812),
    .A2(_08223_),
    .Y(_00639_),
    .B1(_08224_));
 sg13g2_nor2_1 _13680_ (.A(net1641),
    .B(net3811),
    .Y(_08225_));
 sg13g2_and2_1 _13681_ (.A(net4875),
    .B(_05886_),
    .X(_08226_));
 sg13g2_o21ai_1 _13682_ (.B1(net4646),
    .Y(_08227_),
    .A1(_00312_),
    .A2(net4265));
 sg13g2_o21ai_1 _13683_ (.B1(_08227_),
    .Y(_08228_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .A2(net4646));
 sg13g2_nor2_1 _13684_ (.A(net4045),
    .B(_08228_),
    .Y(_08229_));
 sg13g2_a221oi_1 _13685_ (.B2(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .C1(_08229_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .Y(_08230_),
    .A2(net4042));
 sg13g2_a21oi_1 _13686_ (.A1(net3811),
    .A2(_08230_),
    .Y(_00640_),
    .B1(_08225_));
 sg13g2_o21ai_1 _13687_ (.B1(net4645),
    .Y(_08231_),
    .A1(_00313_),
    .A2(net4265));
 sg13g2_o21ai_1 _13688_ (.B1(_08231_),
    .Y(_08232_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .A2(net4645));
 sg13g2_nor2_1 _13689_ (.A(net4045),
    .B(_08232_),
    .Y(_08233_));
 sg13g2_a221oi_1 _13690_ (.B2(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .C1(_08233_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .Y(_08234_),
    .A2(net4041));
 sg13g2_nor2_1 _13691_ (.A(net1320),
    .B(net3810),
    .Y(_08235_));
 sg13g2_a21oi_1 _13692_ (.A1(net3810),
    .A2(_08234_),
    .Y(_00641_),
    .B1(_08235_));
 sg13g2_o21ai_1 _13693_ (.B1(net4645),
    .Y(_08236_),
    .A1(_00314_),
    .A2(net4265));
 sg13g2_o21ai_1 _13694_ (.B1(_08236_),
    .Y(_08237_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .A2(net4645));
 sg13g2_nor2_1 _13695_ (.A(net4045),
    .B(_08237_),
    .Y(_08238_));
 sg13g2_a221oi_1 _13696_ (.B2(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .C1(_08238_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .Y(_08239_),
    .A2(net4042));
 sg13g2_nor2_1 _13697_ (.A(net745),
    .B(net3811),
    .Y(_08240_));
 sg13g2_a21oi_1 _13698_ (.A1(net3811),
    .A2(_08239_),
    .Y(_00642_),
    .B1(_08240_));
 sg13g2_o21ai_1 _13699_ (.B1(net4645),
    .Y(_08241_),
    .A1(_00315_),
    .A2(net4265));
 sg13g2_o21ai_1 _13700_ (.B1(_08241_),
    .Y(_08242_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .A2(net4645));
 sg13g2_nor2_1 _13701_ (.A(net4045),
    .B(_08242_),
    .Y(_08243_));
 sg13g2_a221oi_1 _13702_ (.B2(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .C1(_08243_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .Y(_08244_),
    .A2(net4041));
 sg13g2_nor2_1 _13703_ (.A(net753),
    .B(net3812),
    .Y(_08245_));
 sg13g2_a21oi_1 _13704_ (.A1(net3812),
    .A2(_08244_),
    .Y(_00643_),
    .B1(_08245_));
 sg13g2_o21ai_1 _13705_ (.B1(net4645),
    .Y(_08246_),
    .A1(_00316_),
    .A2(net4265));
 sg13g2_o21ai_1 _13706_ (.B1(_08246_),
    .Y(_08247_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .A2(net4646));
 sg13g2_nor2_1 _13707_ (.A(net4045),
    .B(_08247_),
    .Y(_08248_));
 sg13g2_a221oi_1 _13708_ (.B2(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .C1(_08248_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .Y(_08249_),
    .A2(net4041));
 sg13g2_nor2_1 _13709_ (.A(net551),
    .B(net3811),
    .Y(_08250_));
 sg13g2_a21oi_1 _13710_ (.A1(net3811),
    .A2(_08249_),
    .Y(_00644_),
    .B1(_08250_));
 sg13g2_o21ai_1 _13711_ (.B1(net4645),
    .Y(_08251_),
    .A1(_00317_),
    .A2(net4265));
 sg13g2_o21ai_1 _13712_ (.B1(_08251_),
    .Y(_08252_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .A2(net4647));
 sg13g2_nor2_1 _13713_ (.A(net4045),
    .B(_08252_),
    .Y(_08253_));
 sg13g2_a221oi_1 _13714_ (.B2(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .C1(_08253_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .Y(_08254_),
    .A2(net4041));
 sg13g2_nor2_1 _13715_ (.A(net635),
    .B(net3810),
    .Y(_08255_));
 sg13g2_a21oi_1 _13716_ (.A1(net3810),
    .A2(_08254_),
    .Y(_00645_),
    .B1(_08255_));
 sg13g2_nor2_1 _13717_ (.A(net902),
    .B(net3810),
    .Y(_08256_));
 sg13g2_o21ai_1 _13718_ (.B1(net4646),
    .Y(_08257_),
    .A1(_00318_),
    .A2(net4265));
 sg13g2_o21ai_1 _13719_ (.B1(_08257_),
    .Y(_08258_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .A2(net4646));
 sg13g2_nor2_1 _13720_ (.A(net4045),
    .B(_08258_),
    .Y(_08259_));
 sg13g2_a221oi_1 _13721_ (.B2(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .C1(_08259_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .Y(_08260_),
    .A2(net4041));
 sg13g2_a21oi_1 _13722_ (.A1(net3810),
    .A2(_08260_),
    .Y(_00646_),
    .B1(_08256_));
 sg13g2_o21ai_1 _13723_ (.B1(net4648),
    .Y(_08261_),
    .A1(_00319_),
    .A2(net4267));
 sg13g2_o21ai_1 _13724_ (.B1(_08261_),
    .Y(_08262_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .A2(net4648));
 sg13g2_nor2_1 _13725_ (.A(net4047),
    .B(_08262_),
    .Y(_08263_));
 sg13g2_a21oi_1 _13726_ (.A1(net2353),
    .A2(net4042),
    .Y(_08264_),
    .B1(_08263_));
 sg13g2_nand3_1 _13727_ (.B(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .C(_05886_),
    .A(net4875),
    .Y(_08265_));
 sg13g2_nand3_1 _13728_ (.B(_08264_),
    .C(_08265_),
    .A(net3815),
    .Y(_08266_));
 sg13g2_o21ai_1 _13729_ (.B1(_08266_),
    .Y(_08267_),
    .A1(net2416),
    .A2(net3815));
 sg13g2_inv_1 _13730_ (.Y(_00647_),
    .A(_08267_));
 sg13g2_o21ai_1 _13731_ (.B1(net4650),
    .Y(_08268_),
    .A1(_00320_),
    .A2(net4267));
 sg13g2_o21ai_1 _13732_ (.B1(_08268_),
    .Y(_08269_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .A2(net4650));
 sg13g2_nor2_1 _13733_ (.A(net4047),
    .B(_08269_),
    .Y(_08270_));
 sg13g2_a221oi_1 _13734_ (.B2(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .C1(_08270_),
    .B1(net3977),
    .A1(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .Y(_08271_),
    .A2(net4042));
 sg13g2_nor2_1 _13735_ (.A(net1511),
    .B(net3815),
    .Y(_08272_));
 sg13g2_a21oi_1 _13736_ (.A1(net3815),
    .A2(_08271_),
    .Y(_00648_),
    .B1(_08272_));
 sg13g2_nor2_1 _13737_ (.A(net1540),
    .B(net3815),
    .Y(_08273_));
 sg13g2_o21ai_1 _13738_ (.B1(net4650),
    .Y(_08274_),
    .A1(_00321_),
    .A2(net4267));
 sg13g2_o21ai_1 _13739_ (.B1(_08274_),
    .Y(_08275_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .A2(net4648));
 sg13g2_nor2_1 _13740_ (.A(net4047),
    .B(_08275_),
    .Y(_08276_));
 sg13g2_a221oi_1 _13741_ (.B2(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .C1(_08276_),
    .B1(net3977),
    .A1(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .Y(_08277_),
    .A2(net4042));
 sg13g2_a21oi_1 _13742_ (.A1(net3816),
    .A2(_08277_),
    .Y(_00649_),
    .B1(_08273_));
 sg13g2_nor2_1 _13743_ (.A(net639),
    .B(net3810),
    .Y(_08278_));
 sg13g2_o21ai_1 _13744_ (.B1(net4649),
    .Y(_08279_),
    .A1(_00322_),
    .A2(net4267));
 sg13g2_o21ai_1 _13745_ (.B1(_08279_),
    .Y(_08280_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .A2(net4649));
 sg13g2_nor2_1 _13746_ (.A(net4047),
    .B(_08280_),
    .Y(_08281_));
 sg13g2_a221oi_1 _13747_ (.B2(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .C1(_08281_),
    .B1(net3977),
    .A1(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .Y(_08282_),
    .A2(_08096_));
 sg13g2_a21oi_1 _13748_ (.A1(net3814),
    .A2(_08282_),
    .Y(_00650_),
    .B1(_08278_));
 sg13g2_nor2_1 _13749_ (.A(net1466),
    .B(net3813),
    .Y(_08283_));
 sg13g2_o21ai_1 _13750_ (.B1(net4649),
    .Y(_08284_),
    .A1(_00323_),
    .A2(net4267));
 sg13g2_o21ai_1 _13751_ (.B1(_08284_),
    .Y(_08285_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .A2(net4648));
 sg13g2_nor2_1 _13752_ (.A(net4047),
    .B(_08285_),
    .Y(_08286_));
 sg13g2_a221oi_1 _13753_ (.B2(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .C1(_08286_),
    .B1(net3977),
    .A1(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .Y(_08287_),
    .A2(net4042));
 sg13g2_a21oi_1 _13754_ (.A1(net3813),
    .A2(_08287_),
    .Y(_00651_),
    .B1(_08283_));
 sg13g2_nor2_1 _13755_ (.A(net1179),
    .B(net3811),
    .Y(_08288_));
 sg13g2_o21ai_1 _13756_ (.B1(net4650),
    .Y(_08289_),
    .A1(_00324_),
    .A2(net4267));
 sg13g2_o21ai_1 _13757_ (.B1(_08289_),
    .Y(_08290_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .A2(net4650));
 sg13g2_nor2_1 _13758_ (.A(net4047),
    .B(_08290_),
    .Y(_08291_));
 sg13g2_a221oi_1 _13759_ (.B2(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .C1(_08291_),
    .B1(net3976),
    .A1(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .Y(_08292_),
    .A2(net4041));
 sg13g2_a21oi_1 _13760_ (.A1(net3811),
    .A2(_08292_),
    .Y(_00652_),
    .B1(_08288_));
 sg13g2_o21ai_1 _13761_ (.B1(net4648),
    .Y(_08293_),
    .A1(_00325_),
    .A2(net4267));
 sg13g2_o21ai_1 _13762_ (.B1(_08293_),
    .Y(_08294_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .A2(net4648));
 sg13g2_nor2_1 _13763_ (.A(net4047),
    .B(_08294_),
    .Y(_08295_));
 sg13g2_a221oi_1 _13764_ (.B2(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .C1(_08295_),
    .B1(net3977),
    .A1(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .Y(_08296_),
    .A2(net4042));
 sg13g2_nor2_1 _13765_ (.A(net500),
    .B(net3815),
    .Y(_08297_));
 sg13g2_a21oi_1 _13766_ (.A1(net3815),
    .A2(_08296_),
    .Y(_00653_),
    .B1(_08297_));
 sg13g2_o21ai_1 _13767_ (.B1(net4648),
    .Y(_08298_),
    .A1(_00326_),
    .A2(net4267));
 sg13g2_o21ai_1 _13768_ (.B1(_08298_),
    .Y(_08299_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .A2(net4648));
 sg13g2_nor2_1 _13769_ (.A(net4048),
    .B(_08299_),
    .Y(_08300_));
 sg13g2_a221oi_1 _13770_ (.B2(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .C1(_08300_),
    .B1(net3977),
    .A1(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .Y(_08301_),
    .A2(net4041));
 sg13g2_nor2_1 _13771_ (.A(net1574),
    .B(net3810),
    .Y(_08302_));
 sg13g2_a21oi_1 _13772_ (.A1(net3814),
    .A2(_08301_),
    .Y(_00654_),
    .B1(_08302_));
 sg13g2_nand2_1 _13773_ (.Y(_08303_),
    .A(_05872_),
    .B(_06025_));
 sg13g2_nor2_1 _13774_ (.A(net4779),
    .B(net2566),
    .Y(_08304_));
 sg13g2_nand3_1 _13775_ (.B(_05872_),
    .C(_08304_),
    .A(_00276_),
    .Y(_08305_));
 sg13g2_nand4_1 _13776_ (.B(_06030_),
    .C(_08303_),
    .A(_06019_),
    .Y(_08306_),
    .D(_08305_));
 sg13g2_o21ai_1 _13777_ (.B1(\soc_inst.core_mem_re ),
    .Y(_08307_),
    .A1(net5074),
    .A2(net4779));
 sg13g2_nand2b_1 _13778_ (.Y(_08308_),
    .B(_08304_),
    .A_N(net5075));
 sg13g2_and2_1 _13779_ (.A(_08307_),
    .B(_08308_),
    .X(_08309_));
 sg13g2_nor3_1 _13780_ (.A(_05867_),
    .B(_08306_),
    .C(_08309_),
    .Y(_08310_));
 sg13g2_a21o_1 _13781_ (.A2(_08306_),
    .A1(net599),
    .B1(_08310_),
    .X(_00655_));
 sg13g2_a21oi_1 _13782_ (.A1(_05906_),
    .A2(_07542_),
    .Y(_08311_),
    .B1(_07807_));
 sg13g2_o21ai_1 _13783_ (.B1(_08311_),
    .Y(_08312_),
    .A1(net4017),
    .A2(_07541_));
 sg13g2_o21ai_1 _13784_ (.B1(_08312_),
    .Y(_00656_),
    .A1(_05719_),
    .A2(_08311_));
 sg13g2_nor3_1 _13785_ (.A(_06032_),
    .B(_07538_),
    .C(_07542_),
    .Y(_08313_));
 sg13g2_a21oi_1 _13786_ (.A1(net4772),
    .A2(_06013_),
    .Y(_08314_),
    .B1(\soc_inst.mem_ctrl.access_state[3] ));
 sg13g2_nor2_1 _13787_ (.A(net641),
    .B(_08313_),
    .Y(_08315_));
 sg13g2_a21oi_1 _13788_ (.A1(_08313_),
    .A2(_08314_),
    .Y(_00657_),
    .B1(_08315_));
 sg13g2_nor2_1 _13789_ (.A(net4780),
    .B(_07530_),
    .Y(_08316_));
 sg13g2_nor2_1 _13790_ (.A(_07539_),
    .B(_08316_),
    .Y(_08317_));
 sg13g2_nand3_1 _13791_ (.B(_07545_),
    .C(_08317_),
    .A(_07529_),
    .Y(_08318_));
 sg13g2_nand2_1 _13792_ (.Y(_08319_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[24] ));
 sg13g2_nand2_1 _13793_ (.Y(_08320_),
    .A(net241),
    .B(net3692));
 sg13g2_o21ai_1 _13794_ (.B1(_08320_),
    .Y(_00658_),
    .A1(net3692),
    .A2(_08319_));
 sg13g2_nand2_1 _13795_ (.Y(_08321_),
    .A(net4780),
    .B(\soc_inst.mem_ctrl.spi_data_out[25] ));
 sg13g2_nand2_1 _13796_ (.Y(_08322_),
    .A(net211),
    .B(net3693));
 sg13g2_o21ai_1 _13797_ (.B1(_08322_),
    .Y(_00659_),
    .A1(net3693),
    .A2(_08321_));
 sg13g2_nand2_1 _13798_ (.Y(_08323_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[26] ));
 sg13g2_nand2_1 _13799_ (.Y(_08324_),
    .A(net202),
    .B(net3688));
 sg13g2_o21ai_1 _13800_ (.B1(_08324_),
    .Y(_00660_),
    .A1(net3687),
    .A2(_08323_));
 sg13g2_nand2_1 _13801_ (.Y(_08325_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[27] ));
 sg13g2_nand2_1 _13802_ (.Y(_08326_),
    .A(net108),
    .B(net3688));
 sg13g2_o21ai_1 _13803_ (.B1(_08326_),
    .Y(_00661_),
    .A1(net3687),
    .A2(_08325_));
 sg13g2_nand2_1 _13804_ (.Y(_08327_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[28] ));
 sg13g2_nand2_1 _13805_ (.Y(_08328_),
    .A(net106),
    .B(net3687));
 sg13g2_o21ai_1 _13806_ (.B1(_08328_),
    .Y(_00662_),
    .A1(net3687),
    .A2(_08327_));
 sg13g2_nand2_1 _13807_ (.Y(_08329_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[29] ));
 sg13g2_nand2_1 _13808_ (.Y(_08330_),
    .A(net124),
    .B(net3688));
 sg13g2_o21ai_1 _13809_ (.B1(_08330_),
    .Y(_00663_),
    .A1(net3688),
    .A2(_08329_));
 sg13g2_nand2_1 _13810_ (.Y(_08331_),
    .A(net4781),
    .B(\soc_inst.mem_ctrl.spi_data_out[30] ));
 sg13g2_nand2_1 _13811_ (.Y(_08332_),
    .A(net182),
    .B(net3689));
 sg13g2_o21ai_1 _13812_ (.B1(_08332_),
    .Y(_00664_),
    .A1(net3689),
    .A2(_08331_));
 sg13g2_nand2_1 _13813_ (.Y(_08333_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[31] ));
 sg13g2_nand2_1 _13814_ (.Y(_08334_),
    .A(net282),
    .B(net3687));
 sg13g2_o21ai_1 _13815_ (.B1(_08334_),
    .Y(_00665_),
    .A1(net3688),
    .A2(_08333_));
 sg13g2_nand2_1 _13816_ (.Y(_08335_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[16] ));
 sg13g2_nand2_1 _13817_ (.Y(_08336_),
    .A(net139),
    .B(net3690));
 sg13g2_o21ai_1 _13818_ (.B1(_08336_),
    .Y(_00666_),
    .A1(net3690),
    .A2(_08335_));
 sg13g2_nand2_1 _13819_ (.Y(_08337_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[17] ));
 sg13g2_nand2_1 _13820_ (.Y(_08338_),
    .A(net332),
    .B(net3690));
 sg13g2_o21ai_1 _13821_ (.B1(_08338_),
    .Y(_00667_),
    .A1(net3690),
    .A2(_08337_));
 sg13g2_nand2_1 _13822_ (.Y(_08339_),
    .A(net4776),
    .B(\soc_inst.mem_ctrl.spi_data_out[18] ));
 sg13g2_nand2_1 _13823_ (.Y(_08340_),
    .A(net179),
    .B(net3686));
 sg13g2_o21ai_1 _13824_ (.B1(_08340_),
    .Y(_00668_),
    .A1(net3686),
    .A2(_08339_));
 sg13g2_nand2_1 _13825_ (.Y(_08341_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[19] ));
 sg13g2_nand2_1 _13826_ (.Y(_08342_),
    .A(net200),
    .B(net3690));
 sg13g2_o21ai_1 _13827_ (.B1(_08342_),
    .Y(_00669_),
    .A1(net3690),
    .A2(_08341_));
 sg13g2_nand2_1 _13828_ (.Y(_08343_),
    .A(net4781),
    .B(\soc_inst.mem_ctrl.spi_data_out[20] ));
 sg13g2_nand2_1 _13829_ (.Y(_08344_),
    .A(net228),
    .B(net3691));
 sg13g2_o21ai_1 _13830_ (.B1(_08344_),
    .Y(_00670_),
    .A1(net3691),
    .A2(_08343_));
 sg13g2_nand2_1 _13831_ (.Y(_08345_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[21] ));
 sg13g2_nand2_1 _13832_ (.Y(_08346_),
    .A(net234),
    .B(net3690));
 sg13g2_o21ai_1 _13833_ (.B1(_08346_),
    .Y(_00671_),
    .A1(net3691),
    .A2(_08345_));
 sg13g2_nand2_1 _13834_ (.Y(_08347_),
    .A(net4780),
    .B(\soc_inst.mem_ctrl.spi_data_out[22] ));
 sg13g2_nand2_1 _13835_ (.Y(_08348_),
    .A(net287),
    .B(net3690));
 sg13g2_o21ai_1 _13836_ (.B1(_08348_),
    .Y(_00672_),
    .A1(net3691),
    .A2(_08347_));
 sg13g2_nand2_1 _13837_ (.Y(_08349_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[23] ));
 sg13g2_nand2_1 _13838_ (.Y(_08350_),
    .A(net255),
    .B(net3688));
 sg13g2_o21ai_1 _13839_ (.B1(_08350_),
    .Y(_00673_),
    .A1(net3687),
    .A2(_08349_));
 sg13g2_nand2_1 _13840_ (.Y(_08351_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[8] ));
 sg13g2_nand2_1 _13841_ (.Y(_08352_),
    .A(net204),
    .B(net3684));
 sg13g2_o21ai_1 _13842_ (.B1(_08352_),
    .Y(_00674_),
    .A1(net3684),
    .A2(_08351_));
 sg13g2_nand2_1 _13843_ (.Y(_08353_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[9] ));
 sg13g2_nand2_1 _13844_ (.Y(_08354_),
    .A(net161),
    .B(net3684));
 sg13g2_o21ai_1 _13845_ (.B1(_08354_),
    .Y(_00675_),
    .A1(net3684),
    .A2(_08353_));
 sg13g2_nand2_1 _13846_ (.Y(_08355_),
    .A(net4776),
    .B(\soc_inst.mem_ctrl.spi_data_out[10] ));
 sg13g2_nand2_1 _13847_ (.Y(_08356_),
    .A(net115),
    .B(net3685));
 sg13g2_o21ai_1 _13848_ (.B1(_08356_),
    .Y(_00676_),
    .A1(net3685),
    .A2(_08355_));
 sg13g2_nand2_1 _13849_ (.Y(_08357_),
    .A(net4776),
    .B(\soc_inst.mem_ctrl.spi_data_out[11] ));
 sg13g2_nand2_1 _13850_ (.Y(_08358_),
    .A(net126),
    .B(net3686));
 sg13g2_o21ai_1 _13851_ (.B1(_08358_),
    .Y(_00677_),
    .A1(net3686),
    .A2(_08357_));
 sg13g2_nand2_1 _13852_ (.Y(_08359_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[12] ));
 sg13g2_nand2_1 _13853_ (.Y(_08360_),
    .A(net262),
    .B(net3683));
 sg13g2_o21ai_1 _13854_ (.B1(_08360_),
    .Y(_00678_),
    .A1(net3683),
    .A2(_08359_));
 sg13g2_nand2_1 _13855_ (.Y(_08361_),
    .A(net4776),
    .B(\soc_inst.mem_ctrl.spi_data_out[13] ));
 sg13g2_nand2_1 _13856_ (.Y(_08362_),
    .A(net122),
    .B(net3683));
 sg13g2_o21ai_1 _13857_ (.B1(_08362_),
    .Y(_00679_),
    .A1(net3683),
    .A2(_08361_));
 sg13g2_nand2_1 _13858_ (.Y(_08363_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[14] ));
 sg13g2_nand2_1 _13859_ (.Y(_08364_),
    .A(net251),
    .B(net3683));
 sg13g2_o21ai_1 _13860_ (.B1(_08364_),
    .Y(_00680_),
    .A1(net3683),
    .A2(_08363_));
 sg13g2_nand2_1 _13861_ (.Y(_08365_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[15] ));
 sg13g2_nand2_1 _13862_ (.Y(_08366_),
    .A(net184),
    .B(net3683));
 sg13g2_o21ai_1 _13863_ (.B1(_08366_),
    .Y(_00681_),
    .A1(net3684),
    .A2(_08365_));
 sg13g2_nand2_1 _13864_ (.Y(_08367_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[0] ));
 sg13g2_nand2_1 _13865_ (.Y(_08368_),
    .A(net146),
    .B(net3685));
 sg13g2_o21ai_1 _13866_ (.B1(_08368_),
    .Y(_00682_),
    .A1(net3685),
    .A2(_08367_));
 sg13g2_nand2_1 _13867_ (.Y(_08369_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[1] ));
 sg13g2_nand2_1 _13868_ (.Y(_08370_),
    .A(net298),
    .B(net3692));
 sg13g2_o21ai_1 _13869_ (.B1(_08370_),
    .Y(_00683_),
    .A1(net3692),
    .A2(_08369_));
 sg13g2_nand2_1 _13870_ (.Y(_08371_),
    .A(net4777),
    .B(\soc_inst.mem_ctrl.spi_data_out[2] ));
 sg13g2_nand2_1 _13871_ (.Y(_08372_),
    .A(net230),
    .B(net3687));
 sg13g2_o21ai_1 _13872_ (.B1(_08372_),
    .Y(_00684_),
    .A1(net3687),
    .A2(_08371_));
 sg13g2_nand2_1 _13873_ (.Y(_08373_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[3] ));
 sg13g2_nand2_1 _13874_ (.Y(_08374_),
    .A(net222),
    .B(net3692));
 sg13g2_o21ai_1 _13875_ (.B1(_08374_),
    .Y(_00685_),
    .A1(net3692),
    .A2(_08373_));
 sg13g2_nand2_1 _13876_ (.Y(_08375_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[4] ));
 sg13g2_nand2_1 _13877_ (.Y(_08376_),
    .A(net247),
    .B(net3684));
 sg13g2_o21ai_1 _13878_ (.B1(_08376_),
    .Y(_00686_),
    .A1(net3684),
    .A2(_08375_));
 sg13g2_nand2_1 _13879_ (.Y(_08377_),
    .A(net4778),
    .B(\soc_inst.mem_ctrl.spi_data_out[5] ));
 sg13g2_nand2_1 _13880_ (.Y(_08378_),
    .A(net253),
    .B(net3692));
 sg13g2_o21ai_1 _13881_ (.B1(_08378_),
    .Y(_00687_),
    .A1(net3692),
    .A2(_08377_));
 sg13g2_nand2_1 _13882_ (.Y(_08379_),
    .A(net4776),
    .B(\soc_inst.mem_ctrl.spi_data_out[6] ));
 sg13g2_nand2_1 _13883_ (.Y(_08380_),
    .A(net189),
    .B(net3685));
 sg13g2_o21ai_1 _13884_ (.B1(_08380_),
    .Y(_00688_),
    .A1(net3685),
    .A2(_08379_));
 sg13g2_nand2_1 _13885_ (.Y(_08381_),
    .A(net4775),
    .B(\soc_inst.mem_ctrl.spi_data_out[7] ));
 sg13g2_nand2_1 _13886_ (.Y(_08382_),
    .A(net249),
    .B(net3683));
 sg13g2_o21ai_1 _13887_ (.B1(_08382_),
    .Y(_00689_),
    .A1(net3684),
    .A2(_08381_));
 sg13g2_nor2b_1 _13888_ (.A(_08306_),
    .B_N(_05949_),
    .Y(_08383_));
 sg13g2_o21ai_1 _13889_ (.B1(net2939),
    .Y(_08384_),
    .A1(net5075),
    .A2(net4779));
 sg13g2_o21ai_1 _13890_ (.B1(_08384_),
    .Y(_08385_),
    .A1(_05868_),
    .A2(_08308_));
 sg13g2_mux2_1 _13891_ (.A0(net2968),
    .A1(_08385_),
    .S(_08383_),
    .X(_00690_));
 sg13g2_and3_2 _13892_ (.X(_08386_),
    .A(_06038_),
    .B(_06040_),
    .C(_06151_));
 sg13g2_nand3_1 _13893_ (.B(_06040_),
    .C(_06151_),
    .A(_06038_),
    .Y(_08387_));
 sg13g2_nor2_1 _13894_ (.A(net2491),
    .B(net4219),
    .Y(_08388_));
 sg13g2_nand2_2 _13895_ (.Y(_08389_),
    .A(net5059),
    .B(_06151_));
 sg13g2_nor4_1 _13896_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .B(net4784),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .D(_08389_),
    .Y(_08390_));
 sg13g2_nor2_1 _13897_ (.A(net2543),
    .B(net4218),
    .Y(_08391_));
 sg13g2_a21oi_1 _13898_ (.A1(net2491),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ),
    .Y(_08392_),
    .B1(net4219));
 sg13g2_o21ai_1 _13899_ (.B1(_06149_),
    .Y(_08393_),
    .A1(_08390_),
    .A2(_08392_));
 sg13g2_nor2_2 _13900_ (.A(net2215),
    .B(net504),
    .Y(_08394_));
 sg13g2_or2_1 _13901_ (.X(_08395_),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ));
 sg13g2_nand3_1 _13902_ (.B(net5073),
    .C(_08394_),
    .A(_05495_),
    .Y(_08396_));
 sg13g2_o21ai_1 _13903_ (.B1(net5066),
    .Y(_08397_),
    .A1(net5081),
    .A2(\soc_inst.bus_spi_sclk ));
 sg13g2_a21oi_2 _13904_ (.B1(net5073),
    .Y(_08398_),
    .A2(net408),
    .A1(net2740));
 sg13g2_inv_1 _13905_ (.Y(_08399_),
    .A(_08398_));
 sg13g2_nand4_1 _13906_ (.B(_08396_),
    .C(_08397_),
    .A(_08393_),
    .Y(_08400_),
    .D(_08399_));
 sg13g2_nor2_1 _13907_ (.A(_05495_),
    .B(_08400_),
    .Y(_08401_));
 sg13g2_a22oi_1 _13908_ (.Y(_08402_),
    .B1(net3971),
    .B2(net9),
    .A2(net4036),
    .A1(net1927));
 sg13g2_inv_1 _13909_ (.Y(_00691_),
    .A(_08402_));
 sg13g2_a22oi_1 _13910_ (.Y(_08403_),
    .B1(net3974),
    .B2(net10),
    .A2(net4039),
    .A1(net1954));
 sg13g2_inv_1 _13911_ (.Y(_00692_),
    .A(_08403_));
 sg13g2_a22oi_1 _13912_ (.Y(_08404_),
    .B1(net3974),
    .B2(net11),
    .A2(net4039),
    .A1(net1750));
 sg13g2_inv_1 _13913_ (.Y(_00693_),
    .A(_08404_));
 sg13g2_a22oi_1 _13914_ (.Y(_08405_),
    .B1(net3972),
    .B2(net12),
    .A2(net4037),
    .A1(net1848));
 sg13g2_inv_1 _13915_ (.Y(_00694_),
    .A(_08405_));
 sg13g2_a22oi_1 _13916_ (.Y(_08406_),
    .B1(net3971),
    .B2(net1927),
    .A2(net4036),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ));
 sg13g2_inv_1 _13917_ (.Y(_00695_),
    .A(net1928));
 sg13g2_a22oi_1 _13918_ (.Y(_08407_),
    .B1(net3974),
    .B2(net1954),
    .A2(net4039),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ));
 sg13g2_inv_1 _13919_ (.Y(_00696_),
    .A(net1955));
 sg13g2_a22oi_1 _13920_ (.Y(_08408_),
    .B1(net3973),
    .B2(net1750),
    .A2(net4038),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ));
 sg13g2_inv_1 _13921_ (.Y(_00697_),
    .A(net1751));
 sg13g2_a22oi_1 _13922_ (.Y(_08409_),
    .B1(net3972),
    .B2(net1848),
    .A2(net4037),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ));
 sg13g2_inv_1 _13923_ (.Y(_00698_),
    .A(net1849));
 sg13g2_a22oi_1 _13924_ (.Y(_08410_),
    .B1(net3971),
    .B2(net2491),
    .A2(net4036),
    .A1(net1913));
 sg13g2_inv_1 _13925_ (.Y(_00699_),
    .A(_08410_));
 sg13g2_a22oi_1 _13926_ (.Y(_08411_),
    .B1(net3973),
    .B2(net2543),
    .A2(net4038),
    .A1(net1836));
 sg13g2_inv_1 _13927_ (.Y(_00700_),
    .A(_08411_));
 sg13g2_a22oi_1 _13928_ (.Y(_08412_),
    .B1(net3975),
    .B2(net1929),
    .A2(net4040),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ));
 sg13g2_inv_1 _13929_ (.Y(_00701_),
    .A(net1930));
 sg13g2_a22oi_1 _13930_ (.Y(_08413_),
    .B1(net3972),
    .B2(net1967),
    .A2(net4037),
    .A1(net1865));
 sg13g2_inv_1 _13931_ (.Y(_00702_),
    .A(_08413_));
 sg13g2_a22oi_1 _13932_ (.Y(_08414_),
    .B1(net3971),
    .B2(net1913),
    .A2(net4036),
    .A1(net1399));
 sg13g2_inv_1 _13933_ (.Y(_00703_),
    .A(_08414_));
 sg13g2_a22oi_1 _13934_ (.Y(_08415_),
    .B1(net3973),
    .B2(net1836),
    .A2(net4038),
    .A1(net1096));
 sg13g2_inv_1 _13935_ (.Y(_00704_),
    .A(_08415_));
 sg13g2_a22oi_1 _13936_ (.Y(_08416_),
    .B1(net3975),
    .B2(net2005),
    .A2(net4040),
    .A1(net1499));
 sg13g2_inv_1 _13937_ (.Y(_00705_),
    .A(_08416_));
 sg13g2_a22oi_1 _13938_ (.Y(_08417_),
    .B1(net3972),
    .B2(net1865),
    .A2(net4037),
    .A1(net1388));
 sg13g2_inv_1 _13939_ (.Y(_00706_),
    .A(_08417_));
 sg13g2_a22oi_1 _13940_ (.Y(_08418_),
    .B1(net3971),
    .B2(net1399),
    .A2(net4036),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ));
 sg13g2_inv_1 _13941_ (.Y(_00707_),
    .A(net1400));
 sg13g2_a22oi_1 _13942_ (.Y(_08419_),
    .B1(net3974),
    .B2(net1096),
    .A2(net4039),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ));
 sg13g2_inv_1 _13943_ (.Y(_00708_),
    .A(net1097));
 sg13g2_a22oi_1 _13944_ (.Y(_08420_),
    .B1(net3973),
    .B2(net1499),
    .A2(net4038),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ));
 sg13g2_inv_1 _13945_ (.Y(_00709_),
    .A(net1500));
 sg13g2_a22oi_1 _13946_ (.Y(_08421_),
    .B1(net3972),
    .B2(net1388),
    .A2(net4037),
    .A1(net1341));
 sg13g2_inv_1 _13947_ (.Y(_00710_),
    .A(_08421_));
 sg13g2_a22oi_1 _13948_ (.Y(_08422_),
    .B1(net3971),
    .B2(net1719),
    .A2(net4036),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ));
 sg13g2_inv_1 _13949_ (.Y(_00711_),
    .A(net1720));
 sg13g2_a22oi_1 _13950_ (.Y(_08423_),
    .B1(net3974),
    .B2(net1859),
    .A2(net4039),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ));
 sg13g2_inv_1 _13951_ (.Y(_00712_),
    .A(net1860));
 sg13g2_a22oi_1 _13952_ (.Y(_08424_),
    .B1(net3973),
    .B2(net1600),
    .A2(net4038),
    .A1(net1514));
 sg13g2_inv_1 _13953_ (.Y(_00713_),
    .A(_08424_));
 sg13g2_a22oi_1 _13954_ (.Y(_08425_),
    .B1(net3972),
    .B2(net1341),
    .A2(net4037),
    .A1(net953));
 sg13g2_inv_1 _13955_ (.Y(_00714_),
    .A(_08425_));
 sg13g2_a22oi_1 _13956_ (.Y(_08426_),
    .B1(net3971),
    .B2(net1846),
    .A2(net4036),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ));
 sg13g2_inv_1 _13957_ (.Y(_00715_),
    .A(net1847));
 sg13g2_a22oi_1 _13958_ (.Y(_08427_),
    .B1(net3974),
    .B2(net2040),
    .A2(net4038),
    .A1(net1723));
 sg13g2_inv_1 _13959_ (.Y(_00716_),
    .A(_08427_));
 sg13g2_a22oi_1 _13960_ (.Y(_08428_),
    .B1(net3973),
    .B2(net1514),
    .A2(net4039),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ));
 sg13g2_inv_1 _13961_ (.Y(_00717_),
    .A(net1515));
 sg13g2_a22oi_1 _13962_ (.Y(_08429_),
    .B1(net3975),
    .B2(net953),
    .A2(net4040),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ));
 sg13g2_inv_1 _13963_ (.Y(_00718_),
    .A(net954));
 sg13g2_a22oi_1 _13964_ (.Y(_08430_),
    .B1(net3971),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ),
    .A2(net4036),
    .A1(net866));
 sg13g2_inv_1 _13965_ (.Y(_00719_),
    .A(net867));
 sg13g2_a22oi_1 _13966_ (.Y(_08431_),
    .B1(net3973),
    .B2(net1723),
    .A2(net4038),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ));
 sg13g2_inv_1 _13967_ (.Y(_00720_),
    .A(net1724));
 sg13g2_a22oi_1 _13968_ (.Y(_08432_),
    .B1(net3973),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ),
    .A2(net4038),
    .A1(net1046));
 sg13g2_inv_1 _13969_ (.Y(_00721_),
    .A(net1047));
 sg13g2_a22oi_1 _13970_ (.Y(_08433_),
    .B1(net3975),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ),
    .A2(net4040),
    .A1(net970));
 sg13g2_inv_1 _13971_ (.Y(_00722_),
    .A(net971));
 sg13g2_a21oi_1 _13972_ (.A1(net2203),
    .A2(_08394_),
    .Y(_08434_),
    .B1(_08398_));
 sg13g2_nor2_1 _13973_ (.A(net5081),
    .B(_08434_),
    .Y(_08435_));
 sg13g2_a21oi_1 _13974_ (.A1(_05417_),
    .A2(_08434_),
    .Y(_00723_),
    .B1(_08435_));
 sg13g2_nor2_1 _13975_ (.A(net5061),
    .B(net486),
    .Y(_08436_));
 sg13g2_nor3_1 _13976_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .Y(_08437_));
 sg13g2_nor2b_2 _13977_ (.A(net504),
    .B_N(_08437_),
    .Y(_08438_));
 sg13g2_nand3_1 _13978_ (.B(_08436_),
    .C(_08438_),
    .A(net5073),
    .Y(_08439_));
 sg13g2_or2_1 _13979_ (.X(_08440_),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .A(net5072));
 sg13g2_nor3_1 _13980_ (.A(net5066),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .C(_08440_),
    .Y(_08441_));
 sg13g2_nor2_1 _13981_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .B(net5064),
    .Y(_08442_));
 sg13g2_nand2_1 _13982_ (.Y(_08443_),
    .A(_08441_),
    .B(_08442_));
 sg13g2_nor3_1 _13983_ (.A(net496),
    .B(_08439_),
    .C(_08443_),
    .Y(_08444_));
 sg13g2_o21ai_1 _13984_ (.B1(_06141_),
    .Y(_08445_),
    .A1(_05501_),
    .A2(_06042_));
 sg13g2_nand2_1 _13985_ (.Y(_08446_),
    .A(_08437_),
    .B(_08442_));
 sg13g2_nand4_1 _13986_ (.B(_06048_),
    .C(_08394_),
    .A(_05496_),
    .Y(_08447_),
    .D(_08441_));
 sg13g2_nor2_1 _13987_ (.A(_08446_),
    .B(_08447_),
    .Y(_08448_));
 sg13g2_a21oi_1 _13988_ (.A1(net496),
    .A2(_08445_),
    .Y(_08449_),
    .B1(_08448_));
 sg13g2_nor4_1 _13989_ (.A(net5061),
    .B(net5121),
    .C(net486),
    .D(_08444_),
    .Y(_08450_));
 sg13g2_nor2b_1 _13990_ (.A(net5121),
    .B_N(_08444_),
    .Y(_08451_));
 sg13g2_a22oi_1 _13991_ (.Y(_08452_),
    .B1(_08451_),
    .B2(net2732),
    .A2(_08450_),
    .A1(_08449_));
 sg13g2_inv_1 _13992_ (.Y(_00724_),
    .A(net2733));
 sg13g2_nand3_1 _13993_ (.B(_05495_),
    .C(net5073),
    .A(net2735),
    .Y(_08453_));
 sg13g2_nor3_1 _13994_ (.A(net5081),
    .B(net97),
    .C(_08393_),
    .Y(_08454_));
 sg13g2_nor2_1 _13995_ (.A(net5061),
    .B(_08454_),
    .Y(_08455_));
 sg13g2_nand2_1 _13996_ (.Y(_00725_),
    .A(_08453_),
    .B(_08455_));
 sg13g2_nor2_1 _13997_ (.A(_08439_),
    .B(_08445_),
    .Y(_08456_));
 sg13g2_nor2_1 _13998_ (.A(_08443_),
    .B(_08456_),
    .Y(_08457_));
 sg13g2_nor3_1 _13999_ (.A(net5122),
    .B(_08444_),
    .C(_08457_),
    .Y(_08458_));
 sg13g2_a21o_1 _14000_ (.A2(_08451_),
    .A1(net627),
    .B1(_08458_),
    .X(_00726_));
 sg13g2_nor3_1 _14001_ (.A(net496),
    .B(net5065),
    .C(_08443_),
    .Y(_08459_));
 sg13g2_nand3_1 _14002_ (.B(_08438_),
    .C(_08459_),
    .A(net5073),
    .Y(_08460_));
 sg13g2_nand2_1 _14003_ (.Y(_08461_),
    .A(_06048_),
    .B(_08459_));
 sg13g2_o21ai_1 _14004_ (.B1(_08461_),
    .Y(_08462_),
    .A1(_05501_),
    .A2(_08459_));
 sg13g2_and4_1 _14005_ (.A(_07068_),
    .B(_08438_),
    .C(_08460_),
    .D(_08462_),
    .X(_08463_));
 sg13g2_a21oi_1 _14006_ (.A1(_07068_),
    .A2(_08460_),
    .Y(_08464_),
    .B1(net5077));
 sg13g2_nor2_1 _14007_ (.A(_08463_),
    .B(_08464_),
    .Y(_00727_));
 sg13g2_a21oi_1 _14008_ (.A1(_06665_),
    .A2(net4177),
    .Y(_08465_),
    .B1(_06722_));
 sg13g2_nor2b_1 _14009_ (.A(_06719_),
    .B_N(_08465_),
    .Y(_08466_));
 sg13g2_a21oi_1 _14010_ (.A1(_07609_),
    .A2(net3760),
    .Y(_08467_),
    .B1(net167));
 sg13g2_a21oi_1 _14011_ (.A1(_05415_),
    .A2(_07609_),
    .Y(_08468_),
    .B1(_07605_));
 sg13g2_and2_1 _14012_ (.A(net4698),
    .B(net3757),
    .X(_08469_));
 sg13g2_nand2_2 _14013_ (.Y(_08470_),
    .A(net4698),
    .B(net3758));
 sg13g2_a21oi_1 _14014_ (.A1(_08468_),
    .A2(net3749),
    .Y(_00728_),
    .B1(net168));
 sg13g2_a21oi_1 _14015_ (.A1(_07614_),
    .A2(net3760),
    .Y(_08471_),
    .B1(net163));
 sg13g2_a21oi_1 _14016_ (.A1(net4757),
    .A2(_07614_),
    .Y(_08472_),
    .B1(_07612_));
 sg13g2_a21oi_1 _14017_ (.A1(net3749),
    .A2(_08472_),
    .Y(_00729_),
    .B1(net164));
 sg13g2_nor2b_2 _14018_ (.A(net4869),
    .B_N(net457),
    .Y(_08473_));
 sg13g2_inv_1 _14019_ (.Y(_08474_),
    .A(_08473_));
 sg13g2_a21oi_1 _14020_ (.A1(net3760),
    .A2(_08473_),
    .Y(_08475_),
    .B1(net111));
 sg13g2_o21ai_1 _14021_ (.B1(net4612),
    .Y(_08476_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .A2(net4609));
 sg13g2_a21oi_1 _14022_ (.A1(net4755),
    .A2(_08473_),
    .Y(_08477_),
    .B1(_08476_));
 sg13g2_a21oi_1 _14023_ (.A1(net3749),
    .A2(_08477_),
    .Y(_00730_),
    .B1(net112));
 sg13g2_a21oi_1 _14024_ (.A1(_07618_),
    .A2(net3761),
    .Y(_08478_),
    .B1(net135));
 sg13g2_a21oi_1 _14025_ (.A1(net4755),
    .A2(_07618_),
    .Y(_08479_),
    .B1(_07616_));
 sg13g2_a21oi_1 _14026_ (.A1(net3749),
    .A2(_08479_),
    .Y(_00731_),
    .B1(net136));
 sg13g2_a21oi_1 _14027_ (.A1(_07622_),
    .A2(net3760),
    .Y(_08480_),
    .B1(net154));
 sg13g2_a21oi_1 _14028_ (.A1(net4755),
    .A2(_07622_),
    .Y(_08481_),
    .B1(_07620_));
 sg13g2_a21oi_1 _14029_ (.A1(net3749),
    .A2(_08481_),
    .Y(_00732_),
    .B1(net155));
 sg13g2_a21oi_1 _14030_ (.A1(_07626_),
    .A2(net3761),
    .Y(_08482_),
    .B1(net141));
 sg13g2_a21oi_1 _14031_ (.A1(net4756),
    .A2(_07626_),
    .Y(_08483_),
    .B1(_07624_));
 sg13g2_a21oi_1 _14032_ (.A1(net3750),
    .A2(_08483_),
    .Y(_00733_),
    .B1(net142));
 sg13g2_nor2b_2 _14033_ (.A(net4869),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .Y(_08484_));
 sg13g2_inv_1 _14034_ (.Y(_08485_),
    .A(_08484_));
 sg13g2_a21oi_1 _14035_ (.A1(net3760),
    .A2(_08484_),
    .Y(_08486_),
    .B1(net236));
 sg13g2_o21ai_1 _14036_ (.B1(net4613),
    .Y(_08487_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .A2(net4609));
 sg13g2_a21oi_1 _14037_ (.A1(net4755),
    .A2(_08484_),
    .Y(_08488_),
    .B1(_08487_));
 sg13g2_a21oi_1 _14038_ (.A1(net3749),
    .A2(_08488_),
    .Y(_00734_),
    .B1(net237));
 sg13g2_nor2b_2 _14039_ (.A(net4867),
    .B_N(net2979),
    .Y(_08489_));
 sg13g2_a21oi_1 _14040_ (.A1(net3758),
    .A2(_08489_),
    .Y(_08490_),
    .B1(net209));
 sg13g2_o21ai_1 _14041_ (.B1(net4614),
    .Y(_08491_),
    .A1(net2979),
    .A2(net4610));
 sg13g2_a21oi_1 _14042_ (.A1(net4755),
    .A2(_08489_),
    .Y(_08492_),
    .B1(_08491_));
 sg13g2_a21oi_1 _14043_ (.A1(net3749),
    .A2(_08492_),
    .Y(_00735_),
    .B1(net210));
 sg13g2_nor2b_1 _14044_ (.A(net4866),
    .B_N(net928),
    .Y(_08493_));
 sg13g2_a21oi_1 _14045_ (.A1(net3757),
    .A2(_08493_),
    .Y(_08494_),
    .B1(net219));
 sg13g2_o21ai_1 _14046_ (.B1(net4615),
    .Y(_08495_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .A2(net4609));
 sg13g2_a21oi_1 _14047_ (.A1(net928),
    .A2(net4709),
    .Y(_08496_),
    .B1(_08495_));
 sg13g2_a21oi_1 _14048_ (.A1(net3750),
    .A2(_08496_),
    .Y(_00736_),
    .B1(net220));
 sg13g2_nor2b_1 _14049_ (.A(net4867),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .Y(_08497_));
 sg13g2_a21oi_1 _14050_ (.A1(net3761),
    .A2(_08497_),
    .Y(_08498_),
    .B1(net175));
 sg13g2_o21ai_1 _14051_ (.B1(net4614),
    .Y(_08499_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .A2(net4610));
 sg13g2_a21oi_1 _14052_ (.A1(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .A2(net4709),
    .Y(_08500_),
    .B1(_08499_));
 sg13g2_a21oi_1 _14053_ (.A1(net3749),
    .A2(_08500_),
    .Y(_00737_),
    .B1(net176));
 sg13g2_nor2b_1 _14054_ (.A(net4866),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .Y(_08501_));
 sg13g2_a21oi_1 _14055_ (.A1(net3757),
    .A2(_08501_),
    .Y(_08502_),
    .B1(net132));
 sg13g2_o21ai_1 _14056_ (.B1(net4612),
    .Y(_08503_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .A2(net4608));
 sg13g2_a21oi_1 _14057_ (.A1(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .A2(net4709),
    .Y(_08504_),
    .B1(_08503_));
 sg13g2_a21oi_1 _14058_ (.A1(net3748),
    .A2(_08504_),
    .Y(_00738_),
    .B1(net133));
 sg13g2_nor2b_1 _14059_ (.A(net4867),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .Y(_08505_));
 sg13g2_a21oi_1 _14060_ (.A1(net3758),
    .A2(_08505_),
    .Y(_08506_),
    .B1(net206));
 sg13g2_o21ai_1 _14061_ (.B1(net4613),
    .Y(_08507_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .A2(net4606));
 sg13g2_a21oi_1 _14062_ (.A1(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .A2(net4708),
    .Y(_08508_),
    .B1(_08507_));
 sg13g2_a21oi_1 _14063_ (.A1(net3748),
    .A2(_08508_),
    .Y(_00739_),
    .B1(net207));
 sg13g2_nor2b_1 _14064_ (.A(net4867),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .Y(_08509_));
 sg13g2_a21oi_1 _14065_ (.A1(net3758),
    .A2(_08509_),
    .Y(_08510_),
    .B1(net259));
 sg13g2_o21ai_1 _14066_ (.B1(net4613),
    .Y(_08511_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .A2(net4605));
 sg13g2_a21oi_1 _14067_ (.A1(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .A2(net4708),
    .Y(_08512_),
    .B1(_08511_));
 sg13g2_a21oi_1 _14068_ (.A1(net3748),
    .A2(_08512_),
    .Y(_00740_),
    .B1(net260));
 sg13g2_nor2b_1 _14069_ (.A(net4866),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .Y(_08513_));
 sg13g2_a21oi_1 _14070_ (.A1(net3757),
    .A2(_08513_),
    .Y(_08514_),
    .B1(net193));
 sg13g2_o21ai_1 _14071_ (.B1(net4612),
    .Y(_08515_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .A2(net4603));
 sg13g2_a21oi_1 _14072_ (.A1(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .A2(net4708),
    .Y(_08516_),
    .B1(_08515_));
 sg13g2_a21oi_1 _14073_ (.A1(net3748),
    .A2(_08516_),
    .Y(_00741_),
    .B1(net194));
 sg13g2_nor2b_2 _14074_ (.A(net4866),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .Y(_08517_));
 sg13g2_a21oi_1 _14075_ (.A1(net3757),
    .A2(_08517_),
    .Y(_08518_),
    .B1(net172));
 sg13g2_o21ai_1 _14076_ (.B1(net4612),
    .Y(_08519_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .A2(net4603));
 sg13g2_a21oi_1 _14077_ (.A1(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .A2(net4708),
    .Y(_08520_),
    .B1(_08519_));
 sg13g2_a21oi_1 _14078_ (.A1(net3748),
    .A2(_08520_),
    .Y(_00742_),
    .B1(net173));
 sg13g2_nor2b_1 _14079_ (.A(net4867),
    .B_N(net1576),
    .Y(_08521_));
 sg13g2_a21oi_1 _14080_ (.A1(net3758),
    .A2(_08521_),
    .Y(_08522_),
    .B1(net284));
 sg13g2_o21ai_1 _14081_ (.B1(net4612),
    .Y(_08523_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .A2(net4604));
 sg13g2_a21oi_1 _14082_ (.A1(net1576),
    .A2(net4708),
    .Y(_08524_),
    .B1(_08523_));
 sg13g2_a21oi_1 _14083_ (.A1(net3750),
    .A2(_08524_),
    .Y(_00743_),
    .B1(net285));
 sg13g2_nor2b_1 _14084_ (.A(net4866),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .Y(_08525_));
 sg13g2_a21oi_1 _14085_ (.A1(net3757),
    .A2(_08525_),
    .Y(_08526_),
    .B1(net129));
 sg13g2_o21ai_1 _14086_ (.B1(net4612),
    .Y(_08527_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .A2(net4603));
 sg13g2_a21oi_1 _14087_ (.A1(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .A2(net4708),
    .Y(_08528_),
    .B1(_08527_));
 sg13g2_a21oi_1 _14088_ (.A1(net3748),
    .A2(_08528_),
    .Y(_00744_),
    .B1(net130));
 sg13g2_nor2b_1 _14089_ (.A(net4867),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .Y(_08529_));
 sg13g2_a21oi_1 _14090_ (.A1(net3757),
    .A2(_08529_),
    .Y(_08530_),
    .B1(net291));
 sg13g2_o21ai_1 _14091_ (.B1(net4612),
    .Y(_08531_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .A2(net4604));
 sg13g2_a21oi_1 _14092_ (.A1(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .A2(net4708),
    .Y(_08532_),
    .B1(_08531_));
 sg13g2_a21oi_1 _14093_ (.A1(net3748),
    .A2(_08532_),
    .Y(_00745_),
    .B1(net292));
 sg13g2_nor2b_1 _14094_ (.A(net4866),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .Y(_08533_));
 sg13g2_a21oi_1 _14095_ (.A1(net3757),
    .A2(_08533_),
    .Y(_08534_),
    .B1(net151));
 sg13g2_o21ai_1 _14096_ (.B1(net4612),
    .Y(_08535_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .A2(net4603));
 sg13g2_a21oi_1 _14097_ (.A1(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .A2(net4708),
    .Y(_08536_),
    .B1(_08535_));
 sg13g2_a21oi_1 _14098_ (.A1(net3748),
    .A2(_08536_),
    .Y(_00746_),
    .B1(net152));
 sg13g2_nor2_2 _14099_ (.A(_06673_),
    .B(net4709),
    .Y(_08537_));
 sg13g2_a21oi_2 _14100_ (.B1(net4874),
    .Y(_08538_),
    .A2(net4867),
    .A1(net4877));
 sg13g2_a22oi_1 _14101_ (.Y(_08539_),
    .B1(_08537_),
    .B2(net1344),
    .A2(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .A1(net4754));
 sg13g2_o21ai_1 _14102_ (.B1(net4614),
    .Y(_08540_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .A2(net4607));
 sg13g2_nor2_1 _14103_ (.A(_08538_),
    .B(_08540_),
    .Y(_08541_));
 sg13g2_nor3_1 _14104_ (.A(net3747),
    .B(_08539_),
    .C(_08541_),
    .Y(_08542_));
 sg13g2_a21o_1 _14105_ (.A2(net3747),
    .A1(net1344),
    .B1(_08542_),
    .X(_00747_));
 sg13g2_a22oi_1 _14106_ (.Y(_08543_),
    .B1(_08537_),
    .B2(net1674),
    .A2(net1005),
    .A1(net4754));
 sg13g2_o21ai_1 _14107_ (.B1(net4613),
    .Y(_08544_),
    .A1(net1005),
    .A2(net4605));
 sg13g2_nor2_1 _14108_ (.A(_08538_),
    .B(_08544_),
    .Y(_08545_));
 sg13g2_nor3_1 _14109_ (.A(net3746),
    .B(_08543_),
    .C(_08545_),
    .Y(_08546_));
 sg13g2_a21o_1 _14110_ (.A2(net3746),
    .A1(net1674),
    .B1(_08546_),
    .X(_00748_));
 sg13g2_a22oi_1 _14111_ (.Y(_08547_),
    .B1(_08537_),
    .B2(net1468),
    .A2(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .A1(net4754));
 sg13g2_o21ai_1 _14112_ (.B1(net4614),
    .Y(_08548_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .A2(net4611));
 sg13g2_nor2_1 _14113_ (.A(_08538_),
    .B(_08548_),
    .Y(_08549_));
 sg13g2_nor3_1 _14114_ (.A(net3747),
    .B(_08547_),
    .C(_08549_),
    .Y(_08550_));
 sg13g2_a21o_1 _14115_ (.A2(net3747),
    .A1(net1468),
    .B1(_08550_),
    .X(_00749_));
 sg13g2_a22oi_1 _14116_ (.Y(_08551_),
    .B1(_08537_),
    .B2(net1705),
    .A2(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .A1(net4754));
 sg13g2_o21ai_1 _14117_ (.B1(net4613),
    .Y(_08552_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .A2(net4606));
 sg13g2_nor2_1 _14118_ (.A(_08538_),
    .B(_08552_),
    .Y(_08553_));
 sg13g2_nor3_1 _14119_ (.A(net3746),
    .B(_08551_),
    .C(_08553_),
    .Y(_08554_));
 sg13g2_a21o_1 _14120_ (.A2(net3746),
    .A1(net1705),
    .B1(_08554_),
    .X(_00750_));
 sg13g2_a22oi_1 _14121_ (.Y(_08555_),
    .B1(_08537_),
    .B2(net1572),
    .A2(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .A1(net4754));
 sg13g2_o21ai_1 _14122_ (.B1(net4613),
    .Y(_08556_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .A2(net4606));
 sg13g2_nor2_1 _14123_ (.A(_08538_),
    .B(_08556_),
    .Y(_08557_));
 sg13g2_nor3_1 _14124_ (.A(net3746),
    .B(_08555_),
    .C(_08557_),
    .Y(_08558_));
 sg13g2_a21o_1 _14125_ (.A2(net3746),
    .A1(net1572),
    .B1(_08558_),
    .X(_00751_));
 sg13g2_a22oi_1 _14126_ (.Y(_08559_),
    .B1(_08537_),
    .B2(net1382),
    .A2(net1095),
    .A1(net4754));
 sg13g2_o21ai_1 _14127_ (.B1(net4613),
    .Y(_08560_),
    .A1(net1095),
    .A2(net4605));
 sg13g2_nor2_1 _14128_ (.A(_08538_),
    .B(_08560_),
    .Y(_08561_));
 sg13g2_nor3_1 _14129_ (.A(net3746),
    .B(_08559_),
    .C(_08561_),
    .Y(_08562_));
 sg13g2_a21o_1 _14130_ (.A2(net3746),
    .A1(net1382),
    .B1(_08562_),
    .X(_00752_));
 sg13g2_a22oi_1 _14131_ (.Y(_08563_),
    .B1(_08537_),
    .B2(net1258),
    .A2(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .A1(_05416_));
 sg13g2_o21ai_1 _14132_ (.B1(net4613),
    .Y(_08564_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .A2(net4607));
 sg13g2_nor2_1 _14133_ (.A(_08538_),
    .B(_08564_),
    .Y(_08565_));
 sg13g2_nor3_1 _14134_ (.A(net3747),
    .B(_08563_),
    .C(_08565_),
    .Y(_08566_));
 sg13g2_a21o_1 _14135_ (.A2(net3747),
    .A1(net1258),
    .B1(_08566_),
    .X(_00753_));
 sg13g2_a22oi_1 _14136_ (.Y(_08567_),
    .B1(_08537_),
    .B2(net1332),
    .A2(net4879),
    .A1(_05416_));
 sg13g2_o21ai_1 _14137_ (.B1(net4614),
    .Y(_08568_),
    .A1(net4879),
    .A2(net4607));
 sg13g2_nor2_1 _14138_ (.A(_08538_),
    .B(_08568_),
    .Y(_08569_));
 sg13g2_nor3_1 _14139_ (.A(net3747),
    .B(_08567_),
    .C(_08569_),
    .Y(_08570_));
 sg13g2_a21o_1 _14140_ (.A2(net3747),
    .A1(net1332),
    .B1(_08570_),
    .X(_00754_));
 sg13g2_nand2_1 _14141_ (.Y(_08571_),
    .A(_05501_),
    .B(net5065));
 sg13g2_or2_1 _14142_ (.X(_08572_),
    .B(net5065),
    .A(net5066));
 sg13g2_nor3_1 _14143_ (.A(net5061),
    .B(net474),
    .C(_08572_),
    .Y(_08573_));
 sg13g2_nand4_1 _14144_ (.B(net5073),
    .C(_08438_),
    .A(_05500_),
    .Y(_08574_),
    .D(_08573_));
 sg13g2_a21oi_1 _14145_ (.A1(_08571_),
    .A2(_08574_),
    .Y(_08575_),
    .B1(net2858));
 sg13g2_nand4_1 _14146_ (.B(net2980),
    .C(_06038_),
    .A(_05492_),
    .Y(_08576_),
    .D(_06041_));
 sg13g2_a22oi_1 _14147_ (.Y(_08577_),
    .B1(_05501_),
    .B2(net5065),
    .A2(net5081),
    .A1(net5066));
 sg13g2_nand4_1 _14148_ (.B(_08438_),
    .C(_08576_),
    .A(_05500_),
    .Y(_08578_),
    .D(_08577_));
 sg13g2_a21oi_1 _14149_ (.A1(_08399_),
    .A2(_08573_),
    .Y(_08579_),
    .B1(_08578_));
 sg13g2_nor3_1 _14150_ (.A(net5121),
    .B(net2859),
    .C(_08579_),
    .Y(_00755_));
 sg13g2_nor3_1 _14151_ (.A(net5064),
    .B(_08396_),
    .C(_08440_),
    .Y(_08580_));
 sg13g2_nor2_2 _14152_ (.A(_05495_),
    .B(net5081),
    .Y(_08581_));
 sg13g2_nor2b_1 _14153_ (.A(net5078),
    .B_N(net5072),
    .Y(_08582_));
 sg13g2_or4_1 _14154_ (.A(_08398_),
    .B(_08580_),
    .C(_08581_),
    .D(_08582_),
    .X(_08583_));
 sg13g2_nor2_2 _14155_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .Y(_08584_));
 sg13g2_nor4_2 _14156_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .C(_08395_),
    .Y(_08585_),
    .D(_08440_));
 sg13g2_or4_1 _14157_ (.A(net5066),
    .B(net5064),
    .C(_08395_),
    .D(_08440_),
    .X(_08586_));
 sg13g2_nor2_1 _14158_ (.A(net4280),
    .B(_08586_),
    .Y(_08587_));
 sg13g2_or2_1 _14159_ (.X(_08588_),
    .B(net4152),
    .A(net4159));
 sg13g2_and2_1 _14160_ (.A(net5081),
    .B(_06130_),
    .X(_08589_));
 sg13g2_nand2_2 _14161_ (.Y(_08590_),
    .A(_08394_),
    .B(_08586_));
 sg13g2_a22oi_1 _14162_ (.Y(_08591_),
    .B1(_08590_),
    .B2(net1907),
    .A2(net4149),
    .A1(net696));
 sg13g2_nand2_2 _14163_ (.Y(_08592_),
    .A(_06282_),
    .B(_08584_));
 sg13g2_a21oi_2 _14164_ (.B1(net5080),
    .Y(_08593_),
    .A2(_08584_),
    .A1(_06282_));
 sg13g2_or2_1 _14165_ (.X(_08594_),
    .B(net4144),
    .A(net4159));
 sg13g2_nand2_1 _14166_ (.Y(_08595_),
    .A(net2250),
    .B(net4144));
 sg13g2_a21oi_1 _14167_ (.A1(_08591_),
    .A2(_08595_),
    .Y(_08596_),
    .B1(_08588_));
 sg13g2_a21o_1 _14168_ (.A2(net4159),
    .A1(net2250),
    .B1(_08596_),
    .X(_00756_));
 sg13g2_o21ai_1 _14169_ (.B1(_08394_),
    .Y(_08597_),
    .A1(net4278),
    .A2(_08586_));
 sg13g2_nand2_1 _14170_ (.Y(_08598_),
    .A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .B(net4142));
 sg13g2_a22oi_1 _14171_ (.Y(_08599_),
    .B1(net465),
    .B2(net4149),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .A1(net5069));
 sg13g2_a21oi_1 _14172_ (.A1(_08598_),
    .A2(_08599_),
    .Y(_08600_),
    .B1(net4159));
 sg13g2_a21o_1 _14173_ (.A2(_08594_),
    .A1(net1905),
    .B1(_08600_),
    .X(_00757_));
 sg13g2_nand2_1 _14174_ (.Y(_08601_),
    .A(net389),
    .B(net4149));
 sg13g2_a22oi_1 _14175_ (.Y(_08602_),
    .B1(net4143),
    .B2(\soc_inst.mem_ctrl.spi_addr[2] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ),
    .A1(net5067));
 sg13g2_a21oi_1 _14176_ (.A1(_08601_),
    .A2(_08602_),
    .Y(_08603_),
    .B1(net4157));
 sg13g2_a21o_1 _14177_ (.A2(_08594_),
    .A1(net1628),
    .B1(_08603_),
    .X(_00758_));
 sg13g2_nand2_1 _14178_ (.Y(_08604_),
    .A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .B(net4142));
 sg13g2_a22oi_1 _14179_ (.Y(_08605_),
    .B1(net588),
    .B2(net4149),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .A1(net5069));
 sg13g2_a21oi_1 _14180_ (.A1(_08604_),
    .A2(_08605_),
    .Y(_08606_),
    .B1(net4159));
 sg13g2_a21o_1 _14181_ (.A2(_08594_),
    .A1(net1525),
    .B1(_08606_),
    .X(_00759_));
 sg13g2_mux2_1 _14182_ (.A0(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .S(net5080),
    .X(_08607_));
 sg13g2_a22oi_1 _14183_ (.Y(_08608_),
    .B1(_08592_),
    .B2(_08607_),
    .A2(_08590_),
    .A1(\soc_inst.mem_ctrl.spi_addr[4] ));
 sg13g2_a22oi_1 _14184_ (.Y(_08609_),
    .B1(net530),
    .B2(net4150),
    .A2(net1525),
    .A1(net5069));
 sg13g2_a221oi_1 _14185_ (.B2(_08609_),
    .C1(_08588_),
    .B1(_08608_),
    .A1(_05439_),
    .Y(_08610_),
    .A2(_08585_));
 sg13g2_a21o_1 _14186_ (.A2(net4160),
    .A1(net1774),
    .B1(_08610_),
    .X(_00760_));
 sg13g2_mux2_1 _14187_ (.A0(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ),
    .S(net5080),
    .X(_08611_));
 sg13g2_a22oi_1 _14188_ (.Y(_08612_),
    .B1(_08592_),
    .B2(_08611_),
    .A2(_08590_),
    .A1(\soc_inst.mem_ctrl.spi_addr[5] ));
 sg13g2_a22oi_1 _14189_ (.Y(_08613_),
    .B1(net427),
    .B2(net4148),
    .A2(net1774),
    .A1(net5068));
 sg13g2_a221oi_1 _14190_ (.B2(_08613_),
    .C1(_08588_),
    .B1(_08612_),
    .A1(_05441_),
    .Y(_08614_),
    .A2(_08585_));
 sg13g2_a21o_1 _14191_ (.A2(net4157),
    .A1(net1791),
    .B1(_08614_),
    .X(_00761_));
 sg13g2_mux2_1 _14192_ (.A0(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .S(net5080),
    .X(_08615_));
 sg13g2_a22oi_1 _14193_ (.Y(_08616_),
    .B1(_08592_),
    .B2(_08615_),
    .A2(_08590_),
    .A1(\soc_inst.mem_ctrl.spi_addr[6] ));
 sg13g2_a22oi_1 _14194_ (.Y(_08617_),
    .B1(net429),
    .B2(net4148),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .A1(net5067));
 sg13g2_a221oi_1 _14195_ (.B2(_08617_),
    .C1(_08588_),
    .B1(_08616_),
    .A1(_05443_),
    .Y(_08618_),
    .A2(_08585_));
 sg13g2_a21o_1 _14196_ (.A2(net4158),
    .A1(net1769),
    .B1(_08618_),
    .X(_00762_));
 sg13g2_mux2_1 _14197_ (.A0(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ),
    .S(net5080),
    .X(_08619_));
 sg13g2_a22oi_1 _14198_ (.Y(_08620_),
    .B1(_08592_),
    .B2(_08619_),
    .A2(_08590_),
    .A1(\soc_inst.mem_ctrl.spi_addr[7] ));
 sg13g2_a22oi_1 _14199_ (.Y(_08621_),
    .B1(net412),
    .B2(net4149),
    .A2(net1769),
    .A1(net5067));
 sg13g2_a21oi_1 _14200_ (.A1(_08620_),
    .A2(_08621_),
    .Y(_08622_),
    .B1(_08588_));
 sg13g2_a21o_1 _14201_ (.A2(net4159),
    .A1(net1950),
    .B1(_08622_),
    .X(_00763_));
 sg13g2_nand2_1 _14202_ (.Y(_08623_),
    .A(net553),
    .B(_08594_));
 sg13g2_mux2_1 _14203_ (.A0(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .A1(\soc_inst.mem_ctrl.spi_addr[8] ),
    .S(net4280),
    .X(_08624_));
 sg13g2_a21oi_1 _14204_ (.A1(_06282_),
    .A2(_08584_),
    .Y(_08625_),
    .B1(_05501_));
 sg13g2_nand2_1 _14205_ (.Y(_08626_),
    .A(\soc_inst.mem_ctrl.spi_data_in[8] ),
    .B(net4150));
 sg13g2_a22oi_1 _14206_ (.Y(_08627_),
    .B1(_08395_),
    .B2(\soc_inst.mem_ctrl.spi_addr[8] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .A1(net5068));
 sg13g2_nand2_1 _14207_ (.Y(_08628_),
    .A(_08626_),
    .B(_08627_));
 sg13g2_a221oi_1 _14208_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ),
    .C1(_08628_),
    .B1(net4139),
    .A1(_08585_),
    .Y(_08629_),
    .A2(_08624_));
 sg13g2_o21ai_1 _14209_ (.B1(_08623_),
    .Y(_00764_),
    .A1(net4159),
    .A2(_08629_));
 sg13g2_a22oi_1 _14210_ (.Y(_08630_),
    .B1(net4138),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .A2(net4144),
    .A1(net861));
 sg13g2_nand2_1 _14211_ (.Y(_08631_),
    .A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .B(net4152));
 sg13g2_a221oi_1 _14212_ (.B2(net4148),
    .C1(net4159),
    .B1(net565),
    .A1(net5068),
    .Y(_08632_),
    .A2(net553));
 sg13g2_nand3_1 _14213_ (.B(_08631_),
    .C(_08632_),
    .A(_08630_),
    .Y(_08633_));
 sg13g2_a21oi_1 _14214_ (.A1(\soc_inst.mem_ctrl.spi_addr[9] ),
    .A2(net4142),
    .Y(_08634_),
    .B1(_08633_));
 sg13g2_a21oi_1 _14215_ (.A1(_05842_),
    .A2(net4158),
    .Y(_00765_),
    .B1(_08634_));
 sg13g2_a22oi_1 _14216_ (.Y(_08635_),
    .B1(net4139),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .A2(net4144),
    .A1(net589));
 sg13g2_nand2_1 _14217_ (.Y(_08636_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .B(net4152));
 sg13g2_a221oi_1 _14218_ (.B2(net4148),
    .C1(net4157),
    .B1(\soc_inst.mem_ctrl.spi_data_in[10] ),
    .A1(net5067),
    .Y(_08637_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ));
 sg13g2_nand3_1 _14219_ (.B(_08636_),
    .C(_08637_),
    .A(_08635_),
    .Y(_08638_));
 sg13g2_a21oi_1 _14220_ (.A1(\soc_inst.mem_ctrl.spi_addr[10] ),
    .A2(net4142),
    .Y(_08639_),
    .B1(_08638_));
 sg13g2_a21oi_1 _14221_ (.A1(_05843_),
    .A2(net4158),
    .Y(_00766_),
    .B1(_08639_));
 sg13g2_a22oi_1 _14222_ (.Y(_08640_),
    .B1(net4138),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .A2(net4144),
    .A1(net806));
 sg13g2_nand2_1 _14223_ (.Y(_08641_),
    .A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .B(net4152));
 sg13g2_a221oi_1 _14224_ (.B2(net4148),
    .C1(net4157),
    .B1(net360),
    .A1(net5067),
    .Y(_08642_),
    .A2(net589));
 sg13g2_nand3_1 _14225_ (.B(_08641_),
    .C(_08642_),
    .A(_08640_),
    .Y(_08643_));
 sg13g2_a21oi_1 _14226_ (.A1(\soc_inst.mem_ctrl.spi_addr[11] ),
    .A2(net4142),
    .Y(_08644_),
    .B1(_08643_));
 sg13g2_a21oi_1 _14227_ (.A1(_05844_),
    .A2(net4158),
    .Y(_00767_),
    .B1(_08644_));
 sg13g2_a22oi_1 _14228_ (.Y(_08645_),
    .B1(net4138),
    .B2(net553),
    .A2(net4144),
    .A1(net1395));
 sg13g2_nand2_1 _14229_ (.Y(_08646_),
    .A(\soc_inst.mem_ctrl.spi_addr[4] ),
    .B(net4152));
 sg13g2_a221oi_1 _14230_ (.B2(net4148),
    .C1(net4157),
    .B1(net580),
    .A1(net5067),
    .Y(_08647_),
    .A2(net806));
 sg13g2_nand3_1 _14231_ (.B(_08646_),
    .C(_08647_),
    .A(_08645_),
    .Y(_08648_));
 sg13g2_a21oi_1 _14232_ (.A1(\soc_inst.mem_ctrl.spi_addr[12] ),
    .A2(net4142),
    .Y(_08649_),
    .B1(_08648_));
 sg13g2_a21oi_1 _14233_ (.A1(_05845_),
    .A2(net4158),
    .Y(_00768_),
    .B1(_08649_));
 sg13g2_nand2_1 _14234_ (.Y(_08650_),
    .A(net861),
    .B(net4138));
 sg13g2_a221oi_1 _14235_ (.B2(net4148),
    .C1(net4157),
    .B1(net557),
    .A1(net5067),
    .Y(_08651_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ));
 sg13g2_a22oi_1 _14236_ (.Y(_08652_),
    .B1(net4144),
    .B2(net1031),
    .A2(net4152),
    .A1(\soc_inst.mem_ctrl.spi_addr[5] ));
 sg13g2_nand3_1 _14237_ (.B(_08651_),
    .C(_08652_),
    .A(_08650_),
    .Y(_08653_));
 sg13g2_a21oi_1 _14238_ (.A1(\soc_inst.mem_ctrl.spi_addr[13] ),
    .A2(net4142),
    .Y(_08654_),
    .B1(_08653_));
 sg13g2_a21oi_1 _14239_ (.A1(_05846_),
    .A2(net4158),
    .Y(_00769_),
    .B1(_08654_));
 sg13g2_nand2_1 _14240_ (.Y(_08655_),
    .A(net589),
    .B(net4138));
 sg13g2_a221oi_1 _14241_ (.B2(net4150),
    .C1(net4157),
    .B1(net534),
    .A1(net5068),
    .Y(_08656_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ));
 sg13g2_a22oi_1 _14242_ (.Y(_08657_),
    .B1(net4144),
    .B2(net914),
    .A2(net4152),
    .A1(\soc_inst.mem_ctrl.spi_addr[6] ));
 sg13g2_nand3_1 _14243_ (.B(_08656_),
    .C(_08657_),
    .A(_08655_),
    .Y(_08658_));
 sg13g2_a21oi_1 _14244_ (.A1(\soc_inst.mem_ctrl.spi_addr[14] ),
    .A2(net4142),
    .Y(_08659_),
    .B1(_08658_));
 sg13g2_a21oi_1 _14245_ (.A1(_05847_),
    .A2(net4158),
    .Y(_00770_),
    .B1(_08659_));
 sg13g2_a22oi_1 _14246_ (.Y(_08660_),
    .B1(net4138),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ),
    .A2(net4145),
    .A1(net704));
 sg13g2_nand2_1 _14247_ (.Y(_08661_),
    .A(\soc_inst.mem_ctrl.spi_addr[7] ),
    .B(net4152));
 sg13g2_a221oi_1 _14248_ (.B2(net4148),
    .C1(net4157),
    .B1(net488),
    .A1(net5067),
    .Y(_08662_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ));
 sg13g2_nand3_1 _14249_ (.B(_08661_),
    .C(_08662_),
    .A(_08660_),
    .Y(_08663_));
 sg13g2_a21oi_1 _14250_ (.A1(\soc_inst.mem_ctrl.spi_addr[15] ),
    .A2(net4143),
    .Y(_08664_),
    .B1(_08663_));
 sg13g2_a21oi_1 _14251_ (.A1(_05848_),
    .A2(net4160),
    .Y(_00771_),
    .B1(_08664_));
 sg13g2_nand2_1 _14252_ (.Y(_08665_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .B(net4138));
 sg13g2_a221oi_1 _14253_ (.B2(net4150),
    .C1(net4160),
    .B1(\soc_inst.mem_ctrl.spi_data_in[16] ),
    .A1(net5069),
    .Y(_08666_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ));
 sg13g2_a22oi_1 _14254_ (.Y(_08667_),
    .B1(net4145),
    .B2(net628),
    .A2(net4153),
    .A1(\soc_inst.mem_ctrl.spi_addr[8] ));
 sg13g2_nand3_1 _14255_ (.B(_08666_),
    .C(_08667_),
    .A(_08665_),
    .Y(_08668_));
 sg13g2_a21oi_1 _14256_ (.A1(\soc_inst.mem_ctrl.spi_addr[16] ),
    .A2(net4143),
    .Y(_08669_),
    .B1(_08668_));
 sg13g2_a21oi_1 _14257_ (.A1(_05849_),
    .A2(net4161),
    .Y(_00772_),
    .B1(_08669_));
 sg13g2_nand2_1 _14258_ (.Y(_08670_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ),
    .B(net4138));
 sg13g2_a221oi_1 _14259_ (.B2(net4150),
    .C1(net4156),
    .B1(net692),
    .A1(net5070),
    .Y(_08671_),
    .A2(net628));
 sg13g2_a22oi_1 _14260_ (.Y(_08672_),
    .B1(net4145),
    .B2(net852),
    .A2(net4153),
    .A1(\soc_inst.mem_ctrl.spi_addr[9] ));
 sg13g2_nand3_1 _14261_ (.B(_08671_),
    .C(_08672_),
    .A(_08670_),
    .Y(_08673_));
 sg13g2_a21oi_1 _14262_ (.A1(\soc_inst.mem_ctrl.spi_addr[17] ),
    .A2(net4143),
    .Y(_08674_),
    .B1(_08673_));
 sg13g2_a21oi_1 _14263_ (.A1(_05851_),
    .A2(net4156),
    .Y(_00773_),
    .B1(_08674_));
 sg13g2_nand2_1 _14264_ (.Y(_08675_),
    .A(net549),
    .B(_08594_));
 sg13g2_nor2_1 _14265_ (.A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .B(net4278),
    .Y(_08676_));
 sg13g2_a21oi_1 _14266_ (.A1(_05449_),
    .A2(net4278),
    .Y(_08677_),
    .B1(_08676_));
 sg13g2_nand2_1 _14267_ (.Y(_08678_),
    .A(net406),
    .B(net4149));
 sg13g2_a22oi_1 _14268_ (.Y(_08679_),
    .B1(_08395_),
    .B2(\soc_inst.mem_ctrl.spi_addr[18] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .A1(net5070));
 sg13g2_nand2_1 _14269_ (.Y(_08680_),
    .A(_08678_),
    .B(_08679_));
 sg13g2_a221oi_1 _14270_ (.B2(_08585_),
    .C1(_08680_),
    .B1(_08677_),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ),
    .Y(_08681_),
    .A2(net4139));
 sg13g2_o21ai_1 _14271_ (.B1(_08675_),
    .Y(_00774_),
    .A1(net4160),
    .A2(_08681_));
 sg13g2_nand2_1 _14272_ (.Y(_08682_),
    .A(net704),
    .B(net4139));
 sg13g2_a221oi_1 _14273_ (.B2(net4150),
    .C1(net4160),
    .B1(net414),
    .A1(net5069),
    .Y(_08683_),
    .A2(net549));
 sg13g2_a22oi_1 _14274_ (.Y(_08684_),
    .B1(net4145),
    .B2(net955),
    .A2(net4153),
    .A1(\soc_inst.mem_ctrl.spi_addr[11] ));
 sg13g2_nand3_1 _14275_ (.B(_08683_),
    .C(_08684_),
    .A(_08682_),
    .Y(_08685_));
 sg13g2_a21oi_1 _14276_ (.A1(\soc_inst.mem_ctrl.spi_addr[19] ),
    .A2(net4143),
    .Y(_08686_),
    .B1(_08685_));
 sg13g2_a21oi_1 _14277_ (.A1(_05854_),
    .A2(net4156),
    .Y(_00775_),
    .B1(_08686_));
 sg13g2_a22oi_1 _14278_ (.Y(_08687_),
    .B1(net4140),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ),
    .A2(net4145),
    .A1(net595));
 sg13g2_nand2_1 _14279_ (.Y(_08688_),
    .A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .B(net4153));
 sg13g2_a221oi_1 _14280_ (.B2(net4151),
    .C1(net4156),
    .B1(\soc_inst.mem_ctrl.spi_data_in[20] ),
    .A1(net5070),
    .Y(_08689_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ));
 sg13g2_nand3_1 _14281_ (.B(_08688_),
    .C(_08689_),
    .A(_08687_),
    .Y(_08690_));
 sg13g2_a21oi_1 _14282_ (.A1(\soc_inst.mem_ctrl.spi_addr[20] ),
    .A2(net4143),
    .Y(_08691_),
    .B1(_08690_));
 sg13g2_a21oi_1 _14283_ (.A1(_05856_),
    .A2(net4154),
    .Y(_00776_),
    .B1(_08691_));
 sg13g2_nand2_1 _14284_ (.Y(_08692_),
    .A(net515),
    .B(_08594_));
 sg13g2_mux2_1 _14285_ (.A0(\soc_inst.mem_ctrl.spi_addr[13] ),
    .A1(\soc_inst.mem_ctrl.spi_addr[21] ),
    .S(net4280),
    .X(_08693_));
 sg13g2_nand2_1 _14286_ (.Y(_08694_),
    .A(net436),
    .B(net4149));
 sg13g2_a22oi_1 _14287_ (.Y(_08695_),
    .B1(_08395_),
    .B2(\soc_inst.mem_ctrl.spi_addr[21] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ),
    .A1(net5070));
 sg13g2_nand2_1 _14288_ (.Y(_08696_),
    .A(_08694_),
    .B(_08695_));
 sg13g2_a221oi_1 _14289_ (.B2(_08585_),
    .C1(_08696_),
    .B1(_08693_),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .Y(_08697_),
    .A2(net4140));
 sg13g2_o21ai_1 _14290_ (.B1(_08692_),
    .Y(_00777_),
    .A1(net4156),
    .A2(_08697_));
 sg13g2_a21oi_1 _14291_ (.A1(_05463_),
    .A2(net4280),
    .Y(_08698_),
    .B1(_08586_));
 sg13g2_o21ai_1 _14292_ (.B1(_08698_),
    .Y(_08699_),
    .A1(\soc_inst.mem_ctrl.spi_addr[14] ),
    .A2(net4280));
 sg13g2_nand2_1 _14293_ (.Y(_08700_),
    .A(net5070),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ));
 sg13g2_o21ai_1 _14294_ (.B1(_08700_),
    .Y(_08701_),
    .A1(_05463_),
    .A2(_08394_));
 sg13g2_a221oi_1 _14295_ (.B2(net549),
    .C1(_08701_),
    .B1(net4139),
    .A1(net377),
    .Y(_08702_),
    .A2(net4150));
 sg13g2_a21oi_1 _14296_ (.A1(_08699_),
    .A2(_08702_),
    .Y(_08703_),
    .B1(net4156));
 sg13g2_a21o_1 _14297_ (.A2(_08594_),
    .A1(net1812),
    .B1(_08703_),
    .X(_00778_));
 sg13g2_a22oi_1 _14298_ (.Y(_08704_),
    .B1(net4140),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ),
    .A2(net4146),
    .A1(net740));
 sg13g2_nand2_1 _14299_ (.Y(_08705_),
    .A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .B(net4153));
 sg13g2_a221oi_1 _14300_ (.B2(net4147),
    .C1(net4156),
    .B1(net346),
    .A1(net5070),
    .Y(_08706_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ));
 sg13g2_nand3_1 _14301_ (.B(_08705_),
    .C(_08706_),
    .A(_08704_),
    .Y(_08707_));
 sg13g2_a21oi_1 _14302_ (.A1(\soc_inst.mem_ctrl.spi_addr[23] ),
    .A2(net4143),
    .Y(_08708_),
    .B1(_08707_));
 sg13g2_a21oi_1 _14303_ (.A1(_05860_),
    .A2(net4154),
    .Y(_00779_),
    .B1(_08708_));
 sg13g2_a21oi_2 _14304_ (.B1(_08585_),
    .Y(_08709_),
    .A2(_08395_),
    .A1(_05417_));
 sg13g2_a22oi_1 _14305_ (.Y(_08710_),
    .B1(net296),
    .B2(net4147),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .A1(net5071));
 sg13g2_nand2_1 _14306_ (.Y(_08711_),
    .A(_08709_),
    .B(_08710_));
 sg13g2_a221oi_1 _14307_ (.B2(net595),
    .C1(_08711_),
    .B1(net4141),
    .A1(net1880),
    .Y(_08712_),
    .A2(net4146));
 sg13g2_o21ai_1 _14308_ (.B1(_08585_),
    .Y(_08713_),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .A2(net4278));
 sg13g2_inv_1 _14309_ (.Y(_08714_),
    .A(_08713_));
 sg13g2_a21oi_1 _14310_ (.A1(\soc_inst.mem_ctrl.spi_addr[16] ),
    .A2(net4279),
    .Y(_08715_),
    .B1(_08713_));
 sg13g2_nor3_1 _14311_ (.A(net4154),
    .B(_08712_),
    .C(_08715_),
    .Y(_08716_));
 sg13g2_a21o_1 _14312_ (.A2(net4154),
    .A1(net1880),
    .B1(_08716_),
    .X(_00780_));
 sg13g2_a22oi_1 _14313_ (.Y(_08717_),
    .B1(net327),
    .B2(net4147),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ),
    .A1(net5071));
 sg13g2_nand2_1 _14314_ (.Y(_08718_),
    .A(_08709_),
    .B(_08717_));
 sg13g2_a221oi_1 _14315_ (.B2(net515),
    .C1(_08718_),
    .B1(net4141),
    .A1(net1560),
    .Y(_08719_),
    .A2(net4146));
 sg13g2_a21oi_1 _14316_ (.A1(\soc_inst.mem_ctrl.spi_addr[17] ),
    .A2(net4279),
    .Y(_08720_),
    .B1(_08713_));
 sg13g2_nor3_1 _14317_ (.A(net4154),
    .B(_08719_),
    .C(_08720_),
    .Y(_08721_));
 sg13g2_a21o_1 _14318_ (.A2(net4154),
    .A1(net1560),
    .B1(_08721_),
    .X(_00781_));
 sg13g2_a21o_1 _14319_ (.A2(net1560),
    .A1(net5070),
    .B1(net4155),
    .X(_08722_));
 sg13g2_a221oi_1 _14320_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ),
    .C1(_08722_),
    .B1(net4140),
    .A1(net313),
    .Y(_08723_),
    .A2(net4147));
 sg13g2_a22oi_1 _14321_ (.Y(_08724_),
    .B1(net4145),
    .B2(net1678),
    .A2(net4153),
    .A1(\soc_inst.mem_ctrl.spi_addr[18] ));
 sg13g2_a22oi_1 _14322_ (.Y(_00782_),
    .B1(_08723_),
    .B2(_08724_),
    .A2(net4156),
    .A1(_05862_));
 sg13g2_a22oi_1 _14323_ (.Y(_08725_),
    .B1(net213),
    .B2(net4147),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ),
    .A1(net5071));
 sg13g2_nand2b_1 _14324_ (.Y(_08726_),
    .B(_08725_),
    .A_N(_08590_));
 sg13g2_a221oi_1 _14325_ (.B2(net740),
    .C1(_08726_),
    .B1(net4141),
    .A1(net1779),
    .Y(_08727_),
    .A2(net4146));
 sg13g2_nor3_1 _14326_ (.A(\soc_inst.mem_ctrl.spi_addr[19] ),
    .B(net4280),
    .C(_08586_),
    .Y(_08728_));
 sg13g2_nor3_1 _14327_ (.A(net4154),
    .B(_08727_),
    .C(_08728_),
    .Y(_08729_));
 sg13g2_a21o_1 _14328_ (.A2(net4155),
    .A1(net1779),
    .B1(_08729_),
    .X(_00783_));
 sg13g2_o21ai_1 _14329_ (.B1(_08714_),
    .Y(_08730_),
    .A1(net2513),
    .A2(net4280));
 sg13g2_nand2_1 _14330_ (.Y(_08731_),
    .A(net264),
    .B(net4147));
 sg13g2_a221oi_1 _14331_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .C1(net4155),
    .B1(_08395_),
    .A1(net5071),
    .Y(_08732_),
    .A2(net1779));
 sg13g2_nand2_1 _14332_ (.Y(_08733_),
    .A(_08731_),
    .B(_08732_));
 sg13g2_a221oi_1 _14333_ (.B2(net1880),
    .C1(_08733_),
    .B1(net4141),
    .A1(net2599),
    .Y(_08734_),
    .A2(net4146));
 sg13g2_a22oi_1 _14334_ (.Y(_00784_),
    .B1(_08730_),
    .B2(_08734_),
    .A2(net4155),
    .A1(_05863_));
 sg13g2_a22oi_1 _14335_ (.Y(_08735_),
    .B1(net226),
    .B2(net4151),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .A1(net5071));
 sg13g2_nand2b_1 _14336_ (.Y(_08736_),
    .B(_08735_),
    .A_N(_08590_));
 sg13g2_a221oi_1 _14337_ (.B2(net1560),
    .C1(_08736_),
    .B1(net4141),
    .A1(net2884),
    .Y(_08737_),
    .A2(net4146));
 sg13g2_nor3_1 _14338_ (.A(net2486),
    .B(_06046_),
    .C(_08586_),
    .Y(_08738_));
 sg13g2_nor3_1 _14339_ (.A(net4162),
    .B(_08737_),
    .C(_08738_),
    .Y(_08739_));
 sg13g2_a21o_1 _14340_ (.A2(net4154),
    .A1(net2884),
    .B1(_08739_),
    .X(_00785_));
 sg13g2_a22oi_1 _14341_ (.Y(_08740_),
    .B1(net277),
    .B2(net4147),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .A1(net5071));
 sg13g2_nand2_1 _14342_ (.Y(_08741_),
    .A(_08709_),
    .B(_08740_));
 sg13g2_a221oi_1 _14343_ (.B2(net1678),
    .C1(_08741_),
    .B1(net4141),
    .A1(net2907),
    .Y(_08742_),
    .A2(net4146));
 sg13g2_a21oi_1 _14344_ (.A1(net1777),
    .A2(net4279),
    .Y(_08743_),
    .B1(_08713_));
 sg13g2_nor3_1 _14345_ (.A(net4155),
    .B(_08742_),
    .C(_08743_),
    .Y(_08744_));
 sg13g2_a21o_1 _14346_ (.A2(net4155),
    .A1(net2907),
    .B1(_08744_),
    .X(_00786_));
 sg13g2_nand2_1 _14347_ (.Y(_08745_),
    .A(net354),
    .B(net4147));
 sg13g2_nand2_1 _14348_ (.Y(_08746_),
    .A(net5071),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ));
 sg13g2_nand3_1 _14349_ (.B(_08745_),
    .C(_08746_),
    .A(_08709_),
    .Y(_08747_));
 sg13g2_a221oi_1 _14350_ (.B2(net1779),
    .C1(_08747_),
    .B1(net4141),
    .A1(net2861),
    .Y(_08748_),
    .A2(net4146));
 sg13g2_a21oi_1 _14351_ (.A1(net2427),
    .A2(net4279),
    .Y(_08749_),
    .B1(_08713_));
 sg13g2_nor3_1 _14352_ (.A(net4155),
    .B(_08748_),
    .C(_08749_),
    .Y(_08750_));
 sg13g2_a21o_1 _14353_ (.A2(net4155),
    .A1(net2861),
    .B1(_08750_),
    .X(_00787_));
 sg13g2_nor2_1 _14354_ (.A(net5072),
    .B(net5065),
    .Y(_08751_));
 sg13g2_a21oi_1 _14355_ (.A1(_06142_),
    .A2(_08751_),
    .Y(_08752_),
    .B1(net5077));
 sg13g2_nor2_1 _14356_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ),
    .B(_08572_),
    .Y(_08753_));
 sg13g2_nor4_1 _14357_ (.A(net5061),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .C(_05865_),
    .D(_08395_),
    .Y(_08754_));
 sg13g2_nand2b_1 _14358_ (.Y(_08755_),
    .B(_08754_),
    .A_N(_08572_));
 sg13g2_nor3_1 _14359_ (.A(_08440_),
    .B(_08446_),
    .C(_08755_),
    .Y(_08756_));
 sg13g2_a21o_2 _14360_ (.A2(_08756_),
    .A1(_08753_),
    .B1(_08752_),
    .X(_08757_));
 sg13g2_a21oi_1 _14361_ (.A1(net5066),
    .A2(net5081),
    .Y(_08758_),
    .B1(net5064));
 sg13g2_nand2_2 _14362_ (.Y(_08759_),
    .A(_05497_),
    .B(_08758_));
 sg13g2_inv_1 _14363_ (.Y(_08760_),
    .A(_08759_));
 sg13g2_nor2_1 _14364_ (.A(net5078),
    .B(uio_out[1]),
    .Y(_08761_));
 sg13g2_a21oi_1 _14365_ (.A1(net5079),
    .A2(_05863_),
    .Y(_08762_),
    .B1(_08761_));
 sg13g2_a22oi_1 _14366_ (.Y(_08763_),
    .B1(_08759_),
    .B2(_08762_),
    .A2(net2988),
    .A1(net5072));
 sg13g2_mux2_1 _14367_ (.A0(net4782),
    .A1(net4783),
    .S(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .X(_08764_));
 sg13g2_nand2_2 _14368_ (.Y(_08765_),
    .A(_08756_),
    .B(_08764_));
 sg13g2_a21oi_1 _14369_ (.A1(_08763_),
    .A2(_08765_),
    .Y(_08766_),
    .B1(_08757_));
 sg13g2_a21o_1 _14370_ (.A2(_08757_),
    .A1(net2706),
    .B1(_08766_),
    .X(_00788_));
 sg13g2_mux2_1 _14371_ (.A0(uio_out[2]),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .S(net5079),
    .X(_08767_));
 sg13g2_nand2_1 _14372_ (.Y(_08768_),
    .A(_08759_),
    .B(_08767_));
 sg13g2_nand3_1 _14373_ (.B(_08765_),
    .C(_08768_),
    .A(_08576_),
    .Y(_08769_));
 sg13g2_mux2_1 _14374_ (.A0(_08769_),
    .A1(net2774),
    .S(_08757_),
    .X(_00789_));
 sg13g2_or2_1 _14375_ (.X(_08770_),
    .B(uio_out[4]),
    .A(net5077));
 sg13g2_o21ai_1 _14376_ (.B1(_08770_),
    .Y(_08771_),
    .A1(_05501_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ));
 sg13g2_o21ai_1 _14377_ (.B1(_08765_),
    .Y(_08772_),
    .A1(_08760_),
    .A2(_08771_));
 sg13g2_mux2_1 _14378_ (.A0(_08772_),
    .A1(net2620),
    .S(_08757_),
    .X(_00790_));
 sg13g2_mux2_1 _14379_ (.A0(uio_out[5]),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ),
    .S(net5079),
    .X(_08773_));
 sg13g2_nand2_1 _14380_ (.Y(_08774_),
    .A(_08759_),
    .B(_08773_));
 sg13g2_nand3_1 _14381_ (.B(_08765_),
    .C(_08774_),
    .A(_08576_),
    .Y(_08775_));
 sg13g2_mux2_1 _14382_ (.A0(_08775_),
    .A1(net2779),
    .S(_08757_),
    .X(_00791_));
 sg13g2_or2_1 _14383_ (.X(_00792_),
    .B(net486),
    .A(net408));
 sg13g2_nand2_1 _14384_ (.Y(_08776_),
    .A(_05872_),
    .B(_08316_));
 sg13g2_nand4_1 _14385_ (.B(_05949_),
    .C(_08303_),
    .A(net4066),
    .Y(_08777_),
    .D(_08776_));
 sg13g2_nor4_1 _14386_ (.A(net2748),
    .B(net4779),
    .C(_05870_),
    .D(_08777_),
    .Y(_08778_));
 sg13g2_a21o_1 _14387_ (.A2(_08777_),
    .A1(net5075),
    .B1(_08778_),
    .X(_00793_));
 sg13g2_nor3_2 _14388_ (.A(net5057),
    .B(net4199),
    .C(net3794),
    .Y(_08779_));
 sg13g2_o21ai_1 _14389_ (.B1(net2173),
    .Y(_08780_),
    .A1(net4982),
    .A2(_08779_));
 sg13g2_nor2_1 _14390_ (.A(net4982),
    .B(_05947_),
    .Y(_08781_));
 sg13g2_a21o_2 _14391_ (.A2(_08779_),
    .A1(_05947_),
    .B1(net4982),
    .X(_08782_));
 sg13g2_a21oi_2 _14392_ (.B1(net4982),
    .Y(_08783_),
    .A2(_08779_),
    .A1(_05947_));
 sg13g2_nor2b_1 _14393_ (.A(net5057),
    .B_N(net1559),
    .Y(_08784_));
 sg13g2_a22oi_1 _14394_ (.Y(_08785_),
    .B1(net3794),
    .B2(_08784_),
    .A2(\soc_inst.cpu_core.csr_file.mepc[0] ),
    .A1(net5057));
 sg13g2_o21ai_1 _14395_ (.B1(_08780_),
    .Y(_00794_),
    .A1(net3736),
    .A2(_08785_));
 sg13g2_nor2_2 _14396_ (.A(net5114),
    .B(net5113),
    .Y(_08786_));
 sg13g2_or2_1 _14397_ (.X(_08787_),
    .B(net5113),
    .A(net5114));
 sg13g2_nor2b_2 _14398_ (.A(net5086),
    .B_N(net5084),
    .Y(_08788_));
 sg13g2_nor2_2 _14399_ (.A(net5086),
    .B(net5082),
    .Y(_08789_));
 sg13g2_nor4_1 _14400_ (.A(net5092),
    .B(net5102),
    .C(net5098),
    .D(net5095),
    .Y(_08790_));
 sg13g2_nor4_1 _14401_ (.A(net5102),
    .B(net5099),
    .C(net5098),
    .D(net5095),
    .Y(_08791_));
 sg13g2_or4_1 _14402_ (.A(net5102),
    .B(net5099),
    .C(net5098),
    .D(net5096),
    .X(_08792_));
 sg13g2_nor2_2 _14403_ (.A(net5093),
    .B(_08792_),
    .Y(_08793_));
 sg13g2_or2_1 _14404_ (.X(_08794_),
    .B(net5105),
    .A(net5107));
 sg13g2_nor4_1 _14405_ (.A(net5092),
    .B(net5089),
    .C(_08792_),
    .D(_08794_),
    .Y(_08795_));
 sg13g2_inv_1 _14406_ (.Y(_08796_),
    .A(_08795_));
 sg13g2_a21oi_1 _14407_ (.A1(_08789_),
    .A2(_08796_),
    .Y(_08797_),
    .B1(_08788_));
 sg13g2_nor2b_2 _14408_ (.A(net5082),
    .B_N(net5084),
    .Y(_08798_));
 sg13g2_nand2b_2 _14409_ (.Y(_08799_),
    .B(net5084),
    .A_N(net5083));
 sg13g2_and2_1 _14410_ (.A(net5087),
    .B(_08798_),
    .X(_08800_));
 sg13g2_nand2_1 _14411_ (.Y(_08801_),
    .A(net5086),
    .B(_08798_));
 sg13g2_or2_1 _14412_ (.X(_08802_),
    .B(net5108),
    .A(net5110));
 sg13g2_nor3_2 _14413_ (.A(net5111),
    .B(_08794_),
    .C(_08802_),
    .Y(_08803_));
 sg13g2_inv_1 _14414_ (.Y(_08804_),
    .A(_08803_));
 sg13g2_nor4_1 _14415_ (.A(net5111),
    .B(net5090),
    .C(_08794_),
    .D(_08802_),
    .Y(_08805_));
 sg13g2_nand2_2 _14416_ (.Y(_08806_),
    .A(_08800_),
    .B(net4602));
 sg13g2_nor2_2 _14417_ (.A(net5088),
    .B(net5085),
    .Y(_08807_));
 sg13g2_and2_1 _14418_ (.A(net5083),
    .B(_08807_),
    .X(_08808_));
 sg13g2_nand2_2 _14419_ (.Y(_08809_),
    .A(net5082),
    .B(_08807_));
 sg13g2_nand2_2 _14420_ (.Y(_08810_),
    .A(net5092),
    .B(net5096));
 sg13g2_nor2_1 _14421_ (.A(_08809_),
    .B(_08810_),
    .Y(_08811_));
 sg13g2_nor3_2 _14422_ (.A(_05650_),
    .B(_08809_),
    .C(_08810_),
    .Y(_08812_));
 sg13g2_nand4_1 _14423_ (.B(net5096),
    .C(net5091),
    .A(net5093),
    .Y(_08813_),
    .D(net4600));
 sg13g2_nor2b_1 _14424_ (.A(net5113),
    .B_N(net5114),
    .Y(_08814_));
 sg13g2_nand2b_2 _14425_ (.Y(_08815_),
    .B(net5114),
    .A_N(net5113));
 sg13g2_nand3_1 _14426_ (.B(_08813_),
    .C(net4694),
    .A(_08806_),
    .Y(_08816_));
 sg13g2_o21ai_1 _14427_ (.B1(_08816_),
    .Y(_08817_),
    .A1(net4696),
    .A2(net4137));
 sg13g2_nor2b_2 _14428_ (.A(net5114),
    .B_N(net5113),
    .Y(_08818_));
 sg13g2_nand2b_2 _14429_ (.Y(_08819_),
    .B(net5113),
    .A_N(net5114));
 sg13g2_nor2_1 _14430_ (.A(net5086),
    .B(_08799_),
    .Y(_08820_));
 sg13g2_and2_1 _14431_ (.A(_08793_),
    .B(net4598),
    .X(_08821_));
 sg13g2_nor2_2 _14432_ (.A(net5088),
    .B(_08821_),
    .Y(_08822_));
 sg13g2_or2_1 _14433_ (.X(_08823_),
    .B(_08821_),
    .A(net5088));
 sg13g2_nand3_1 _14434_ (.B(net4602),
    .C(net4599),
    .A(_08791_),
    .Y(_08824_));
 sg13g2_nor2_2 _14435_ (.A(net5094),
    .B(_08824_),
    .Y(_08825_));
 sg13g2_or4_1 _14436_ (.A(net5092),
    .B(net5089),
    .C(_08792_),
    .D(_08809_),
    .X(_08826_));
 sg13g2_nor2_2 _14437_ (.A(_08823_),
    .B(_08825_),
    .Y(_08827_));
 sg13g2_a21oi_2 _14438_ (.B1(_08817_),
    .Y(_08828_),
    .A2(_08827_),
    .A1(net4692));
 sg13g2_a21o_1 _14439_ (.A2(_08827_),
    .A1(net4692),
    .B1(_08817_),
    .X(_08829_));
 sg13g2_nor2_2 _14440_ (.A(\soc_inst.core_instr_addr[1] ),
    .B(_08828_),
    .Y(_08830_));
 sg13g2_xnor2_1 _14441_ (.Y(_08831_),
    .A(_05436_),
    .B(_08828_));
 sg13g2_a21oi_1 _14442_ (.A1(net2441),
    .A2(net4201),
    .Y(_08832_),
    .B1(net3793));
 sg13g2_o21ai_1 _14443_ (.B1(_08832_),
    .Y(_08833_),
    .A1(net4201),
    .A2(_08831_));
 sg13g2_a21oi_1 _14444_ (.A1(_05613_),
    .A2(net3794),
    .Y(_08834_),
    .B1(net5057));
 sg13g2_a221oi_1 _14445_ (.B2(_08834_),
    .C1(net3736),
    .B1(_08833_),
    .A1(net5057),
    .Y(_08835_),
    .A2(\soc_inst.cpu_core.csr_file.mepc[1] ));
 sg13g2_a21oi_1 _14446_ (.A1(_05436_),
    .A2(net3736),
    .Y(_00795_),
    .B1(_08835_));
 sg13g2_nor2_1 _14447_ (.A(_05437_),
    .B(_08830_),
    .Y(_08836_));
 sg13g2_xnor2_1 _14448_ (.Y(_08837_),
    .A(\soc_inst.core_instr_addr[2] ),
    .B(_08830_));
 sg13g2_a21oi_1 _14449_ (.A1(_05707_),
    .A2(net4201),
    .Y(_08838_),
    .B1(net3793));
 sg13g2_o21ai_1 _14450_ (.B1(_08838_),
    .Y(_08839_),
    .A1(net4199),
    .A2(_08837_));
 sg13g2_a21oi_1 _14451_ (.A1(net1605),
    .A2(net3794),
    .Y(_08840_),
    .B1(net5055));
 sg13g2_a221oi_1 _14452_ (.B2(_08840_),
    .C1(net3736),
    .B1(_08839_),
    .A1(net5055),
    .Y(_08841_),
    .A2(_05614_));
 sg13g2_a21o_1 _14453_ (.A2(net3734),
    .A1(net2726),
    .B1(_08841_),
    .X(_00796_));
 sg13g2_nand2_1 _14454_ (.Y(_08842_),
    .A(net2496),
    .B(net3736));
 sg13g2_nor3_1 _14455_ (.A(_05437_),
    .B(_05438_),
    .C(_08830_),
    .Y(_08843_));
 sg13g2_nor2_1 _14456_ (.A(\soc_inst.core_instr_addr[3] ),
    .B(_08836_),
    .Y(_08844_));
 sg13g2_o21ai_1 _14457_ (.B1(_06628_),
    .Y(_08845_),
    .A1(_08843_),
    .A2(_08844_));
 sg13g2_a21oi_1 _14458_ (.A1(_05708_),
    .A2(net4201),
    .Y(_08846_),
    .B1(net3793));
 sg13g2_a221oi_1 _14459_ (.B2(_08846_),
    .C1(net5057),
    .B1(_08845_),
    .A1(net499),
    .Y(_08847_),
    .A2(net3794));
 sg13g2_o21ai_1 _14460_ (.B1(_08783_),
    .Y(_08848_),
    .A1(_05474_),
    .A2(\soc_inst.cpu_core.csr_file.mepc[3] ));
 sg13g2_o21ai_1 _14461_ (.B1(_08842_),
    .Y(_00797_),
    .A1(_08847_),
    .A2(_08848_));
 sg13g2_nor4_1 _14462_ (.A(_05437_),
    .B(_05438_),
    .C(_05440_),
    .D(_08830_),
    .Y(_08849_));
 sg13g2_xnor2_1 _14463_ (.Y(_08850_),
    .A(_05440_),
    .B(_08843_));
 sg13g2_a21oi_1 _14464_ (.A1(_05709_),
    .A2(net4201),
    .Y(_08851_),
    .B1(net3793));
 sg13g2_o21ai_1 _14465_ (.B1(_08851_),
    .Y(_08852_),
    .A1(net4199),
    .A2(_08850_));
 sg13g2_a21oi_1 _14466_ (.A1(net1533),
    .A2(net3796),
    .Y(_08853_),
    .B1(net5055));
 sg13g2_o21ai_1 _14467_ (.B1(_08783_),
    .Y(_08854_),
    .A1(_05474_),
    .A2(\soc_inst.cpu_core.csr_file.mepc[4] ));
 sg13g2_a21oi_1 _14468_ (.A1(_08852_),
    .A2(_08853_),
    .Y(_08855_),
    .B1(_08854_));
 sg13g2_a21o_1 _14469_ (.A2(net3734),
    .A1(net2537),
    .B1(_08855_),
    .X(_00798_));
 sg13g2_nor2_1 _14470_ (.A(\soc_inst.core_instr_addr[5] ),
    .B(_08849_),
    .Y(_08856_));
 sg13g2_nand2_1 _14471_ (.Y(_08857_),
    .A(\soc_inst.core_instr_addr[5] ),
    .B(_08849_));
 sg13g2_nor2_1 _14472_ (.A(net4199),
    .B(_08856_),
    .Y(_08858_));
 sg13g2_a221oi_1 _14473_ (.B2(_08858_),
    .C1(net3794),
    .B1(_08857_),
    .A1(net1037),
    .Y(_08859_),
    .A2(net4201));
 sg13g2_o21ai_1 _14474_ (.B1(_05474_),
    .Y(_08860_),
    .A1(net387),
    .A2(net3800));
 sg13g2_or2_1 _14475_ (.X(_08861_),
    .B(_08860_),
    .A(_08859_));
 sg13g2_a21oi_1 _14476_ (.A1(net5055),
    .A2(net1090),
    .Y(_08862_),
    .B1(net3735));
 sg13g2_a22oi_1 _14477_ (.Y(_00799_),
    .B1(_08861_),
    .B2(_08862_),
    .A2(net3735),
    .A1(_05442_));
 sg13g2_nand3_1 _14478_ (.B(\soc_inst.core_instr_addr[6] ),
    .C(_08849_),
    .A(\soc_inst.core_instr_addr[5] ),
    .Y(_08863_));
 sg13g2_xnor2_1 _14479_ (.Y(_08864_),
    .A(_05444_),
    .B(_08857_));
 sg13g2_a21oi_1 _14480_ (.A1(net2728),
    .A2(net4201),
    .Y(_08865_),
    .B1(net3794));
 sg13g2_o21ai_1 _14481_ (.B1(_08865_),
    .Y(_08866_),
    .A1(net4199),
    .A2(_08864_));
 sg13g2_a21oi_1 _14482_ (.A1(_05617_),
    .A2(net3796),
    .Y(_08867_),
    .B1(net5055));
 sg13g2_a221oi_1 _14483_ (.B2(_08867_),
    .C1(net3734),
    .B1(_08866_),
    .A1(net5055),
    .Y(_08868_),
    .A2(net1435));
 sg13g2_a21oi_1 _14484_ (.A1(_05444_),
    .A2(net3735),
    .Y(_00800_),
    .B1(_08868_));
 sg13g2_nand4_1 _14485_ (.B(\soc_inst.core_instr_addr[6] ),
    .C(\soc_inst.core_instr_addr[7] ),
    .A(\soc_inst.core_instr_addr[5] ),
    .Y(_08869_),
    .D(_08849_));
 sg13g2_a21oi_1 _14486_ (.A1(_05445_),
    .A2(_08863_),
    .Y(_08870_),
    .B1(net4199));
 sg13g2_a22oi_1 _14487_ (.Y(_08871_),
    .B1(_08869_),
    .B2(_08870_),
    .A2(net4199),
    .A1(net2516));
 sg13g2_o21ai_1 _14488_ (.B1(_05474_),
    .Y(_08872_),
    .A1(net547),
    .A2(net3800));
 sg13g2_a21o_1 _14489_ (.A2(_08871_),
    .A1(net3800),
    .B1(_08872_),
    .X(_08873_));
 sg13g2_a21oi_1 _14490_ (.A1(net5055),
    .A2(net2683),
    .Y(_08874_),
    .B1(net3734));
 sg13g2_a22oi_1 _14491_ (.Y(_00801_),
    .B1(_08873_),
    .B2(_08874_),
    .A2(net3735),
    .A1(_05445_));
 sg13g2_and2_1 _14492_ (.A(_05446_),
    .B(_08869_),
    .X(_08875_));
 sg13g2_nor2_1 _14493_ (.A(_05446_),
    .B(_08869_),
    .Y(_08876_));
 sg13g2_nor3_1 _14494_ (.A(net4200),
    .B(_08875_),
    .C(_08876_),
    .Y(_08877_));
 sg13g2_a21oi_1 _14495_ (.A1(net1461),
    .A2(net4199),
    .Y(_08878_),
    .B1(_08877_));
 sg13g2_o21ai_1 _14496_ (.B1(_05474_),
    .Y(_08879_),
    .A1(net506),
    .A2(net3800));
 sg13g2_a21o_1 _14497_ (.A2(_08878_),
    .A1(net3800),
    .B1(_08879_),
    .X(_08880_));
 sg13g2_a21oi_1 _14498_ (.A1(net5056),
    .A2(net1016),
    .Y(_08881_),
    .B1(net3734));
 sg13g2_a22oi_1 _14499_ (.Y(_00802_),
    .B1(_08880_),
    .B2(_08881_),
    .A2(net3734),
    .A1(_05446_));
 sg13g2_nor3_1 _14500_ (.A(_05446_),
    .B(_05448_),
    .C(_08869_),
    .Y(_08882_));
 sg13g2_o21ai_1 _14501_ (.B1(_06628_),
    .Y(_08883_),
    .A1(\soc_inst.core_instr_addr[9] ),
    .A2(_08876_));
 sg13g2_nor2_1 _14502_ (.A(_08882_),
    .B(_08883_),
    .Y(_08884_));
 sg13g2_a21oi_1 _14503_ (.A1(net2208),
    .A2(net4200),
    .Y(_08885_),
    .B1(_08884_));
 sg13g2_o21ai_1 _14504_ (.B1(_05474_),
    .Y(_08886_),
    .A1(net664),
    .A2(net3800));
 sg13g2_a21o_1 _14505_ (.A2(_08885_),
    .A1(net3801),
    .B1(_08886_),
    .X(_08887_));
 sg13g2_a21oi_1 _14506_ (.A1(net5054),
    .A2(net999),
    .Y(_08888_),
    .B1(net3734));
 sg13g2_a22oi_1 _14507_ (.Y(_00803_),
    .B1(_08887_),
    .B2(_08888_),
    .A2(net3734),
    .A1(_05448_));
 sg13g2_nor2_1 _14508_ (.A(net2771),
    .B(_08783_),
    .Y(_08889_));
 sg13g2_nor4_1 _14509_ (.A(_05446_),
    .B(_05448_),
    .C(_05450_),
    .D(_08869_),
    .Y(_08890_));
 sg13g2_xnor2_1 _14510_ (.Y(_08891_),
    .A(\soc_inst.core_instr_addr[10] ),
    .B(_08882_));
 sg13g2_a21oi_1 _14511_ (.A1(net2263),
    .A2(net4200),
    .Y(_08892_),
    .B1(net3795));
 sg13g2_o21ai_1 _14512_ (.B1(_08892_),
    .Y(_08893_),
    .A1(net4200),
    .A2(_08891_));
 sg13g2_a21oi_1 _14513_ (.A1(_05622_),
    .A2(net3796),
    .Y(_08894_),
    .B1(net5055));
 sg13g2_a22oi_1 _14514_ (.Y(_08895_),
    .B1(_08893_),
    .B2(_08894_),
    .A2(net1208),
    .A1(net5056));
 sg13g2_a21oi_1 _14515_ (.A1(_08783_),
    .A2(_08895_),
    .Y(_00804_),
    .B1(_08889_));
 sg13g2_and2_1 _14516_ (.A(\soc_inst.core_instr_addr[11] ),
    .B(_08890_),
    .X(_08896_));
 sg13g2_o21ai_1 _14517_ (.B1(_06628_),
    .Y(_08897_),
    .A1(\soc_inst.core_instr_addr[11] ),
    .A2(_08890_));
 sg13g2_nor2_1 _14518_ (.A(_08896_),
    .B(_08897_),
    .Y(_08898_));
 sg13g2_a21oi_1 _14519_ (.A1(net1825),
    .A2(net4200),
    .Y(_08899_),
    .B1(_08898_));
 sg13g2_o21ai_1 _14520_ (.B1(_05474_),
    .Y(_08900_),
    .A1(net450),
    .A2(net3800));
 sg13g2_a21o_1 _14521_ (.A2(_08899_),
    .A1(net3799),
    .B1(_08900_),
    .X(_08901_));
 sg13g2_a21oi_1 _14522_ (.A1(net5057),
    .A2(net2484),
    .Y(_08902_),
    .B1(net3736));
 sg13g2_a22oi_1 _14523_ (.Y(_00805_),
    .B1(_08901_),
    .B2(_08902_),
    .A2(net3736),
    .A1(_05452_));
 sg13g2_xnor2_1 _14524_ (.Y(_08903_),
    .A(\soc_inst.core_instr_addr[12] ),
    .B(_08896_));
 sg13g2_a21oi_1 _14525_ (.A1(net1322),
    .A2(net4196),
    .Y(_08904_),
    .B1(net3792));
 sg13g2_o21ai_1 _14526_ (.B1(_08904_),
    .Y(_08905_),
    .A1(net4197),
    .A2(_08903_));
 sg13g2_a21oi_1 _14527_ (.A1(_05625_),
    .A2(net3792),
    .Y(_08906_),
    .B1(net5053));
 sg13g2_a221oi_1 _14528_ (.B2(_08906_),
    .C1(net3733),
    .B1(_08905_),
    .A1(net5053),
    .Y(_08907_),
    .A2(net2559));
 sg13g2_a21oi_1 _14529_ (.A1(_05453_),
    .A2(net3733),
    .Y(_00806_),
    .B1(_08907_));
 sg13g2_a21oi_1 _14530_ (.A1(\soc_inst.core_instr_addr[12] ),
    .A2(_08896_),
    .Y(_08908_),
    .B1(\soc_inst.core_instr_addr[13] ));
 sg13g2_nand3_1 _14531_ (.B(\soc_inst.core_instr_addr[13] ),
    .C(_08896_),
    .A(\soc_inst.core_instr_addr[12] ),
    .Y(_08909_));
 sg13g2_nor2_1 _14532_ (.A(net4200),
    .B(_08908_),
    .Y(_08910_));
 sg13g2_a22oi_1 _14533_ (.Y(_08911_),
    .B1(_08909_),
    .B2(_08910_),
    .A2(net4197),
    .A1(net2352));
 sg13g2_o21ai_1 _14534_ (.B1(_05474_),
    .Y(_08912_),
    .A1(net945),
    .A2(net3799));
 sg13g2_a21o_1 _14535_ (.A2(_08911_),
    .A1(net3799),
    .B1(_08912_),
    .X(_08913_));
 sg13g2_a21oi_1 _14536_ (.A1(net5058),
    .A2(net789),
    .Y(_08914_),
    .B1(net3731));
 sg13g2_a22oi_1 _14537_ (.Y(_00807_),
    .B1(_08913_),
    .B2(_08914_),
    .A2(net3731),
    .A1(_05454_));
 sg13g2_nor2_1 _14538_ (.A(net2762),
    .B(_08783_),
    .Y(_08915_));
 sg13g2_and4_1 _14539_ (.A(\soc_inst.core_instr_addr[12] ),
    .B(\soc_inst.core_instr_addr[13] ),
    .C(\soc_inst.core_instr_addr[14] ),
    .D(_08896_),
    .X(_08916_));
 sg13g2_xnor2_1 _14540_ (.Y(_08917_),
    .A(_05455_),
    .B(_08909_));
 sg13g2_a21oi_1 _14541_ (.A1(\soc_inst.cpu_core.ex_branch_target[14] ),
    .A2(net4196),
    .Y(_08918_),
    .B1(net3795));
 sg13g2_o21ai_1 _14542_ (.B1(_08918_),
    .Y(_08919_),
    .A1(net4200),
    .A2(_08917_));
 sg13g2_a21oi_1 _14543_ (.A1(_05628_),
    .A2(net3796),
    .Y(_08920_),
    .B1(net5054));
 sg13g2_a22oi_1 _14544_ (.Y(_08921_),
    .B1(_08919_),
    .B2(_08920_),
    .A2(net1914),
    .A1(net5054));
 sg13g2_a21oi_1 _14545_ (.A1(_08783_),
    .A2(_08921_),
    .Y(_00808_),
    .B1(_08915_));
 sg13g2_nand2_1 _14546_ (.Y(_08922_),
    .A(\soc_inst.core_instr_addr[15] ),
    .B(_08916_));
 sg13g2_xnor2_1 _14547_ (.Y(_08923_),
    .A(\soc_inst.core_instr_addr[15] ),
    .B(_08916_));
 sg13g2_a21oi_1 _14548_ (.A1(net508),
    .A2(net4198),
    .Y(_08924_),
    .B1(net3792));
 sg13g2_o21ai_1 _14549_ (.B1(_08924_),
    .Y(_08925_),
    .A1(net4198),
    .A2(_08923_));
 sg13g2_a21oi_1 _14550_ (.A1(_05630_),
    .A2(net3792),
    .Y(_08926_),
    .B1(net5053));
 sg13g2_a221oi_1 _14551_ (.B2(_08926_),
    .C1(net3731),
    .B1(_08925_),
    .A1(net5053),
    .Y(_08927_),
    .A2(net832));
 sg13g2_a21oi_1 _14552_ (.A1(_05456_),
    .A2(net3731),
    .Y(_00809_),
    .B1(_08927_));
 sg13g2_nand3_1 _14553_ (.B(\soc_inst.core_instr_addr[16] ),
    .C(_08916_),
    .A(\soc_inst.core_instr_addr[15] ),
    .Y(_08928_));
 sg13g2_xnor2_1 _14554_ (.Y(_08929_),
    .A(_05457_),
    .B(_08922_));
 sg13g2_a21oi_1 _14555_ (.A1(net2746),
    .A2(net4195),
    .Y(_08930_),
    .B1(net3790));
 sg13g2_o21ai_1 _14556_ (.B1(_08930_),
    .Y(_08931_),
    .A1(net4197),
    .A2(_08929_));
 sg13g2_a21oi_1 _14557_ (.A1(_05632_),
    .A2(net3797),
    .Y(_08932_),
    .B1(net5052));
 sg13g2_a221oi_1 _14558_ (.B2(_08932_),
    .C1(net3732),
    .B1(_08931_),
    .A1(net5052),
    .Y(_08933_),
    .A2(net2061));
 sg13g2_a21oi_1 _14559_ (.A1(_05457_),
    .A2(net3732),
    .Y(_00810_),
    .B1(_08933_));
 sg13g2_and4_1 _14560_ (.A(\soc_inst.core_instr_addr[15] ),
    .B(\soc_inst.core_instr_addr[16] ),
    .C(\soc_inst.core_instr_addr[17] ),
    .D(_08916_),
    .X(_08934_));
 sg13g2_xnor2_1 _14561_ (.Y(_08935_),
    .A(_05458_),
    .B(_08928_));
 sg13g2_a21oi_1 _14562_ (.A1(net1301),
    .A2(net4195),
    .Y(_08936_),
    .B1(net3790));
 sg13g2_o21ai_1 _14563_ (.B1(_08936_),
    .Y(_08937_),
    .A1(net4197),
    .A2(_08935_));
 sg13g2_a21oi_1 _14564_ (.A1(_05634_),
    .A2(net3792),
    .Y(_08938_),
    .B1(net5052));
 sg13g2_a221oi_1 _14565_ (.B2(_08938_),
    .C1(net3732),
    .B1(_08937_),
    .A1(net5053),
    .Y(_08939_),
    .A2(net2115));
 sg13g2_a21oi_1 _14566_ (.A1(_05458_),
    .A2(net3732),
    .Y(_00811_),
    .B1(_08939_));
 sg13g2_xnor2_1 _14567_ (.Y(_08940_),
    .A(\soc_inst.core_instr_addr[18] ),
    .B(_08934_));
 sg13g2_a21oi_1 _14568_ (.A1(net2520),
    .A2(net4195),
    .Y(_08941_),
    .B1(net3791));
 sg13g2_o21ai_1 _14569_ (.B1(_08941_),
    .Y(_08942_),
    .A1(net4197),
    .A2(_08940_));
 sg13g2_a21oi_1 _14570_ (.A1(_05636_),
    .A2(net3791),
    .Y(_08943_),
    .B1(net5051));
 sg13g2_a221oi_1 _14571_ (.B2(_08943_),
    .C1(net3730),
    .B1(_08942_),
    .A1(net5051),
    .Y(_08944_),
    .A2(net1104));
 sg13g2_a21oi_1 _14572_ (.A1(_05459_),
    .A2(net3730),
    .Y(_00812_),
    .B1(_08944_));
 sg13g2_a21oi_1 _14573_ (.A1(\soc_inst.core_instr_addr[18] ),
    .A2(_08934_),
    .Y(_08945_),
    .B1(\soc_inst.core_instr_addr[19] ));
 sg13g2_nand3_1 _14574_ (.B(\soc_inst.core_instr_addr[19] ),
    .C(_08934_),
    .A(\soc_inst.core_instr_addr[18] ),
    .Y(_08946_));
 sg13g2_nand2_1 _14575_ (.Y(_08947_),
    .A(_06628_),
    .B(_08946_));
 sg13g2_a21oi_1 _14576_ (.A1(net2062),
    .A2(net4195),
    .Y(_08948_),
    .B1(net3790));
 sg13g2_o21ai_1 _14577_ (.B1(_08948_),
    .Y(_08949_),
    .A1(_08945_),
    .A2(_08947_));
 sg13g2_a21oi_1 _14578_ (.A1(_05638_),
    .A2(net3791),
    .Y(_08950_),
    .B1(net5052));
 sg13g2_a221oi_1 _14579_ (.B2(_08950_),
    .C1(net3730),
    .B1(_08949_),
    .A1(net5051),
    .Y(_08951_),
    .A2(net1307));
 sg13g2_a21oi_1 _14580_ (.A1(_05460_),
    .A2(net3730),
    .Y(_00813_),
    .B1(_08951_));
 sg13g2_and4_1 _14581_ (.A(\soc_inst.core_instr_addr[18] ),
    .B(\soc_inst.core_instr_addr[19] ),
    .C(\soc_inst.core_instr_addr[20] ),
    .D(_08934_),
    .X(_08952_));
 sg13g2_xnor2_1 _14582_ (.Y(_08953_),
    .A(_05461_),
    .B(_08946_));
 sg13g2_a21oi_1 _14583_ (.A1(net2225),
    .A2(net4197),
    .Y(_08954_),
    .B1(net3790));
 sg13g2_o21ai_1 _14584_ (.B1(_08954_),
    .Y(_08955_),
    .A1(net4197),
    .A2(_08953_));
 sg13g2_a21oi_1 _14585_ (.A1(_05640_),
    .A2(net3797),
    .Y(_08956_),
    .B1(net5052));
 sg13g2_a221oi_1 _14586_ (.B2(_08956_),
    .C1(net3732),
    .B1(_08955_),
    .A1(net5052),
    .Y(_08957_),
    .A2(net1634));
 sg13g2_a21oi_1 _14587_ (.A1(_05461_),
    .A2(net3732),
    .Y(_00814_),
    .B1(_08957_));
 sg13g2_xnor2_1 _14588_ (.Y(_08958_),
    .A(\soc_inst.core_instr_addr[21] ),
    .B(_08952_));
 sg13g2_a21oi_1 _14589_ (.A1(net2350),
    .A2(net4195),
    .Y(_08959_),
    .B1(net3790));
 sg13g2_o21ai_1 _14590_ (.B1(_08959_),
    .Y(_08960_),
    .A1(net4195),
    .A2(_08958_));
 sg13g2_a21oi_1 _14591_ (.A1(_05642_),
    .A2(net3790),
    .Y(_08961_),
    .B1(net5051));
 sg13g2_a221oi_1 _14592_ (.B2(_08961_),
    .C1(net3730),
    .B1(_08960_),
    .A1(net5051),
    .Y(_08962_),
    .A2(net1713));
 sg13g2_a21oi_1 _14593_ (.A1(_05462_),
    .A2(net3730),
    .Y(_00815_),
    .B1(_08962_));
 sg13g2_a21oi_1 _14594_ (.A1(\soc_inst.core_instr_addr[21] ),
    .A2(_08952_),
    .Y(_08963_),
    .B1(net2854));
 sg13g2_nand3_1 _14595_ (.B(\soc_inst.core_instr_addr[22] ),
    .C(_08952_),
    .A(\soc_inst.core_instr_addr[21] ),
    .Y(_08964_));
 sg13g2_nand2_1 _14596_ (.Y(_08965_),
    .A(_06628_),
    .B(_08964_));
 sg13g2_a21oi_1 _14597_ (.A1(net2768),
    .A2(net4195),
    .Y(_08966_),
    .B1(net3790));
 sg13g2_o21ai_1 _14598_ (.B1(_08966_),
    .Y(_08967_),
    .A1(_08963_),
    .A2(_08965_));
 sg13g2_a21oi_1 _14599_ (.A1(_05644_),
    .A2(net3792),
    .Y(_08968_),
    .B1(net5052));
 sg13g2_a221oi_1 _14600_ (.B2(_08968_),
    .C1(net3732),
    .B1(_08967_),
    .A1(net5052),
    .Y(_08969_),
    .A2(net925));
 sg13g2_a21oi_1 _14601_ (.A1(_05464_),
    .A2(net3732),
    .Y(_00816_),
    .B1(_08969_));
 sg13g2_xnor2_1 _14602_ (.Y(_08970_),
    .A(_05465_),
    .B(_08964_));
 sg13g2_a21oi_1 _14603_ (.A1(net1069),
    .A2(net4195),
    .Y(_08971_),
    .B1(net3790));
 sg13g2_o21ai_1 _14604_ (.B1(_08971_),
    .Y(_08972_),
    .A1(net4197),
    .A2(_08970_));
 sg13g2_a21oi_1 _14605_ (.A1(_05646_),
    .A2(net3791),
    .Y(_08973_),
    .B1(net5051));
 sg13g2_a221oi_1 _14606_ (.B2(_08973_),
    .C1(net3730),
    .B1(_08972_),
    .A1(net5051),
    .Y(_08974_),
    .A2(net1949));
 sg13g2_a21oi_1 _14607_ (.A1(_05465_),
    .A2(net3730),
    .Y(_00817_),
    .B1(_08974_));
 sg13g2_a21oi_1 _14608_ (.A1(net4872),
    .A2(net2334),
    .Y(_08975_),
    .B1(_06755_));
 sg13g2_nand4_1 _14609_ (.B(net4255),
    .C(net4707),
    .A(net2334),
    .Y(_08976_),
    .D(_06754_));
 sg13g2_o21ai_1 _14610_ (.B1(_08976_),
    .Y(_08977_),
    .A1(net4231),
    .A2(_08975_));
 sg13g2_mux2_1 _14611_ (.A0(_08977_),
    .A1(net2334),
    .S(net3855),
    .X(_00818_));
 sg13g2_a21oi_1 _14612_ (.A1(net4872),
    .A2(net2395),
    .Y(_08978_),
    .B1(_06767_));
 sg13g2_nand4_1 _14613_ (.B(net4255),
    .C(net4707),
    .A(net2395),
    .Y(_08979_),
    .D(_06766_));
 sg13g2_o21ai_1 _14614_ (.B1(_08979_),
    .Y(_08980_),
    .A1(net4231),
    .A2(_08978_));
 sg13g2_mux2_1 _14615_ (.A0(_08980_),
    .A1(net2395),
    .S(net3855),
    .X(_00819_));
 sg13g2_a21oi_1 _14616_ (.A1(net4871),
    .A2(net2011),
    .Y(_08981_),
    .B1(_06775_));
 sg13g2_nand4_1 _14617_ (.B(net4255),
    .C(net4707),
    .A(net2011),
    .Y(_08982_),
    .D(_06774_));
 sg13g2_o21ai_1 _14618_ (.B1(_08982_),
    .Y(_08983_),
    .A1(net4230),
    .A2(_08981_));
 sg13g2_mux2_1 _14619_ (.A0(_08983_),
    .A1(net2011),
    .S(net3855),
    .X(_00820_));
 sg13g2_a21oi_1 _14620_ (.A1(net4872),
    .A2(net2401),
    .Y(_08984_),
    .B1(_06788_));
 sg13g2_nand4_1 _14621_ (.B(net4255),
    .C(net4707),
    .A(net2401),
    .Y(_08985_),
    .D(_06787_));
 sg13g2_o21ai_1 _14622_ (.B1(_08985_),
    .Y(_08986_),
    .A1(net4231),
    .A2(_08984_));
 sg13g2_mux2_1 _14623_ (.A0(_08986_),
    .A1(net2401),
    .S(net3855),
    .X(_00821_));
 sg13g2_nor2_1 _14624_ (.A(net2059),
    .B(net1801),
    .Y(_08987_));
 sg13g2_nand3b_1 _14625_ (.B(net517),
    .C(_08987_),
    .Y(_08988_),
    .A_N(net2972));
 sg13g2_nand3_1 _14626_ (.B(net5060),
    .C(_08988_),
    .A(net2738),
    .Y(_08989_));
 sg13g2_and2_1 _14627_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ),
    .B(_07850_),
    .X(_08990_));
 sg13g2_nand2_1 _14628_ (.Y(_08991_),
    .A(net2880),
    .B(_07850_));
 sg13g2_nand4_1 _14629_ (.B(_05393_),
    .C(net5060),
    .A(net869),
    .Y(_08992_),
    .D(_08987_));
 sg13g2_nand3_1 _14630_ (.B(net4596),
    .C(_08992_),
    .A(_08989_),
    .Y(_08993_));
 sg13g2_nand2_1 _14631_ (.Y(_08994_),
    .A(net5480),
    .B(_08993_));
 sg13g2_nand2b_1 _14632_ (.Y(_08995_),
    .B(net2738),
    .A_N(net5060));
 sg13g2_xor2_1 _14633_ (.B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ),
    .A(_00330_),
    .X(_08996_));
 sg13g2_or2_1 _14634_ (.X(_08997_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .A(_00329_));
 sg13g2_xnor2_1 _14635_ (.Y(_08998_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ));
 sg13g2_nand2b_1 _14636_ (.Y(_08999_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ),
    .A_N(net4759));
 sg13g2_o21ai_1 _14637_ (.B1(_08999_),
    .Y(_09000_),
    .A1(_00327_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ));
 sg13g2_a221oi_1 _14638_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .C1(_09000_),
    .B1(_05392_),
    .A1(_00329_),
    .Y(_09001_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ));
 sg13g2_a22oi_1 _14639_ (.Y(_09002_),
    .B1(_05413_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ),
    .A2(_05412_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ));
 sg13g2_xnor2_1 _14640_ (.Y(_09003_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ));
 sg13g2_xnor2_1 _14641_ (.Y(_09004_),
    .A(_00328_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ));
 sg13g2_o21ai_1 _14642_ (.B1(_08997_),
    .Y(_09005_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .A2(_05412_));
 sg13g2_nand3_1 _14643_ (.B(_08998_),
    .C(_09003_),
    .A(_08996_),
    .Y(_09006_));
 sg13g2_a22oi_1 _14644_ (.Y(_09007_),
    .B1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .B2(_05411_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ),
    .A1(_00327_));
 sg13g2_a221oi_1 _14645_ (.B2(_05390_),
    .C1(_09005_),
    .B1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .A1(_05391_),
    .Y(_09008_),
    .A2(net4759));
 sg13g2_nand4_1 _14646_ (.B(_09002_),
    .C(_09007_),
    .A(_09001_),
    .Y(_09009_),
    .D(_09008_));
 sg13g2_nor3_2 _14647_ (.A(_09004_),
    .B(_09006_),
    .C(_09009_),
    .Y(_09010_));
 sg13g2_nand2b_2 _14648_ (.Y(_09011_),
    .B(net5472),
    .A_N(_09010_));
 sg13g2_o21ai_1 _14649_ (.B1(_08994_),
    .Y(_00822_),
    .A1(_08995_),
    .A2(_09011_));
 sg13g2_nand2_1 _14650_ (.Y(_09012_),
    .A(_05410_),
    .B(net5060));
 sg13g2_nand2b_1 _14651_ (.Y(_09013_),
    .B(_09010_),
    .A_N(_08995_));
 sg13g2_nand3_1 _14652_ (.B(_09012_),
    .C(_09013_),
    .A(_08989_),
    .Y(_09014_));
 sg13g2_and2_1 _14653_ (.A(net5480),
    .B(_09014_),
    .X(_00823_));
 sg13g2_nor2_1 _14654_ (.A(net1369),
    .B(net3759),
    .Y(_09015_));
 sg13g2_nand2b_1 _14655_ (.Y(_09016_),
    .B(_06754_),
    .A_N(net1369));
 sg13g2_a21oi_1 _14656_ (.A1(_06757_),
    .A2(_09016_),
    .Y(_09017_),
    .B1(_07632_));
 sg13g2_a21oi_1 _14657_ (.A1(net3759),
    .A2(_09017_),
    .Y(_00824_),
    .B1(_09015_));
 sg13g2_nor2_1 _14658_ (.A(net1406),
    .B(net3760),
    .Y(_09018_));
 sg13g2_nand2b_1 _14659_ (.Y(_09019_),
    .B(_06766_),
    .A_N(net1406));
 sg13g2_a21oi_1 _14660_ (.A1(_06769_),
    .A2(_09019_),
    .Y(_09020_),
    .B1(_07636_));
 sg13g2_a21oi_1 _14661_ (.A1(net3760),
    .A2(_09020_),
    .Y(_00825_),
    .B1(_09018_));
 sg13g2_nor2_1 _14662_ (.A(net843),
    .B(net3759),
    .Y(_09021_));
 sg13g2_nand2b_1 _14663_ (.Y(_09022_),
    .B(_06774_),
    .A_N(net843));
 sg13g2_a21oi_1 _14664_ (.A1(_06777_),
    .A2(_09022_),
    .Y(_09023_),
    .B1(_07640_));
 sg13g2_a21oi_1 _14665_ (.A1(net3759),
    .A2(_09023_),
    .Y(_00826_),
    .B1(_09021_));
 sg13g2_a21oi_1 _14666_ (.A1(_06741_),
    .A2(net3759),
    .Y(_09024_),
    .B1(net356));
 sg13g2_a21oi_1 _14667_ (.A1(_06743_),
    .A2(net3759),
    .Y(_00827_),
    .B1(_09024_));
 sg13g2_nor2_1 _14668_ (.A(net759),
    .B(net3759),
    .Y(_09025_));
 sg13g2_nand2b_1 _14669_ (.Y(_09026_),
    .B(_06787_),
    .A_N(net759));
 sg13g2_a21oi_1 _14670_ (.A1(_06790_),
    .A2(_09026_),
    .Y(_09027_),
    .B1(_07645_));
 sg13g2_a21oi_1 _14671_ (.A1(net3759),
    .A2(_09027_),
    .Y(_00828_),
    .B1(_09025_));
 sg13g2_nand2_1 _14672_ (.Y(_09028_),
    .A(_08459_),
    .B(_08754_));
 sg13g2_nand2_1 _14673_ (.Y(_09029_),
    .A(_07068_),
    .B(_09028_));
 sg13g2_a21o_2 _14674_ (.A2(_08581_),
    .A1(net97),
    .B1(_09029_),
    .X(_09030_));
 sg13g2_nand2_1 _14675_ (.Y(_09031_),
    .A(_06122_),
    .B(_06282_));
 sg13g2_nor2_1 _14676_ (.A(net5081),
    .B(_09031_),
    .Y(_09032_));
 sg13g2_nor2_1 _14677_ (.A(net5077),
    .B(_09032_),
    .Y(_09033_));
 sg13g2_o21ai_1 _14678_ (.B1(net2899),
    .Y(_09034_),
    .A1(net5077),
    .A2(_09032_));
 sg13g2_nor3_1 _14679_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .B(net5078),
    .C(_08581_),
    .Y(_09035_));
 sg13g2_nor2_1 _14680_ (.A(net5066),
    .B(_09031_),
    .Y(_09036_));
 sg13g2_nor2_1 _14681_ (.A(_09035_),
    .B(_09036_),
    .Y(_09037_));
 sg13g2_nor3_2 _14682_ (.A(net5064),
    .B(_08440_),
    .C(_08755_),
    .Y(_09038_));
 sg13g2_inv_1 _14683_ (.Y(_09039_),
    .A(_09038_));
 sg13g2_nand2_1 _14684_ (.Y(_09040_),
    .A(_06128_),
    .B(_09039_));
 sg13g2_or2_1 _14685_ (.X(_09041_),
    .B(_09040_),
    .A(net5072));
 sg13g2_nand3_1 _14686_ (.B(net4783),
    .C(net5077),
    .A(net4782),
    .Y(_09042_));
 sg13g2_xnor2_1 _14687_ (.Y(_09043_),
    .A(net2899),
    .B(_09042_));
 sg13g2_a221oi_1 _14688_ (.B2(_09043_),
    .C1(_09030_),
    .B1(_09041_),
    .A1(_09034_),
    .Y(_09044_),
    .A2(_09037_));
 sg13g2_a21oi_1 _14689_ (.A1(_05491_),
    .A2(_09030_),
    .Y(_00829_),
    .B1(_09044_));
 sg13g2_o21ai_1 _14690_ (.B1(_05492_),
    .Y(_09045_),
    .A1(_05491_),
    .A2(_09042_));
 sg13g2_and3_1 _14691_ (.X(_09046_),
    .A(net4782),
    .B(net4783),
    .C(_06151_));
 sg13g2_nor2_1 _14692_ (.A(net5065),
    .B(_09038_),
    .Y(_09047_));
 sg13g2_a22oi_1 _14693_ (.Y(_09048_),
    .B1(_09047_),
    .B2(_06043_),
    .A2(_09046_),
    .A1(net5077));
 sg13g2_o21ai_1 _14694_ (.B1(_09045_),
    .Y(_09049_),
    .A1(_09030_),
    .A2(_09048_));
 sg13g2_nor3_1 _14695_ (.A(_06037_),
    .B(_06125_),
    .C(_09033_),
    .Y(_09050_));
 sg13g2_a21o_1 _14696_ (.A2(_08581_),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .B1(net5078),
    .X(_09051_));
 sg13g2_nor2_1 _14697_ (.A(_09036_),
    .B(_09050_),
    .Y(_09052_));
 sg13g2_o21ai_1 _14698_ (.B1(_09052_),
    .Y(_09053_),
    .A1(net2868),
    .A2(_09051_));
 sg13g2_a22oi_1 _14699_ (.Y(_00830_),
    .B1(_09049_),
    .B2(_09053_),
    .A2(_09030_),
    .A1(_05492_));
 sg13g2_nand2_1 _14700_ (.Y(_09054_),
    .A(_05494_),
    .B(_05501_));
 sg13g2_nor2b_2 _14701_ (.A(_09038_),
    .B_N(_08751_),
    .Y(_09055_));
 sg13g2_a21oi_1 _14702_ (.A1(net5059),
    .A2(_09046_),
    .Y(_09056_),
    .B1(_09055_));
 sg13g2_o21ai_1 _14703_ (.B1(_09056_),
    .Y(_09057_),
    .A1(net5059),
    .A2(_09046_));
 sg13g2_o21ai_1 _14704_ (.B1(_09039_),
    .Y(_09058_),
    .A1(net5059),
    .A2(_06151_));
 sg13g2_nor2b_1 _14705_ (.A(_09058_),
    .B_N(_08389_),
    .Y(_09059_));
 sg13g2_inv_1 _14706_ (.Y(_09060_),
    .A(_09059_));
 sg13g2_a22oi_1 _14707_ (.Y(_09061_),
    .B1(_09060_),
    .B2(net5078),
    .A2(_08758_),
    .A1(_06282_));
 sg13g2_o21ai_1 _14708_ (.B1(_09057_),
    .Y(_09062_),
    .A1(net5077),
    .A2(_09055_));
 sg13g2_or2_1 _14709_ (.X(_09063_),
    .B(_09062_),
    .A(_09061_));
 sg13g2_nand3_1 _14710_ (.B(_08581_),
    .C(_09059_),
    .A(_08393_),
    .Y(_09064_));
 sg13g2_a21oi_1 _14711_ (.A1(_09054_),
    .A2(_09063_),
    .Y(_09065_),
    .B1(_09030_));
 sg13g2_a22oi_1 _14712_ (.Y(_00831_),
    .B1(_09064_),
    .B2(_09065_),
    .A2(_09030_),
    .A1(_05494_));
 sg13g2_a21oi_1 _14713_ (.A1(_08760_),
    .A2(_09055_),
    .Y(_09066_),
    .B1(net5079));
 sg13g2_nor3_1 _14714_ (.A(_09030_),
    .B(_09056_),
    .C(_09066_),
    .Y(_09067_));
 sg13g2_nand2b_1 _14715_ (.Y(_09068_),
    .B(net2373),
    .A_N(_09067_));
 sg13g2_nand2_1 _14716_ (.Y(_09069_),
    .A(_05493_),
    .B(_05501_));
 sg13g2_a22oi_1 _14717_ (.Y(_09070_),
    .B1(_08759_),
    .B2(_09069_),
    .A2(_08581_),
    .A1(_08393_));
 sg13g2_xnor2_1 _14718_ (.Y(_09071_),
    .A(_05493_),
    .B(_08389_));
 sg13g2_nor3_1 _14719_ (.A(_09038_),
    .B(_09070_),
    .C(_09071_),
    .Y(_09072_));
 sg13g2_nor4_1 _14720_ (.A(net2373),
    .B(_08389_),
    .C(_09042_),
    .D(_09055_),
    .Y(_09073_));
 sg13g2_nor2_1 _14721_ (.A(_09072_),
    .B(_09073_),
    .Y(_09074_));
 sg13g2_o21ai_1 _14722_ (.B1(_09068_),
    .Y(_00832_),
    .A1(_09030_),
    .A2(_09074_));
 sg13g2_xor2_1 _14723_ (.B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ),
    .A(net460),
    .X(_00833_));
 sg13g2_nand3_1 _14724_ (.B(net2844),
    .C(net2578),
    .A(net460),
    .Y(_09075_));
 sg13g2_a21o_1 _14725_ (.A2(net2578),
    .A1(net460),
    .B1(net2844),
    .X(_09076_));
 sg13g2_and2_1 _14726_ (.A(_09075_),
    .B(_09076_),
    .X(_00834_));
 sg13g2_nand4_1 _14727_ (.B(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .Y(_09077_),
    .D(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ));
 sg13g2_xnor2_1 _14728_ (.Y(_00835_),
    .A(net401),
    .B(_09075_));
 sg13g2_nor2_2 _14729_ (.A(_05506_),
    .B(_06135_),
    .Y(_09078_));
 sg13g2_a21oi_1 _14730_ (.A1(_05504_),
    .A2(_09077_),
    .Y(_00836_),
    .B1(_09078_));
 sg13g2_and2_1 _14731_ (.A(net217),
    .B(_09078_),
    .X(_09079_));
 sg13g2_xor2_1 _14732_ (.B(_09078_),
    .A(net217),
    .X(_00837_));
 sg13g2_xor2_1 _14733_ (.B(_09079_),
    .A(net245),
    .X(_00838_));
 sg13g2_nand3_1 _14734_ (.B(net2727),
    .C(_09079_),
    .A(net245),
    .Y(_09080_));
 sg13g2_a21o_1 _14735_ (.A2(_09079_),
    .A1(net245),
    .B1(net2727),
    .X(_09081_));
 sg13g2_and2_1 _14736_ (.A(_09080_),
    .B(_09081_),
    .X(_00839_));
 sg13g2_nor2_1 _14737_ (.A(_05505_),
    .B(_09080_),
    .Y(_09082_));
 sg13g2_xnor2_1 _14738_ (.Y(_00840_),
    .A(net418),
    .B(_09080_));
 sg13g2_and2_1 _14739_ (.A(net368),
    .B(_09082_),
    .X(_09083_));
 sg13g2_xor2_1 _14740_ (.B(_09082_),
    .A(net368),
    .X(_00841_));
 sg13g2_xor2_1 _14741_ (.B(_09083_),
    .A(net303),
    .X(_00842_));
 sg13g2_nand3_1 _14742_ (.B(net2794),
    .C(_09083_),
    .A(net303),
    .Y(_09084_));
 sg13g2_a21o_1 _14743_ (.A2(_09083_),
    .A1(net303),
    .B1(net2794),
    .X(_09085_));
 sg13g2_and2_1 _14744_ (.A(_09084_),
    .B(_09085_),
    .X(_00843_));
 sg13g2_xnor2_1 _14745_ (.Y(_00844_),
    .A(net144),
    .B(_09084_));
 sg13g2_a21o_1 _14746_ (.A2(_06127_),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .B1(net334),
    .X(_00845_));
 sg13g2_nor2_1 _14747_ (.A(_05495_),
    .B(_08454_),
    .Y(_09086_));
 sg13g2_nor2_1 _14748_ (.A(_08455_),
    .B(_09086_),
    .Y(_09087_));
 sg13g2_nor2b_2 _14749_ (.A(net2862),
    .B_N(net5061),
    .Y(_09088_));
 sg13g2_nor2_2 _14750_ (.A(net5063),
    .B(net4221),
    .Y(_09089_));
 sg13g2_a22oi_1 _14751_ (.Y(_09090_),
    .B1(net4135),
    .B2(net9),
    .A2(net4686),
    .A1(net1927));
 sg13g2_nor2_1 _14752_ (.A(net2807),
    .B(net3882),
    .Y(_09091_));
 sg13g2_a21oi_1 _14753_ (.A1(net3882),
    .A2(_09090_),
    .Y(_00846_),
    .B1(_09091_));
 sg13g2_a22oi_1 _14754_ (.Y(_09092_),
    .B1(net4134),
    .B2(net10),
    .A2(net4688),
    .A1(net1954));
 sg13g2_nor2_1 _14755_ (.A(net2874),
    .B(net3890),
    .Y(_09093_));
 sg13g2_a21oi_1 _14756_ (.A1(net3888),
    .A2(_09092_),
    .Y(_00847_),
    .B1(_09093_));
 sg13g2_a22oi_1 _14757_ (.Y(_09094_),
    .B1(net4134),
    .B2(net11),
    .A2(net4689),
    .A1(net1750));
 sg13g2_nor2_1 _14758_ (.A(net2877),
    .B(net3888),
    .Y(_09095_));
 sg13g2_a21oi_1 _14759_ (.A1(net3888),
    .A2(_09094_),
    .Y(_00848_),
    .B1(_09095_));
 sg13g2_a22oi_1 _14760_ (.Y(_09096_),
    .B1(net4135),
    .B2(net12),
    .A2(net4686),
    .A1(net1848));
 sg13g2_nor2_1 _14761_ (.A(net2816),
    .B(net3882),
    .Y(_09097_));
 sg13g2_a21oi_1 _14762_ (.A1(net3883),
    .A2(_09096_),
    .Y(_00849_),
    .B1(_09097_));
 sg13g2_a22oi_1 _14763_ (.Y(_09098_),
    .B1(net4135),
    .B2(net1927),
    .A2(net4686),
    .A1(net2491));
 sg13g2_nor2_1 _14764_ (.A(net2635),
    .B(net3882),
    .Y(_09099_));
 sg13g2_a21oi_1 _14765_ (.A1(net3882),
    .A2(_09098_),
    .Y(_00850_),
    .B1(_09099_));
 sg13g2_a22oi_1 _14766_ (.Y(_09100_),
    .B1(net4134),
    .B2(net1954),
    .A2(net4689),
    .A1(net2543));
 sg13g2_nor2_1 _14767_ (.A(net2704),
    .B(net3888),
    .Y(_09101_));
 sg13g2_a21oi_1 _14768_ (.A1(net3888),
    .A2(_09100_),
    .Y(_00851_),
    .B1(_09101_));
 sg13g2_a22oi_1 _14769_ (.Y(_09102_),
    .B1(net4134),
    .B2(net1750),
    .A2(net4690),
    .A1(net1929));
 sg13g2_nor2_1 _14770_ (.A(net2820),
    .B(net3886),
    .Y(_09103_));
 sg13g2_a21oi_1 _14771_ (.A1(net3885),
    .A2(_09102_),
    .Y(_00852_),
    .B1(_09103_));
 sg13g2_a22oi_1 _14772_ (.Y(_09104_),
    .B1(net4135),
    .B2(net1848),
    .A2(net4687),
    .A1(net1967));
 sg13g2_nor2_1 _14773_ (.A(net2714),
    .B(net3884),
    .Y(_09105_));
 sg13g2_a21oi_1 _14774_ (.A1(net3883),
    .A2(_09104_),
    .Y(_00853_),
    .B1(_09105_));
 sg13g2_a22oi_1 _14775_ (.Y(_09106_),
    .B1(net4135),
    .B2(net2491),
    .A2(net4686),
    .A1(net1913));
 sg13g2_nor2_1 _14776_ (.A(net2788),
    .B(net3882),
    .Y(_09107_));
 sg13g2_a21oi_1 _14777_ (.A1(net3883),
    .A2(_09106_),
    .Y(_00854_),
    .B1(_09107_));
 sg13g2_a22oi_1 _14778_ (.Y(_09108_),
    .B1(net4134),
    .B2(net2543),
    .A2(net4689),
    .A1(net1836));
 sg13g2_nor2_1 _14779_ (.A(net2917),
    .B(net3885),
    .Y(_09109_));
 sg13g2_a21oi_1 _14780_ (.A1(net3886),
    .A2(_09108_),
    .Y(_00855_),
    .B1(_09109_));
 sg13g2_a22oi_1 _14781_ (.Y(_09110_),
    .B1(net4134),
    .B2(net1929),
    .A2(net4690),
    .A1(net2005));
 sg13g2_nor2_1 _14782_ (.A(net2669),
    .B(net3885),
    .Y(_09111_));
 sg13g2_a21oi_1 _14783_ (.A1(net3885),
    .A2(_09110_),
    .Y(_00856_),
    .B1(_09111_));
 sg13g2_a22oi_1 _14784_ (.Y(_09112_),
    .B1(net4134),
    .B2(net1967),
    .A2(net4687),
    .A1(net1865));
 sg13g2_nor2_1 _14785_ (.A(net2656),
    .B(net3884),
    .Y(_09113_));
 sg13g2_a21oi_1 _14786_ (.A1(net3884),
    .A2(_09112_),
    .Y(_00857_),
    .B1(_09113_));
 sg13g2_a22oi_1 _14787_ (.Y(_09114_),
    .B1(net4135),
    .B2(net1913),
    .A2(net4686),
    .A1(net1399));
 sg13g2_nor2_1 _14788_ (.A(net2553),
    .B(net3882),
    .Y(_09115_));
 sg13g2_a21oi_1 _14789_ (.A1(net3882),
    .A2(_09114_),
    .Y(_00858_),
    .B1(_09115_));
 sg13g2_a22oi_1 _14790_ (.Y(_09116_),
    .B1(_09089_),
    .B2(net1836),
    .A2(net4688),
    .A1(net1096));
 sg13g2_nor2_1 _14791_ (.A(net2856),
    .B(net3890),
    .Y(_09117_));
 sg13g2_a21oi_1 _14792_ (.A1(net3888),
    .A2(_09116_),
    .Y(_00859_),
    .B1(_09117_));
 sg13g2_a22oi_1 _14793_ (.Y(_09118_),
    .B1(net4134),
    .B2(net2005),
    .A2(net4690),
    .A1(net1499));
 sg13g2_nor2_1 _14794_ (.A(net2811),
    .B(net3886),
    .Y(_09119_));
 sg13g2_a21oi_1 _14795_ (.A1(net3886),
    .A2(_09118_),
    .Y(_00860_),
    .B1(_09119_));
 sg13g2_a22oi_1 _14796_ (.Y(_09120_),
    .B1(net4135),
    .B2(net1865),
    .A2(net4687),
    .A1(net1388));
 sg13g2_nor2_1 _14797_ (.A(net2693),
    .B(net3884),
    .Y(_09121_));
 sg13g2_a21oi_1 _14798_ (.A1(net3884),
    .A2(_09120_),
    .Y(_00861_),
    .B1(_09121_));
 sg13g2_nor2_1 _14799_ (.A(net9),
    .B(net4219),
    .Y(_09122_));
 sg13g2_nor2_1 _14800_ (.A(net1399),
    .B(net4221),
    .Y(_09123_));
 sg13g2_nor3_1 _14801_ (.A(net5061),
    .B(_09122_),
    .C(_09123_),
    .Y(_09124_));
 sg13g2_a21oi_1 _14802_ (.A1(net1719),
    .A2(net4686),
    .Y(_09125_),
    .B1(_09124_));
 sg13g2_nor2_1 _14803_ (.A(net2677),
    .B(net3884),
    .Y(_09126_));
 sg13g2_a21oi_1 _14804_ (.A1(net3883),
    .A2(_09125_),
    .Y(_00862_),
    .B1(_09126_));
 sg13g2_nor2_1 _14805_ (.A(net10),
    .B(net4218),
    .Y(_09127_));
 sg13g2_nor2_1 _14806_ (.A(net1096),
    .B(net4220),
    .Y(_09128_));
 sg13g2_nor3_1 _14807_ (.A(net5062),
    .B(_09127_),
    .C(_09128_),
    .Y(_09129_));
 sg13g2_a21oi_1 _14808_ (.A1(net1859),
    .A2(net4688),
    .Y(_09130_),
    .B1(_09129_));
 sg13g2_nor2_1 _14809_ (.A(net2611),
    .B(net3891),
    .Y(_09131_));
 sg13g2_a21oi_1 _14810_ (.A1(net3889),
    .A2(_09130_),
    .Y(_00863_),
    .B1(_09131_));
 sg13g2_nor2_1 _14811_ (.A(net11),
    .B(net4218),
    .Y(_09132_));
 sg13g2_nor2_1 _14812_ (.A(net1499),
    .B(net4220),
    .Y(_09133_));
 sg13g2_nor3_1 _14813_ (.A(net5062),
    .B(_09132_),
    .C(_09133_),
    .Y(_09134_));
 sg13g2_a21oi_1 _14814_ (.A1(net1600),
    .A2(net4689),
    .Y(_09135_),
    .B1(_09134_));
 sg13g2_nor2_1 _14815_ (.A(net2647),
    .B(net3885),
    .Y(_09136_));
 sg13g2_a21oi_1 _14816_ (.A1(net3885),
    .A2(_09135_),
    .Y(_00864_),
    .B1(_09136_));
 sg13g2_nor2_1 _14817_ (.A(net12),
    .B(net4219),
    .Y(_09137_));
 sg13g2_nor2_1 _14818_ (.A(net1388),
    .B(net4221),
    .Y(_09138_));
 sg13g2_nor3_1 _14819_ (.A(net5063),
    .B(_09137_),
    .C(_09138_),
    .Y(_09139_));
 sg13g2_a21oi_1 _14820_ (.A1(net1341),
    .A2(net4687),
    .Y(_09140_),
    .B1(_09139_));
 sg13g2_nor2_1 _14821_ (.A(net2881),
    .B(net3887),
    .Y(_09141_));
 sg13g2_a21oi_1 _14822_ (.A1(net3887),
    .A2(_09140_),
    .Y(_00865_),
    .B1(_09141_));
 sg13g2_nor2_1 _14823_ (.A(net1927),
    .B(net4219),
    .Y(_09142_));
 sg13g2_nor2_1 _14824_ (.A(net1719),
    .B(net4221),
    .Y(_09143_));
 sg13g2_nor3_1 _14825_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(_09142_),
    .C(_09143_),
    .Y(_09144_));
 sg13g2_a21oi_1 _14826_ (.A1(net1846),
    .A2(net4686),
    .Y(_09145_),
    .B1(_09144_));
 sg13g2_nor2_1 _14827_ (.A(net2848),
    .B(net3890),
    .Y(_09146_));
 sg13g2_a21oi_1 _14828_ (.A1(net3890),
    .A2(_09145_),
    .Y(_00866_),
    .B1(_09146_));
 sg13g2_nor2_1 _14829_ (.A(net1954),
    .B(net4218),
    .Y(_09147_));
 sg13g2_nor2_1 _14830_ (.A(net1859),
    .B(net4220),
    .Y(_09148_));
 sg13g2_nor3_1 _14831_ (.A(net5062),
    .B(_09147_),
    .C(_09148_),
    .Y(_09149_));
 sg13g2_a21oi_1 _14832_ (.A1(net2040),
    .A2(net4688),
    .Y(_09150_),
    .B1(_09149_));
 sg13g2_nor2_1 _14833_ (.A(net2564),
    .B(net3889),
    .Y(_09151_));
 sg13g2_a21oi_1 _14834_ (.A1(net3891),
    .A2(_09150_),
    .Y(_00867_),
    .B1(_09151_));
 sg13g2_nor2_1 _14835_ (.A(net1750),
    .B(net4218),
    .Y(_09152_));
 sg13g2_nor2_1 _14836_ (.A(net1600),
    .B(net4220),
    .Y(_09153_));
 sg13g2_nor3_1 _14837_ (.A(net5062),
    .B(_09152_),
    .C(_09153_),
    .Y(_09154_));
 sg13g2_a21oi_1 _14838_ (.A1(net1514),
    .A2(net4688),
    .Y(_09155_),
    .B1(_09154_));
 sg13g2_nor2_1 _14839_ (.A(net2565),
    .B(net3890),
    .Y(_09156_));
 sg13g2_a21oi_1 _14840_ (.A1(net3889),
    .A2(_09155_),
    .Y(_00868_),
    .B1(_09156_));
 sg13g2_nor2_1 _14841_ (.A(net1848),
    .B(net4219),
    .Y(_09157_));
 sg13g2_nor2_1 _14842_ (.A(net1341),
    .B(net4221),
    .Y(_09158_));
 sg13g2_nor3_1 _14843_ (.A(net5063),
    .B(_09157_),
    .C(_09158_),
    .Y(_09159_));
 sg13g2_a21oi_1 _14844_ (.A1(net953),
    .A2(net4687),
    .Y(_09160_),
    .B1(_09159_));
 sg13g2_nor2_1 _14845_ (.A(net2666),
    .B(net3884),
    .Y(_09161_));
 sg13g2_a21oi_1 _14846_ (.A1(net3892),
    .A2(_09160_),
    .Y(_00869_),
    .B1(_09161_));
 sg13g2_nor2_1 _14847_ (.A(net1846),
    .B(net4221),
    .Y(_09162_));
 sg13g2_nor3_1 _14848_ (.A(net5063),
    .B(_08388_),
    .C(_09162_),
    .Y(_09163_));
 sg13g2_a21oi_1 _14849_ (.A1(net2903),
    .A2(net4687),
    .Y(_09164_),
    .B1(_09163_));
 sg13g2_nor2_1 _14850_ (.A(net2879),
    .B(net3887),
    .Y(_09165_));
 sg13g2_a21oi_1 _14851_ (.A1(net3885),
    .A2(net2904),
    .Y(_00870_),
    .B1(_09165_));
 sg13g2_nor2_1 _14852_ (.A(net2040),
    .B(_08386_),
    .Y(_09166_));
 sg13g2_nor3_1 _14853_ (.A(net5063),
    .B(_08391_),
    .C(_09166_),
    .Y(_09167_));
 sg13g2_a21oi_1 _14854_ (.A1(net1723),
    .A2(net4688),
    .Y(_09168_),
    .B1(_09167_));
 sg13g2_nor2_1 _14855_ (.A(net2641),
    .B(net3889),
    .Y(_09169_));
 sg13g2_a21oi_1 _14856_ (.A1(net3889),
    .A2(_09168_),
    .Y(_00871_),
    .B1(_09169_));
 sg13g2_nor2_1 _14857_ (.A(net1929),
    .B(net4218),
    .Y(_09170_));
 sg13g2_nor2_1 _14858_ (.A(net1514),
    .B(_08386_),
    .Y(_09171_));
 sg13g2_nor3_1 _14859_ (.A(net5062),
    .B(_09170_),
    .C(_09171_),
    .Y(_09172_));
 sg13g2_a21oi_1 _14860_ (.A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ),
    .A2(net4688),
    .Y(_09173_),
    .B1(_09172_));
 sg13g2_nor2_1 _14861_ (.A(net2072),
    .B(net3888),
    .Y(_09174_));
 sg13g2_a21oi_1 _14862_ (.A1(net3891),
    .A2(_09173_),
    .Y(_00872_),
    .B1(_09174_));
 sg13g2_nor2_1 _14863_ (.A(net1967),
    .B(net4218),
    .Y(_09175_));
 sg13g2_nor2_1 _14864_ (.A(net953),
    .B(net4220),
    .Y(_09176_));
 sg13g2_nor3_1 _14865_ (.A(net5062),
    .B(_09175_),
    .C(_09176_),
    .Y(_09177_));
 sg13g2_a21oi_1 _14866_ (.A1(net2840),
    .A2(net4690),
    .Y(_09178_),
    .B1(_09177_));
 sg13g2_nor2_1 _14867_ (.A(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .B(net3890),
    .Y(_09179_));
 sg13g2_a21oi_1 _14868_ (.A1(net3886),
    .A2(net2841),
    .Y(_00873_),
    .B1(_09179_));
 sg13g2_nor2_1 _14869_ (.A(net1913),
    .B(net4219),
    .Y(_09180_));
 sg13g2_nor2_1 _14870_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ),
    .B(net4221),
    .Y(_09181_));
 sg13g2_nor3_1 _14871_ (.A(net5063),
    .B(_09180_),
    .C(_09181_),
    .Y(_09182_));
 sg13g2_a21oi_1 _14872_ (.A1(net866),
    .A2(net4686),
    .Y(_09183_),
    .B1(_09182_));
 sg13g2_nor2_1 _14873_ (.A(net2615),
    .B(net3885),
    .Y(_09184_));
 sg13g2_a21oi_1 _14874_ (.A1(net3884),
    .A2(_09183_),
    .Y(_00874_),
    .B1(_09184_));
 sg13g2_nor2_1 _14875_ (.A(net1836),
    .B(_08387_),
    .Y(_09185_));
 sg13g2_nor2_1 _14876_ (.A(net1723),
    .B(net4220),
    .Y(_09186_));
 sg13g2_nor3_1 _14877_ (.A(net5063),
    .B(_09185_),
    .C(_09186_),
    .Y(_09187_));
 sg13g2_a21oi_1 _14878_ (.A1(net2462),
    .A2(net4689),
    .Y(_09188_),
    .B1(_09187_));
 sg13g2_nor2_1 _14879_ (.A(\soc_inst.mem_ctrl.spi_data_out[29] ),
    .B(net3889),
    .Y(_09189_));
 sg13g2_a21oi_1 _14880_ (.A1(net3888),
    .A2(net2463),
    .Y(_00875_),
    .B1(_09189_));
 sg13g2_nor2_1 _14881_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ),
    .B(_08387_),
    .Y(_09190_));
 sg13g2_nor2_1 _14882_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ),
    .B(net4220),
    .Y(_09191_));
 sg13g2_nor3_1 _14883_ (.A(net5062),
    .B(_09190_),
    .C(_09191_),
    .Y(_09192_));
 sg13g2_a21oi_1 _14884_ (.A1(net1046),
    .A2(net4688),
    .Y(_09193_),
    .B1(_09192_));
 sg13g2_nor2_1 _14885_ (.A(net2000),
    .B(net3890),
    .Y(_09194_));
 sg13g2_a21oi_1 _14886_ (.A1(net3889),
    .A2(_09193_),
    .Y(_00876_),
    .B1(_09194_));
 sg13g2_nor2_1 _14887_ (.A(net1865),
    .B(net4218),
    .Y(_09195_));
 sg13g2_nor2_1 _14888_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ),
    .B(net4220),
    .Y(_09196_));
 sg13g2_nor3_1 _14889_ (.A(net5062),
    .B(_09195_),
    .C(_09196_),
    .Y(_09197_));
 sg13g2_a21oi_1 _14890_ (.A1(net970),
    .A2(net4690),
    .Y(_09198_),
    .B1(_09197_));
 sg13g2_nor2_1 _14891_ (.A(net2097),
    .B(net3889),
    .Y(_09199_));
 sg13g2_a21oi_1 _14892_ (.A1(net3891),
    .A2(_09198_),
    .Y(_00877_),
    .B1(_09199_));
 sg13g2_nand2_2 _14893_ (.Y(_09200_),
    .A(\soc_inst.cpu_core.csr_file.mie[11] ),
    .B(\soc_inst.cpu_core.csr_file.mip_eip ));
 sg13g2_nand4_1 _14894_ (.B(\soc_inst.cpu_core.if_pc[5] ),
    .C(\soc_inst.cpu_core.if_pc[6] ),
    .A(\soc_inst.cpu_core.if_pc[4] ),
    .Y(_09201_),
    .D(\soc_inst.cpu_core.if_pc[7] ));
 sg13g2_nand3_1 _14895_ (.B(\soc_inst.cpu_core.if_pc[0] ),
    .C(\soc_inst.cpu_core.if_pc[3] ),
    .A(\soc_inst.cpu_core.if_pc[1] ),
    .Y(_09202_));
 sg13g2_nor3_1 _14896_ (.A(_05522_),
    .B(_09201_),
    .C(_09202_),
    .Y(_09203_));
 sg13g2_nand4_1 _14897_ (.B(\soc_inst.cpu_core.if_pc[13] ),
    .C(\soc_inst.cpu_core.if_pc[14] ),
    .A(\soc_inst.cpu_core.if_pc[12] ),
    .Y(_09204_),
    .D(\soc_inst.cpu_core.if_pc[15] ));
 sg13g2_nand4_1 _14898_ (.B(\soc_inst.cpu_core.if_pc[9] ),
    .C(\soc_inst.cpu_core.if_pc[10] ),
    .A(\soc_inst.cpu_core.if_pc[8] ),
    .Y(_09205_),
    .D(\soc_inst.cpu_core.if_pc[11] ));
 sg13g2_nand4_1 _14899_ (.B(\soc_inst.cpu_core.if_pc[17] ),
    .C(\soc_inst.cpu_core.if_pc[18] ),
    .A(\soc_inst.cpu_core.if_pc[16] ),
    .Y(_09206_),
    .D(\soc_inst.cpu_core.if_pc[19] ));
 sg13g2_nand4_1 _14900_ (.B(\soc_inst.cpu_core.if_pc[21] ),
    .C(\soc_inst.cpu_core.if_pc[22] ),
    .A(\soc_inst.cpu_core.if_pc[20] ),
    .Y(_09207_),
    .D(\soc_inst.cpu_core.if_pc[23] ));
 sg13g2_nor4_1 _14901_ (.A(_09204_),
    .B(_09205_),
    .C(_09206_),
    .D(_09207_),
    .Y(_09208_));
 sg13g2_a221oi_1 _14902_ (.B2(_09208_),
    .C1(_05518_),
    .B1(_09203_),
    .A1(_06805_),
    .Y(_09209_),
    .A2(_09200_));
 sg13g2_nor2_1 _14903_ (.A(net4972),
    .B(_09209_),
    .Y(_09210_));
 sg13g2_or2_1 _14904_ (.X(_09211_),
    .B(_09209_),
    .A(net4903));
 sg13g2_a21oi_1 _14905_ (.A1(_05479_),
    .A2(net4960),
    .Y(_00878_),
    .B1(net4129));
 sg13g2_nand2_2 _14906_ (.Y(_09212_),
    .A(net4752),
    .B(net541));
 sg13g2_nor2_1 _14907_ (.A(_00268_),
    .B(_00267_),
    .Y(_09213_));
 sg13g2_nand2_2 _14908_ (.Y(_09214_),
    .A(_00269_),
    .B(_09213_));
 sg13g2_nor3_2 _14909_ (.A(\soc_inst.cpu_core.id_instr[3] ),
    .B(\soc_inst.cpu_core.id_instr[2] ),
    .C(_09214_),
    .Y(_09215_));
 sg13g2_nor2b_1 _14910_ (.A(net4878),
    .B_N(_09215_),
    .Y(_09216_));
 sg13g2_nand2b_1 _14911_ (.Y(_09217_),
    .B(_09215_),
    .A_N(net4878));
 sg13g2_o21ai_1 _14912_ (.B1(_09212_),
    .Y(_09218_),
    .A1(net4970),
    .A2(_09216_));
 sg13g2_nor4_1 _14913_ (.A(\soc_inst.cpu_core.id_instr[8] ),
    .B(\soc_inst.cpu_core.id_instr[7] ),
    .C(\soc_inst.cpu_core.id_instr[10] ),
    .D(\soc_inst.cpu_core.id_instr[11] ),
    .Y(_09219_));
 sg13g2_nor2b_2 _14914_ (.A(\soc_inst.cpu_core.id_instr[9] ),
    .B_N(_09219_),
    .Y(_09220_));
 sg13g2_nor4_1 _14915_ (.A(_00269_),
    .B(_00268_),
    .C(_00267_),
    .D(\soc_inst.cpu_core.id_instr[3] ),
    .Y(_09221_));
 sg13g2_nand4_1 _14916_ (.B(net541),
    .C(net4878),
    .A(_05517_),
    .Y(_09222_),
    .D(_09221_));
 sg13g2_nor2_1 _14917_ (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[1] ),
    .Y(_09223_));
 sg13g2_nor3_2 _14918_ (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[0] ),
    .C(\soc_inst.cpu_core.id_funct3[1] ),
    .Y(_09224_));
 sg13g2_nor3_1 _14919_ (.A(_09220_),
    .B(_09222_),
    .C(_09224_),
    .Y(_09225_));
 sg13g2_nand3_1 _14920_ (.B(\soc_inst.cpu_core.id_instr[5] ),
    .C(net4878),
    .A(\soc_inst.cpu_core.id_instr[2] ),
    .Y(_09226_));
 sg13g2_nor2_2 _14921_ (.A(_09214_),
    .B(_09226_),
    .Y(_09227_));
 sg13g2_nor2b_1 _14922_ (.A(net4878),
    .B_N(_09221_),
    .Y(_09228_));
 sg13g2_nor3_1 _14923_ (.A(\soc_inst.cpu_core.id_instr[3] ),
    .B(_09214_),
    .C(_09226_),
    .Y(_09229_));
 sg13g2_nand2b_2 _14924_ (.Y(_09230_),
    .B(_09227_),
    .A_N(\soc_inst.cpu_core.id_instr[3] ));
 sg13g2_and2_1 _14925_ (.A(\soc_inst.cpu_core.id_instr[3] ),
    .B(_09227_),
    .X(_09231_));
 sg13g2_nand2_2 _14926_ (.Y(_09232_),
    .A(\soc_inst.cpu_core.id_instr[3] ),
    .B(_09227_));
 sg13g2_nor3_1 _14927_ (.A(_09225_),
    .B(_09227_),
    .C(_09228_),
    .Y(_09233_));
 sg13g2_a22oi_1 _14928_ (.Y(_00879_),
    .B1(_09218_),
    .B2(_09233_),
    .A2(_05543_),
    .A1(net4970));
 sg13g2_nand2_1 _14929_ (.Y(_09234_),
    .A(net5051),
    .B(net4964));
 sg13g2_nor4_1 _14930_ (.A(net720),
    .B(net2354),
    .C(net2358),
    .D(net2139),
    .Y(_09235_));
 sg13g2_nor2_1 _14931_ (.A(net2505),
    .B(net583),
    .Y(_09236_));
 sg13g2_and2_1 _14932_ (.A(net2631),
    .B(net567),
    .X(_09237_));
 sg13g2_nand4_1 _14933_ (.B(_09235_),
    .C(_09236_),
    .A(net2307),
    .Y(_09238_),
    .D(_09237_));
 sg13g2_nor2_1 _14934_ (.A(net4956),
    .B(\soc_inst.cpu_core.id_imm12[3] ),
    .Y(_09239_));
 sg13g2_nor2b_2 _14935_ (.A(_09222_),
    .B_N(_09224_),
    .Y(_09240_));
 sg13g2_nor4_1 _14936_ (.A(net4955),
    .B(net2702),
    .C(net2585),
    .D(net2330),
    .Y(_09241_));
 sg13g2_nand2_1 _14937_ (.Y(_09242_),
    .A(_09240_),
    .B(_09241_));
 sg13g2_o21ai_1 _14938_ (.B1(_09234_),
    .Y(_00880_),
    .A1(_09238_),
    .A2(_09242_));
 sg13g2_nor3_1 _14939_ (.A(\soc_inst.cpu_core.id_imm12[1] ),
    .B(\soc_inst.cpu_core.id_imm12[8] ),
    .C(net567),
    .Y(_09243_));
 sg13g2_nand3_1 _14940_ (.B(_09236_),
    .C(_09243_),
    .A(_09235_),
    .Y(_09244_));
 sg13g2_nand2_1 _14941_ (.Y(_09245_),
    .A(\soc_inst.cpu_core.id_imm12[0] ),
    .B(_09239_));
 sg13g2_nor3_1 _14942_ (.A(\soc_inst.cpu_core.id_imm12[2] ),
    .B(_09244_),
    .C(_09245_),
    .Y(_09246_));
 sg13g2_a22oi_1 _14943_ (.Y(_09247_),
    .B1(_09240_),
    .B2(_09246_),
    .A2(net4960),
    .A1(net1911));
 sg13g2_inv_1 _14944_ (.Y(_00881_),
    .A(net1912));
 sg13g2_mux2_1 _14945_ (.A0(net336),
    .A1(net5050),
    .S(net4978),
    .X(_00882_));
 sg13g2_mux2_1 _14946_ (.A0(net896),
    .A1(\soc_inst.core_mem_wdata[1] ),
    .S(net4934),
    .X(_00883_));
 sg13g2_mux2_1 _14947_ (.A0(net1265),
    .A1(\soc_inst.core_mem_wdata[2] ),
    .S(net4979),
    .X(_00884_));
 sg13g2_mux2_1 _14948_ (.A0(net783),
    .A1(\soc_inst.core_mem_wdata[3] ),
    .S(net4947),
    .X(_00885_));
 sg13g2_mux2_1 _14949_ (.A0(net399),
    .A1(net957),
    .S(net4947),
    .X(_00886_));
 sg13g2_mux2_1 _14950_ (.A0(net364),
    .A1(net1023),
    .S(net4947),
    .X(_00887_));
 sg13g2_mux2_1 _14951_ (.A0(net1147),
    .A1(\soc_inst.core_mem_wdata[6] ),
    .S(net4979),
    .X(_00888_));
 sg13g2_mux2_1 _14952_ (.A0(net1201),
    .A1(net5030),
    .S(net4978),
    .X(_00889_));
 sg13g2_mux2_1 _14953_ (.A0(net707),
    .A1(net5027),
    .S(net4985),
    .X(_00890_));
 sg13g2_mux2_1 _14954_ (.A0(net940),
    .A1(net5025),
    .S(net4979),
    .X(_00891_));
 sg13g2_mux2_1 _14955_ (.A0(net717),
    .A1(net5023),
    .S(net4985),
    .X(_00892_));
 sg13g2_mux2_1 _14956_ (.A0(net1476),
    .A1(net5022),
    .S(net4979),
    .X(_00893_));
 sg13g2_mux2_1 _14957_ (.A0(net1102),
    .A1(net5021),
    .S(net4979),
    .X(_00894_));
 sg13g2_mux2_1 _14958_ (.A0(net2162),
    .A1(net5020),
    .S(net4922),
    .X(_00895_));
 sg13g2_mux2_1 _14959_ (.A0(net1293),
    .A1(net5019),
    .S(net4962),
    .X(_00896_));
 sg13g2_mux2_1 _14960_ (.A0(net372),
    .A1(net5018),
    .S(net4946),
    .X(_00897_));
 sg13g2_mux2_1 _14961_ (.A0(net1066),
    .A1(\soc_inst.core_mem_wdata[16] ),
    .S(net4989),
    .X(_00898_));
 sg13g2_mux2_1 _14962_ (.A0(net2870),
    .A1(\soc_inst.core_mem_wdata[17] ),
    .S(net4991),
    .X(_00899_));
 sg13g2_mux2_1 _14963_ (.A0(net1085),
    .A1(net1170),
    .S(net4989),
    .X(_00900_));
 sg13g2_mux2_1 _14964_ (.A0(net311),
    .A1(net1021),
    .S(net4995),
    .X(_00901_));
 sg13g2_mux2_1 _14965_ (.A0(net2851),
    .A1(\soc_inst.core_mem_wdata[20] ),
    .S(net4991),
    .X(_00902_));
 sg13g2_mux2_1 _14966_ (.A0(net1174),
    .A1(\soc_inst.core_mem_wdata[21] ),
    .S(net4989),
    .X(_00903_));
 sg13g2_mux2_1 _14967_ (.A0(\soc_inst.cpu_core.ex_rs2_data[22] ),
    .A1(net2754),
    .S(net4995),
    .X(_00904_));
 sg13g2_mux2_1 _14968_ (.A0(net1972),
    .A1(net2758),
    .S(net4989),
    .X(_00905_));
 sg13g2_mux2_1 _14969_ (.A0(net497),
    .A1(net962),
    .S(net4979),
    .X(_00906_));
 sg13g2_mux2_1 _14970_ (.A0(net1172),
    .A1(\soc_inst.core_mem_wdata[25] ),
    .S(net4981),
    .X(_00907_));
 sg13g2_mux2_1 _14971_ (.A0(net2397),
    .A1(net532),
    .S(net4995),
    .X(_00908_));
 sg13g2_mux2_1 _14972_ (.A0(net316),
    .A1(net480),
    .S(net4995),
    .X(_00909_));
 sg13g2_mux2_1 _14973_ (.A0(net1874),
    .A1(net610),
    .S(net4996),
    .X(_00910_));
 sg13g2_mux2_1 _14974_ (.A0(net713),
    .A1(\soc_inst.core_mem_wdata[29] ),
    .S(net4940),
    .X(_00911_));
 sg13g2_mux2_1 _14975_ (.A0(net2466),
    .A1(net383),
    .S(net4995),
    .X(_00912_));
 sg13g2_mux2_1 _14976_ (.A0(net863),
    .A1(net422),
    .S(net4995),
    .X(_00913_));
 sg13g2_nand2_1 _14977_ (.Y(_09248_),
    .A(net574),
    .B(net4960));
 sg13g2_o21ai_1 _14978_ (.B1(_09248_),
    .Y(_00914_),
    .A1(_09242_),
    .A2(_09244_));
 sg13g2_a21o_1 _14979_ (.A2(net4059),
    .A1(net4749),
    .B1(net525),
    .X(_00915_));
 sg13g2_and2_1 _14980_ (.A(_08779_),
    .B(_08781_),
    .X(_09249_));
 sg13g2_nand2_2 _14981_ (.Y(_09250_),
    .A(_08779_),
    .B(_08781_));
 sg13g2_nor3_1 _14982_ (.A(net5114),
    .B(net4031),
    .C(net3720),
    .Y(_09251_));
 sg13g2_a21o_1 _14983_ (.A2(net4943),
    .A1(net1676),
    .B1(_09251_),
    .X(_00916_));
 sg13g2_nor3_1 _14984_ (.A(net5113),
    .B(_08817_),
    .C(net3720),
    .Y(_09252_));
 sg13g2_a21o_1 _14985_ (.A2(net4934),
    .A1(net1426),
    .B1(_09252_),
    .X(_00917_));
 sg13g2_nor2b_1 _14986_ (.A(net5084),
    .B_N(net5086),
    .Y(_09253_));
 sg13g2_nand2b_2 _14987_ (.Y(_09254_),
    .B(net5087),
    .A_N(net5085));
 sg13g2_nand2_1 _14988_ (.Y(_09255_),
    .A(net5099),
    .B(_08790_));
 sg13g2_nor2_1 _14989_ (.A(net4601),
    .B(net4595),
    .Y(_09256_));
 sg13g2_o21ai_1 _14990_ (.B1(_08800_),
    .Y(_09257_),
    .A1(net4602),
    .A2(_09255_));
 sg13g2_o21ai_1 _14991_ (.B1(_09257_),
    .Y(_09258_),
    .A1(net5082),
    .A2(_09254_));
 sg13g2_nand3_1 _14992_ (.B(_09254_),
    .C(_09257_),
    .A(_08813_),
    .Y(_09259_));
 sg13g2_nand2_1 _14993_ (.Y(_09260_),
    .A(_08803_),
    .B(net4599));
 sg13g2_inv_1 _14994_ (.Y(_09261_),
    .A(_09260_));
 sg13g2_a21oi_1 _14995_ (.A1(\soc_inst.core_instr_data[12] ),
    .A2(_08793_),
    .Y(_09262_),
    .B1(_09260_));
 sg13g2_nand2b_1 _14996_ (.Y(_09263_),
    .B(_08822_),
    .A_N(_09262_));
 sg13g2_a21oi_1 _14997_ (.A1(_08822_),
    .A2(_09260_),
    .Y(_09264_),
    .B1(net4691));
 sg13g2_a22oi_1 _14998_ (.Y(_09265_),
    .B1(_09263_),
    .B2(_08818_),
    .A2(_09259_),
    .A1(net4695));
 sg13g2_nor2_1 _14999_ (.A(net5112),
    .B(net4028),
    .Y(_09266_));
 sg13g2_a21oi_1 _15000_ (.A1(net4030),
    .A2(_09265_),
    .Y(_09267_),
    .B1(_09266_));
 sg13g2_a22oi_1 _15001_ (.Y(_09268_),
    .B1(net3722),
    .B2(_09267_),
    .A2(net2580),
    .A1(net4934));
 sg13g2_inv_1 _15002_ (.Y(_00918_),
    .A(_09268_));
 sg13g2_nand2_1 _15003_ (.Y(_09269_),
    .A(net5110),
    .B(net4032));
 sg13g2_o21ai_1 _15004_ (.B1(_09269_),
    .Y(_09270_),
    .A1(net4033),
    .A2(_09254_));
 sg13g2_a22oi_1 _15005_ (.Y(_09271_),
    .B1(net3723),
    .B2(_09270_),
    .A2(net2798),
    .A1(net4934));
 sg13g2_inv_1 _15006_ (.Y(_00919_),
    .A(_09271_));
 sg13g2_nor2_2 _15007_ (.A(net4696),
    .B(_08788_),
    .Y(_09272_));
 sg13g2_and2_1 _15008_ (.A(net5085),
    .B(net5083),
    .X(_09273_));
 sg13g2_nand2_1 _15009_ (.Y(_09274_),
    .A(net5084),
    .B(net5083));
 sg13g2_nor2_1 _15010_ (.A(net4684),
    .B(net4683),
    .Y(_09275_));
 sg13g2_nor3_2 _15011_ (.A(net5088),
    .B(net5085),
    .C(net5083),
    .Y(_09276_));
 sg13g2_nand2_1 _15012_ (.Y(_09277_),
    .A(_05648_),
    .B(_08807_));
 sg13g2_nor2_1 _15013_ (.A(_08803_),
    .B(_08809_),
    .Y(_09278_));
 sg13g2_o21ai_1 _15014_ (.B1(net4599),
    .Y(_09279_),
    .A1(_08793_),
    .A2(_08804_));
 sg13g2_nand3_1 _15015_ (.B(net4594),
    .C(_09279_),
    .A(_08822_),
    .Y(_09280_));
 sg13g2_a221oi_1 _15016_ (.B2(net4692),
    .C1(_09272_),
    .B1(_09280_),
    .A1(net4694),
    .Y(_09281_),
    .A2(_09275_));
 sg13g2_nor2_1 _15017_ (.A(net4032),
    .B(_09281_),
    .Y(_09282_));
 sg13g2_a21oi_1 _15018_ (.A1(net5108),
    .A2(net4033),
    .Y(_09283_),
    .B1(_09282_));
 sg13g2_a22oi_1 _15019_ (.Y(_09284_),
    .B1(net3722),
    .B2(_09283_),
    .A2(net4934),
    .A1(net5017));
 sg13g2_inv_1 _15020_ (.Y(_00920_),
    .A(_09284_));
 sg13g2_nor2_1 _15021_ (.A(net5106),
    .B(net4025),
    .Y(_09285_));
 sg13g2_nand3_1 _15022_ (.B(_08810_),
    .C(_08819_),
    .A(_08807_),
    .Y(_09286_));
 sg13g2_a221oi_1 _15023_ (.B2(net5083),
    .C1(_09258_),
    .B1(_09286_),
    .A1(net4692),
    .Y(_09287_),
    .A2(_08823_));
 sg13g2_a21oi_1 _15024_ (.A1(net4028),
    .A2(_09287_),
    .Y(_09288_),
    .B1(_09285_));
 sg13g2_a22oi_1 _15025_ (.Y(_09289_),
    .B1(net3722),
    .B2(_09288_),
    .A2(net2608),
    .A1(net4950));
 sg13g2_inv_1 _15026_ (.Y(_00921_),
    .A(_09289_));
 sg13g2_nand2_1 _15027_ (.Y(_09290_),
    .A(net5104),
    .B(net4035));
 sg13g2_o21ai_1 _15028_ (.B1(_08806_),
    .Y(_09291_),
    .A1(net5082),
    .A2(_09254_));
 sg13g2_nand4_1 _15029_ (.B(_08813_),
    .C(_09254_),
    .A(_08806_),
    .Y(_09292_),
    .D(_09274_));
 sg13g2_a21oi_1 _15030_ (.A1(net4695),
    .A2(_09292_),
    .Y(_09293_),
    .B1(_09264_));
 sg13g2_o21ai_1 _15031_ (.B1(_09290_),
    .Y(_09294_),
    .A1(net4035),
    .A2(_09293_));
 sg13g2_a22oi_1 _15032_ (.Y(_09295_),
    .B1(net3729),
    .B2(_09294_),
    .A2(net5016),
    .A1(net4936));
 sg13g2_inv_1 _15033_ (.Y(_00922_),
    .A(_09295_));
 sg13g2_nand2_1 _15034_ (.Y(_09296_),
    .A(net4927),
    .B(net905));
 sg13g2_o21ai_1 _15035_ (.B1(net4692),
    .Y(_09297_),
    .A1(net4598),
    .A2(_09278_));
 sg13g2_nand2_1 _15036_ (.Y(_09298_),
    .A(net4028),
    .B(_09297_));
 sg13g2_a21oi_1 _15037_ (.A1(net5111),
    .A2(_08789_),
    .Y(_09299_),
    .B1(net4137));
 sg13g2_a21oi_1 _15038_ (.A1(net5103),
    .A2(_09276_),
    .Y(_09300_),
    .B1(_08823_));
 sg13g2_o21ai_1 _15039_ (.B1(_09262_),
    .Y(_09301_),
    .A1(net5091),
    .A2(_08793_));
 sg13g2_a21oi_1 _15040_ (.A1(_09300_),
    .A2(_09301_),
    .Y(_09302_),
    .B1(net4691));
 sg13g2_nand2_1 _15041_ (.Y(_09303_),
    .A(net5102),
    .B(net4599));
 sg13g2_a22oi_1 _15042_ (.Y(_09304_),
    .B1(net4682),
    .B2(net5091),
    .A2(_08798_),
    .A1(net5102));
 sg13g2_nand4_1 _15043_ (.B(net4594),
    .C(_09303_),
    .A(_08813_),
    .Y(_09305_),
    .D(_09304_));
 sg13g2_nor2_2 _15044_ (.A(_08815_),
    .B(_09276_),
    .Y(_09306_));
 sg13g2_inv_2 _15045_ (.Y(_09307_),
    .A(_09306_));
 sg13g2_a21o_1 _15046_ (.A2(net4694),
    .A1(net5103),
    .B1(_09306_),
    .X(_09308_));
 sg13g2_o21ai_1 _15047_ (.B1(_09308_),
    .Y(_09309_),
    .A1(_09291_),
    .A2(_09305_));
 sg13g2_o21ai_1 _15048_ (.B1(_09309_),
    .Y(_09310_),
    .A1(net4696),
    .A2(_09299_));
 sg13g2_or2_1 _15049_ (.X(_09311_),
    .B(_09310_),
    .A(_09302_));
 sg13g2_a22oi_1 _15050_ (.Y(_09312_),
    .B1(_09311_),
    .B2(net4028),
    .A2(_09298_),
    .A1(net5103));
 sg13g2_o21ai_1 _15051_ (.B1(_09296_),
    .Y(_00923_),
    .A1(net3721),
    .A2(_09312_));
 sg13g2_nand2_1 _15052_ (.Y(_09313_),
    .A(net4932),
    .B(net568));
 sg13g2_a21oi_1 _15053_ (.A1(net5110),
    .A2(_08789_),
    .Y(_09314_),
    .B1(net4137));
 sg13g2_nor2_2 _15054_ (.A(net4691),
    .B(_08827_),
    .Y(_09315_));
 sg13g2_a21o_1 _15055_ (.A2(net4694),
    .A1(net5099),
    .B1(_09306_),
    .X(_09316_));
 sg13g2_nand2_1 _15056_ (.Y(_09317_),
    .A(_08806_),
    .B(net4594));
 sg13g2_a21oi_1 _15057_ (.A1(net5100),
    .A2(net4599),
    .Y(_09318_),
    .B1(_08812_));
 sg13g2_a22oi_1 _15058_ (.Y(_09319_),
    .B1(net4682),
    .B2(\soc_inst.core_instr_data[3] ),
    .A2(_08800_),
    .A1(net5100));
 sg13g2_nand4_1 _15059_ (.B(net4594),
    .C(_09318_),
    .A(_08806_),
    .Y(_09320_),
    .D(_09319_));
 sg13g2_a21oi_1 _15060_ (.A1(_09316_),
    .A2(_09320_),
    .Y(_09321_),
    .B1(_09315_));
 sg13g2_o21ai_1 _15061_ (.B1(_09321_),
    .Y(_09322_),
    .A1(_08787_),
    .A2(_09314_));
 sg13g2_nand2_1 _15062_ (.Y(_09323_),
    .A(_08820_),
    .B(_09316_));
 sg13g2_o21ai_1 _15063_ (.B1(net4692),
    .Y(_09324_),
    .A1(_08789_),
    .A2(_09278_));
 sg13g2_nand3_1 _15064_ (.B(_09323_),
    .C(_09324_),
    .A(net4028),
    .Y(_09325_));
 sg13g2_a22oi_1 _15065_ (.Y(_09326_),
    .B1(_09325_),
    .B2(net5099),
    .A2(_09322_),
    .A1(net4028));
 sg13g2_o21ai_1 _15066_ (.B1(_09313_),
    .Y(_00924_),
    .A1(net3720),
    .A2(_09326_));
 sg13g2_nand2_1 _15067_ (.Y(_09327_),
    .A(net4692),
    .B(net4683));
 sg13g2_nand3_1 _15068_ (.B(_09324_),
    .C(_09327_),
    .A(net4029),
    .Y(_09328_));
 sg13g2_nand2_1 _15069_ (.Y(_09329_),
    .A(net5097),
    .B(_09328_));
 sg13g2_nor2_2 _15070_ (.A(net5086),
    .B(_09274_),
    .Y(_09330_));
 sg13g2_a221oi_1 _15071_ (.B2(net5104),
    .C1(net4137),
    .B1(_09330_),
    .A1(net5108),
    .Y(_09331_),
    .A2(_08789_));
 sg13g2_nand2_1 _15072_ (.Y(_09332_),
    .A(net5097),
    .B(net4600));
 sg13g2_a22oi_1 _15073_ (.Y(_09333_),
    .B1(net4682),
    .B2(net5109),
    .A2(_08798_),
    .A1(net5097));
 sg13g2_nand3_1 _15074_ (.B(_09332_),
    .C(_09333_),
    .A(_08813_),
    .Y(_09334_));
 sg13g2_a21o_1 _15075_ (.A2(net4694),
    .A1(net5097),
    .B1(_09306_),
    .X(_09335_));
 sg13g2_o21ai_1 _15076_ (.B1(_09335_),
    .Y(_09336_),
    .A1(_09317_),
    .A2(_09334_));
 sg13g2_o21ai_1 _15077_ (.B1(_09336_),
    .Y(_09337_),
    .A1(_08787_),
    .A2(_09331_));
 sg13g2_o21ai_1 _15078_ (.B1(net4031),
    .Y(_09338_),
    .A1(_09315_),
    .A2(_09337_));
 sg13g2_a21oi_1 _15079_ (.A1(_09329_),
    .A2(_09338_),
    .Y(_09339_),
    .B1(_09250_));
 sg13g2_a21o_1 _15080_ (.A2(net1457),
    .A1(net4932),
    .B1(_09339_),
    .X(_00925_));
 sg13g2_nand2_1 _15081_ (.Y(_09340_),
    .A(net4932),
    .B(net667));
 sg13g2_a21oi_1 _15082_ (.A1(_05649_),
    .A2(_09330_),
    .Y(_09341_),
    .B1(net4696));
 sg13g2_a21oi_1 _15083_ (.A1(net5085),
    .A2(net5096),
    .Y(_09342_),
    .B1(_08807_));
 sg13g2_o21ai_1 _15084_ (.B1(net4694),
    .Y(_09343_),
    .A1(net5095),
    .A2(net4594));
 sg13g2_a21oi_1 _15085_ (.A1(_08806_),
    .A2(_09342_),
    .Y(_09344_),
    .B1(_09343_));
 sg13g2_or3_1 _15086_ (.A(_09315_),
    .B(_09341_),
    .C(_09344_),
    .X(_09345_));
 sg13g2_a22oi_1 _15087_ (.Y(_09346_),
    .B1(_09345_),
    .B2(net4028),
    .A2(_09328_),
    .A1(net5095));
 sg13g2_o21ai_1 _15088_ (.B1(_09340_),
    .Y(_00926_),
    .A1(net3720),
    .A2(_09346_));
 sg13g2_nand2_1 _15089_ (.Y(_09347_),
    .A(net4932),
    .B(net706));
 sg13g2_a22oi_1 _15090_ (.Y(_09348_),
    .B1(net4598),
    .B2(net5093),
    .A2(net4602),
    .A1(_08800_));
 sg13g2_a21o_1 _15091_ (.A2(_08798_),
    .A1(_08791_),
    .B1(net5087),
    .X(_09349_));
 sg13g2_o21ai_1 _15092_ (.B1(net4692),
    .Y(_09350_),
    .A1(_08825_),
    .A2(_09349_));
 sg13g2_o21ai_1 _15093_ (.B1(_09350_),
    .Y(_09351_),
    .A1(_09307_),
    .A2(_09348_));
 sg13g2_nor2_1 _15094_ (.A(net5090),
    .B(_08810_),
    .Y(_09352_));
 sg13g2_nor2_1 _15095_ (.A(_08809_),
    .B(_09352_),
    .Y(_09353_));
 sg13g2_nand2_1 _15096_ (.Y(_09354_),
    .A(net5092),
    .B(_05649_));
 sg13g2_nand2_1 _15097_ (.Y(_09355_),
    .A(net5096),
    .B(net4599));
 sg13g2_a22oi_1 _15098_ (.Y(_09356_),
    .B1(_09353_),
    .B2(_09354_),
    .A2(net5084),
    .A1(net5087));
 sg13g2_a21oi_1 _15099_ (.A1(net4594),
    .A2(_09356_),
    .Y(_09357_),
    .B1(_08815_));
 sg13g2_nor2_1 _15100_ (.A(_09330_),
    .B(_09357_),
    .Y(_09358_));
 sg13g2_nand3_1 _15101_ (.B(_09324_),
    .C(_09358_),
    .A(net4028),
    .Y(_09359_));
 sg13g2_a22oi_1 _15102_ (.Y(_09360_),
    .B1(_09359_),
    .B2(net5093),
    .A2(_09351_),
    .A1(net4029));
 sg13g2_o21ai_1 _15103_ (.B1(_09347_),
    .Y(_00927_),
    .A1(net3720),
    .A2(_09360_));
 sg13g2_nor2_1 _15104_ (.A(net5111),
    .B(net4602),
    .Y(_09361_));
 sg13g2_a21o_1 _15105_ (.A2(net4684),
    .A1(net5090),
    .B1(_09353_),
    .X(_09362_));
 sg13g2_and2_1 _15106_ (.A(net5106),
    .B(net5105),
    .X(_09363_));
 sg13g2_a221oi_1 _15107_ (.B2(net4600),
    .C1(_09362_),
    .B1(_09363_),
    .A1(net5087),
    .Y(_09364_),
    .A2(net4683));
 sg13g2_o21ai_1 _15108_ (.B1(_09364_),
    .Y(_09365_),
    .A1(_09257_),
    .A2(_09361_));
 sg13g2_a221oi_1 _15109_ (.B2(net4695),
    .C1(net4035),
    .B1(_09365_),
    .A1(_08818_),
    .Y(_09366_),
    .A2(_09276_));
 sg13g2_a21oi_1 _15110_ (.A1(_05650_),
    .A2(net4035),
    .Y(_09367_),
    .B1(_09366_));
 sg13g2_a22oi_1 _15111_ (.Y(_09368_),
    .B1(net3723),
    .B2(_09367_),
    .A2(net1986),
    .A1(net4931));
 sg13g2_inv_1 _15112_ (.Y(_00928_),
    .A(_09368_));
 sg13g2_nand2_1 _15113_ (.Y(_09369_),
    .A(net4930),
    .B(net2276));
 sg13g2_nor2b_1 _15114_ (.A(_08825_),
    .B_N(_08807_),
    .Y(_09370_));
 sg13g2_nand2_2 _15115_ (.Y(_09371_),
    .A(_08796_),
    .B(net4681));
 sg13g2_nor2_1 _15116_ (.A(\soc_inst.core_instr_data[3] ),
    .B(net4602),
    .Y(_09372_));
 sg13g2_nor3_1 _15117_ (.A(net5104),
    .B(_05649_),
    .C(net5090),
    .Y(_09373_));
 sg13g2_a22oi_1 _15118_ (.Y(_09374_),
    .B1(net4685),
    .B2(net5090),
    .A2(net4599),
    .A1(net5092));
 sg13g2_or2_1 _15119_ (.X(_09375_),
    .B(_09374_),
    .A(_09373_));
 sg13g2_o21ai_1 _15120_ (.B1(_09375_),
    .Y(_09376_),
    .A1(_09257_),
    .A2(_09372_));
 sg13g2_a22oi_1 _15121_ (.Y(_09377_),
    .B1(_09376_),
    .B2(net4694),
    .A2(_09371_),
    .A1(_08786_));
 sg13g2_o21ai_1 _15122_ (.B1(_09377_),
    .Y(_09378_),
    .A1(_08817_),
    .A2(_09370_));
 sg13g2_o21ai_1 _15123_ (.B1(_09378_),
    .Y(_09379_),
    .A1(net5086),
    .A2(net4029));
 sg13g2_o21ai_1 _15124_ (.B1(_09369_),
    .Y(_00929_),
    .A1(net3720),
    .A2(_09379_));
 sg13g2_nand2_1 _15125_ (.Y(_09380_),
    .A(net4930),
    .B(net2222));
 sg13g2_nor2_1 _15126_ (.A(net5108),
    .B(net4602),
    .Y(_09381_));
 sg13g2_a21oi_1 _15127_ (.A1(_08794_),
    .A2(net4600),
    .Y(_09382_),
    .B1(_09362_));
 sg13g2_o21ai_1 _15128_ (.B1(_09382_),
    .Y(_09383_),
    .A1(_09257_),
    .A2(_09381_));
 sg13g2_a21o_1 _15129_ (.A2(_09383_),
    .A1(net4695),
    .B1(net4032),
    .X(_09384_));
 sg13g2_o21ai_1 _15130_ (.B1(_09384_),
    .Y(_09385_),
    .A1(net5084),
    .A2(net4029));
 sg13g2_o21ai_1 _15131_ (.B1(_09380_),
    .Y(_00930_),
    .A1(net3720),
    .A2(_09385_));
 sg13g2_nor2_2 _15132_ (.A(net5091),
    .B(_08803_),
    .Y(_09386_));
 sg13g2_a21o_1 _15133_ (.A2(_09303_),
    .A1(_08826_),
    .B1(_09386_),
    .X(_09387_));
 sg13g2_a21oi_1 _15134_ (.A1(_09300_),
    .A2(_09387_),
    .Y(_09388_),
    .B1(net4691));
 sg13g2_nor2_1 _15135_ (.A(net5106),
    .B(net4601),
    .Y(_09389_));
 sg13g2_nor2_1 _15136_ (.A(_09257_),
    .B(_09389_),
    .Y(_09390_));
 sg13g2_a21oi_1 _15137_ (.A1(net5089),
    .A2(net4684),
    .Y(_09391_),
    .B1(net4681));
 sg13g2_nand2_1 _15138_ (.Y(_09392_),
    .A(net5103),
    .B(net4682));
 sg13g2_nand4_1 _15139_ (.B(_09303_),
    .C(_09391_),
    .A(_08813_),
    .Y(_09393_),
    .D(_09392_));
 sg13g2_o21ai_1 _15140_ (.B1(_09308_),
    .Y(_09394_),
    .A1(_09390_),
    .A2(_09393_));
 sg13g2_a21oi_1 _15141_ (.A1(net5102),
    .A2(_08788_),
    .Y(_09395_),
    .B1(net4136));
 sg13g2_o21ai_1 _15142_ (.B1(_09394_),
    .Y(_09396_),
    .A1(net4696),
    .A2(_09395_));
 sg13g2_o21ai_1 _15143_ (.B1(net4026),
    .Y(_09397_),
    .A1(_09388_),
    .A2(_09396_));
 sg13g2_o21ai_1 _15144_ (.B1(_09397_),
    .Y(_09398_),
    .A1(_05648_),
    .A2(net4025));
 sg13g2_a22oi_1 _15145_ (.Y(_09399_),
    .B1(net3723),
    .B2(_09398_),
    .A2(net1126),
    .A1(net4927));
 sg13g2_inv_1 _15146_ (.Y(_00931_),
    .A(_09399_));
 sg13g2_nand2_1 _15147_ (.Y(_09400_),
    .A(net4893),
    .B(net2366));
 sg13g2_o21ai_1 _15148_ (.B1(net4594),
    .Y(_09401_),
    .A1(_08809_),
    .A2(_09386_));
 sg13g2_nand2_1 _15149_ (.Y(_09402_),
    .A(net5101),
    .B(_09401_));
 sg13g2_a21o_1 _15150_ (.A2(_09402_),
    .A1(_09370_),
    .B1(_08819_),
    .X(_09403_));
 sg13g2_a21oi_1 _15151_ (.A1(net5099),
    .A2(_08786_),
    .Y(_09404_),
    .B1(_09272_));
 sg13g2_nor2_1 _15152_ (.A(net5105),
    .B(net4601),
    .Y(_09405_));
 sg13g2_nand2_1 _15153_ (.Y(_09406_),
    .A(net5100),
    .B(net4682));
 sg13g2_a21oi_1 _15154_ (.A1(net4595),
    .A2(_09405_),
    .Y(_09407_),
    .B1(_08801_));
 sg13g2_nand3_1 _15155_ (.B(_09391_),
    .C(_09406_),
    .A(_09318_),
    .Y(_09408_));
 sg13g2_o21ai_1 _15156_ (.B1(_09316_),
    .Y(_09409_),
    .A1(_09407_),
    .A2(_09408_));
 sg13g2_nand4_1 _15157_ (.B(_09403_),
    .C(_09404_),
    .A(net4025),
    .Y(_09410_),
    .D(_09409_));
 sg13g2_o21ai_1 _15158_ (.B1(_09410_),
    .Y(_09411_),
    .A1(net198),
    .A2(net4024));
 sg13g2_o21ai_1 _15159_ (.B1(_09400_),
    .Y(_00932_),
    .A1(net3721),
    .A2(_09411_));
 sg13g2_nand2_1 _15160_ (.Y(_09412_),
    .A(net4929),
    .B(net1239));
 sg13g2_a21o_2 _15161_ (.A2(_09386_),
    .A1(net4595),
    .B1(_08801_),
    .X(_09413_));
 sg13g2_nor2_2 _15162_ (.A(_09256_),
    .B(_09413_),
    .Y(_09414_));
 sg13g2_inv_1 _15163_ (.Y(_09415_),
    .A(_09414_));
 sg13g2_nor2_1 _15164_ (.A(_08812_),
    .B(_09414_),
    .Y(_09416_));
 sg13g2_and2_1 _15165_ (.A(_09391_),
    .B(_09416_),
    .X(_09417_));
 sg13g2_nand3_1 _15166_ (.B(net5097),
    .C(_09254_),
    .A(net5082),
    .Y(_09418_));
 sg13g2_nand2_1 _15167_ (.Y(_09419_),
    .A(_09417_),
    .B(_09418_));
 sg13g2_a21oi_1 _15168_ (.A1(_08826_),
    .A2(_09332_),
    .Y(_09420_),
    .B1(_09386_));
 sg13g2_a21oi_1 _15169_ (.A1(net5098),
    .A2(net4681),
    .Y(_09421_),
    .B1(_09420_));
 sg13g2_nand2_1 _15170_ (.Y(_09422_),
    .A(_08822_),
    .B(_09421_));
 sg13g2_a21oi_1 _15171_ (.A1(net5097),
    .A2(_08788_),
    .Y(_09423_),
    .B1(net4136));
 sg13g2_o21ai_1 _15172_ (.B1(net4025),
    .Y(_09424_),
    .A1(net4696),
    .A2(_09423_));
 sg13g2_a221oi_1 _15173_ (.B2(net4693),
    .C1(_09424_),
    .B1(_09422_),
    .A1(_09335_),
    .Y(_09425_),
    .A2(_09419_));
 sg13g2_o21ai_1 _15174_ (.B1(net3722),
    .Y(_09426_),
    .A1(net391),
    .A2(net4024));
 sg13g2_o21ai_1 _15175_ (.B1(_09412_),
    .Y(_00933_),
    .A1(_09425_),
    .A2(_09426_));
 sg13g2_nand2_1 _15176_ (.Y(_09427_),
    .A(net362),
    .B(net4032));
 sg13g2_a21oi_1 _15177_ (.A1(_08826_),
    .A2(_09355_),
    .Y(_09428_),
    .B1(_09386_));
 sg13g2_o21ai_1 _15178_ (.B1(_08799_),
    .Y(_09429_),
    .A1(net5091),
    .A2(_09254_));
 sg13g2_a21oi_1 _15179_ (.A1(_09415_),
    .A2(_09429_),
    .Y(_09430_),
    .B1(_09343_));
 sg13g2_a21oi_1 _15180_ (.A1(net5095),
    .A2(net4681),
    .Y(_09431_),
    .B1(_09428_));
 sg13g2_nand2_1 _15181_ (.Y(_09432_),
    .A(_08822_),
    .B(_09431_));
 sg13g2_a221oi_1 _15182_ (.B2(net4693),
    .C1(_09430_),
    .B1(_09432_),
    .A1(_08786_),
    .Y(_09433_),
    .A2(_09371_));
 sg13g2_o21ai_1 _15183_ (.B1(_09427_),
    .Y(_09434_),
    .A1(net4034),
    .A2(_09433_));
 sg13g2_a22oi_1 _15184_ (.Y(_09435_),
    .B1(net3722),
    .B2(_09434_),
    .A2(net2783),
    .A1(net4932));
 sg13g2_inv_1 _15185_ (.Y(_00934_),
    .A(_09435_));
 sg13g2_nand2_1 _15186_ (.Y(_09436_),
    .A(net4927),
    .B(net1587));
 sg13g2_o21ai_1 _15187_ (.B1(net4694),
    .Y(_09437_),
    .A1(net5093),
    .A2(net4594));
 sg13g2_nand2b_1 _15188_ (.Y(_09438_),
    .B(_08824_),
    .A_N(net5094));
 sg13g2_a21oi_1 _15189_ (.A1(_09401_),
    .A2(_09438_),
    .Y(_09439_),
    .B1(_08823_));
 sg13g2_nor2_1 _15190_ (.A(net4691),
    .B(_09439_),
    .Y(_09440_));
 sg13g2_nor2_1 _15191_ (.A(net4033),
    .B(_09440_),
    .Y(_09441_));
 sg13g2_o21ai_1 _15192_ (.B1(_09441_),
    .Y(_09442_),
    .A1(_09417_),
    .A2(_09437_));
 sg13g2_o21ai_1 _15193_ (.B1(_09442_),
    .Y(_09443_),
    .A1(net395),
    .A2(net4027));
 sg13g2_o21ai_1 _15194_ (.B1(_09436_),
    .Y(_00935_),
    .A1(net3721),
    .A2(_09443_));
 sg13g2_nand2_1 _15195_ (.Y(_09444_),
    .A(net4929),
    .B(net5006));
 sg13g2_nand2_1 _15196_ (.Y(_09445_),
    .A(net5111),
    .B(net4598));
 sg13g2_o21ai_1 _15197_ (.B1(net5112),
    .Y(_09446_),
    .A1(net4599),
    .A2(net4598));
 sg13g2_nor2_2 _15198_ (.A(_08793_),
    .B(_08815_),
    .Y(_09447_));
 sg13g2_nand2_1 _15199_ (.Y(_09448_),
    .A(net5112),
    .B(_09447_));
 sg13g2_a22oi_1 _15200_ (.Y(_09449_),
    .B1(_09448_),
    .B2(_09307_),
    .A2(_09446_),
    .A1(_09417_));
 sg13g2_a22oi_1 _15201_ (.Y(_09450_),
    .B1(_09261_),
    .B2(_08793_),
    .A2(_08799_),
    .A1(net5112));
 sg13g2_a21oi_1 _15202_ (.A1(_08822_),
    .A2(_09450_),
    .Y(_09451_),
    .B1(net4691));
 sg13g2_a21oi_1 _15203_ (.A1(net5111),
    .A2(_09330_),
    .Y(_09452_),
    .B1(net4136));
 sg13g2_nor2_1 _15204_ (.A(net4696),
    .B(_09452_),
    .Y(_09453_));
 sg13g2_nor4_1 _15205_ (.A(net4032),
    .B(_09449_),
    .C(_09451_),
    .D(_09453_),
    .Y(_09454_));
 sg13g2_o21ai_1 _15206_ (.B1(net3722),
    .Y(_09455_),
    .A1(net370),
    .A2(net4024));
 sg13g2_o21ai_1 _15207_ (.B1(_09444_),
    .Y(_00936_),
    .A1(_09454_),
    .A2(_09455_));
 sg13g2_nand2_1 _15208_ (.Y(_09456_),
    .A(net4893),
    .B(net5004));
 sg13g2_a21o_1 _15209_ (.A2(_09330_),
    .A1(net5110),
    .B1(net4136),
    .X(_09457_));
 sg13g2_and2_1 _15210_ (.A(\soc_inst.core_instr_data[3] ),
    .B(_08799_),
    .X(_09458_));
 sg13g2_a221oi_1 _15211_ (.B2(net4693),
    .C1(_09315_),
    .B1(_09458_),
    .A1(_08786_),
    .Y(_09459_),
    .A2(_09457_));
 sg13g2_o21ai_1 _15212_ (.B1(_09306_),
    .Y(_09460_),
    .A1(_08812_),
    .A2(_09414_));
 sg13g2_o21ai_1 _15213_ (.B1(net5084),
    .Y(_09461_),
    .A1(net5086),
    .A2(net5082));
 sg13g2_nor3_1 _15214_ (.A(_08812_),
    .B(_09414_),
    .C(_09461_),
    .Y(_09462_));
 sg13g2_o21ai_1 _15215_ (.B1(net5110),
    .Y(_09463_),
    .A1(_09306_),
    .A2(_09447_));
 sg13g2_or2_1 _15216_ (.X(_09464_),
    .B(_09463_),
    .A(_09462_));
 sg13g2_nand4_1 _15217_ (.B(_09459_),
    .C(_09460_),
    .A(net4025),
    .Y(_09465_),
    .D(_09464_));
 sg13g2_o21ai_1 _15218_ (.B1(_09465_),
    .Y(_09466_),
    .A1(net309),
    .A2(net4024));
 sg13g2_o21ai_1 _15219_ (.B1(_09456_),
    .Y(_00937_),
    .A1(net3721),
    .A2(_09466_));
 sg13g2_a21oi_1 _15220_ (.A1(net5108),
    .A2(_09461_),
    .Y(_09467_),
    .B1(net4681));
 sg13g2_nand2_1 _15221_ (.Y(_09468_),
    .A(net5108),
    .B(_09447_));
 sg13g2_a22oi_1 _15222_ (.Y(_09469_),
    .B1(_09468_),
    .B2(_09307_),
    .A2(_09467_),
    .A1(_09416_));
 sg13g2_a221oi_1 _15223_ (.B2(net5108),
    .C1(net4136),
    .B1(_09330_),
    .A1(net5104),
    .Y(_09470_),
    .A2(_08789_));
 sg13g2_a21oi_1 _15224_ (.A1(net5108),
    .A2(net4693),
    .Y(_09471_),
    .B1(_09315_));
 sg13g2_o21ai_1 _15225_ (.B1(_09471_),
    .Y(_09472_),
    .A1(net4696),
    .A2(_09470_));
 sg13g2_o21ai_1 _15226_ (.B1(net4027),
    .Y(_09473_),
    .A1(_09469_),
    .A2(_09472_));
 sg13g2_o21ai_1 _15227_ (.B1(_09473_),
    .Y(_09474_),
    .A1(_05733_),
    .A2(net4024));
 sg13g2_a22oi_1 _15228_ (.Y(_09475_),
    .B1(net3723),
    .B2(_09474_),
    .A2(net5002),
    .A1(net4928));
 sg13g2_inv_1 _15229_ (.Y(_00938_),
    .A(_09475_));
 sg13g2_and2_1 _15230_ (.A(net5106),
    .B(_09461_),
    .X(_09476_));
 sg13g2_nor4_1 _15231_ (.A(_08811_),
    .B(net4681),
    .C(_09414_),
    .D(_09476_),
    .Y(_09477_));
 sg13g2_a21oi_1 _15232_ (.A1(net5106),
    .A2(_09447_),
    .Y(_09478_),
    .B1(_09306_));
 sg13g2_nor2_1 _15233_ (.A(net5106),
    .B(_09371_),
    .Y(_09479_));
 sg13g2_a21oi_1 _15234_ (.A1(_05649_),
    .A2(net4598),
    .Y(_09480_),
    .B1(_09479_));
 sg13g2_a221oi_1 _15235_ (.B2(_08786_),
    .C1(_09315_),
    .B1(_09480_),
    .A1(net5106),
    .Y(_09481_),
    .A2(net4693));
 sg13g2_o21ai_1 _15236_ (.B1(_09481_),
    .Y(_09482_),
    .A1(_09477_),
    .A2(_09478_));
 sg13g2_mux2_1 _15237_ (.A0(net191),
    .A1(_09482_),
    .S(net4027),
    .X(_09483_));
 sg13g2_a22oi_1 _15238_ (.Y(_09484_),
    .B1(net3723),
    .B2(_09483_),
    .A2(net5000),
    .A1(net4931));
 sg13g2_inv_1 _15239_ (.Y(_00939_),
    .A(_09484_));
 sg13g2_nand2_1 _15240_ (.Y(_09485_),
    .A(net266),
    .B(net4032));
 sg13g2_or4_1 _15241_ (.A(net5088),
    .B(net5104),
    .C(_08821_),
    .D(_08825_),
    .X(_09486_));
 sg13g2_nor3_1 _15242_ (.A(net5105),
    .B(net4601),
    .C(net4595),
    .Y(_09487_));
 sg13g2_nor2_1 _15243_ (.A(_09413_),
    .B(_09487_),
    .Y(_09488_));
 sg13g2_a221oi_1 _15244_ (.B2(net5092),
    .C1(net4681),
    .B1(net4684),
    .A1(net5104),
    .Y(_09489_),
    .A2(_08789_));
 sg13g2_nand2b_1 _15245_ (.Y(_09490_),
    .B(_08810_),
    .A_N(net5105));
 sg13g2_a21oi_1 _15246_ (.A1(_09353_),
    .A2(_09490_),
    .Y(_09491_),
    .B1(_09488_));
 sg13g2_nand2_1 _15247_ (.Y(_09492_),
    .A(net5104),
    .B(_09447_));
 sg13g2_a22oi_1 _15248_ (.Y(_09493_),
    .B1(_09492_),
    .B2(_09307_),
    .A2(_09491_),
    .A1(_09489_));
 sg13g2_a21o_1 _15249_ (.A2(_08789_),
    .A1(net5092),
    .B1(net4136),
    .X(_09494_));
 sg13g2_a221oi_1 _15250_ (.B2(_08786_),
    .C1(_09493_),
    .B1(_09494_),
    .A1(net4693),
    .Y(_09495_),
    .A2(_09486_));
 sg13g2_o21ai_1 _15251_ (.B1(_09485_),
    .Y(_09496_),
    .A1(net4032),
    .A2(_09495_));
 sg13g2_a22oi_1 _15252_ (.Y(_09497_),
    .B1(net3722),
    .B2(_09496_),
    .A2(net2717),
    .A1(net4929));
 sg13g2_inv_1 _15253_ (.Y(_00940_),
    .A(_09497_));
 sg13g2_nand2_1 _15254_ (.Y(_09498_),
    .A(net4927),
    .B(net2251));
 sg13g2_o21ai_1 _15255_ (.B1(_08786_),
    .Y(_09499_),
    .A1(net5089),
    .A2(net4136));
 sg13g2_a21oi_2 _15256_ (.B1(_09306_),
    .Y(_09500_),
    .A2(_09447_),
    .A1(net5089));
 sg13g2_inv_1 _15257_ (.Y(_09501_),
    .A(_09500_));
 sg13g2_nor3_1 _15258_ (.A(net5111),
    .B(net4601),
    .C(net4595),
    .Y(_09502_));
 sg13g2_a21oi_1 _15259_ (.A1(net5093),
    .A2(net4600),
    .Y(_09503_),
    .B1(net4598));
 sg13g2_o21ai_1 _15260_ (.B1(_09277_),
    .Y(_09504_),
    .A1(_05650_),
    .A2(_09503_));
 sg13g2_o21ai_1 _15261_ (.B1(net5111),
    .Y(_09505_),
    .A1(net4685),
    .A2(net4682));
 sg13g2_o21ai_1 _15262_ (.B1(_09505_),
    .Y(_09506_),
    .A1(_09413_),
    .A2(_09502_));
 sg13g2_o21ai_1 _15263_ (.B1(_09501_),
    .Y(_09507_),
    .A1(_09504_),
    .A2(_09506_));
 sg13g2_o21ai_1 _15264_ (.B1(net5089),
    .Y(_09508_),
    .A1(_08788_),
    .A2(net4683));
 sg13g2_nand2b_1 _15265_ (.Y(_09509_),
    .B(net4693),
    .A_N(_09508_));
 sg13g2_nand4_1 _15266_ (.B(_09499_),
    .C(_09507_),
    .A(net4025),
    .Y(_09510_),
    .D(_09509_));
 sg13g2_o21ai_1 _15267_ (.B1(_09510_),
    .Y(_09511_),
    .A1(net2096),
    .A2(net4025));
 sg13g2_o21ai_1 _15268_ (.B1(_09498_),
    .Y(_00941_),
    .A1(net3720),
    .A2(_09511_));
 sg13g2_nand2_1 _15269_ (.Y(_09512_),
    .A(net4929),
    .B(net1597));
 sg13g2_a221oi_1 _15270_ (.B2(net5102),
    .C1(net4136),
    .B1(net4681),
    .A1(net5106),
    .Y(_09513_),
    .A2(_08788_));
 sg13g2_nand2b_1 _15271_ (.Y(_09514_),
    .B(_08786_),
    .A_N(_09513_));
 sg13g2_nor3_1 _15272_ (.A(net5107),
    .B(net4601),
    .C(net4595),
    .Y(_09515_));
 sg13g2_a221oi_1 _15273_ (.B2(net5107),
    .C1(_09504_),
    .B1(net4682),
    .A1(net5102),
    .Y(_09516_),
    .A2(net4685));
 sg13g2_o21ai_1 _15274_ (.B1(_09516_),
    .Y(_09517_),
    .A1(_09413_),
    .A2(_09515_));
 sg13g2_a21oi_1 _15275_ (.A1(_09392_),
    .A2(_09445_),
    .Y(_09518_),
    .B1(net4691));
 sg13g2_a21oi_1 _15276_ (.A1(_09501_),
    .A2(_09517_),
    .Y(_09519_),
    .B1(_09518_));
 sg13g2_nand3_1 _15277_ (.B(_09514_),
    .C(_09519_),
    .A(net4025),
    .Y(_09520_));
 sg13g2_o21ai_1 _15278_ (.B1(_09520_),
    .Y(_09521_),
    .A1(net275),
    .A2(net4024));
 sg13g2_o21ai_1 _15279_ (.B1(_09512_),
    .Y(_00942_),
    .A1(net3721),
    .A2(_09521_));
 sg13g2_nor3_1 _15280_ (.A(net5110),
    .B(net4601),
    .C(net4595),
    .Y(_09522_));
 sg13g2_o21ai_1 _15281_ (.B1(net5104),
    .Y(_09523_),
    .A1(net4685),
    .A2(net4682));
 sg13g2_o21ai_1 _15282_ (.B1(_09523_),
    .Y(_09524_),
    .A1(_09413_),
    .A2(_09522_));
 sg13g2_o21ai_1 _15283_ (.B1(_09501_),
    .Y(_09525_),
    .A1(_09504_),
    .A2(_09524_));
 sg13g2_a22oi_1 _15284_ (.Y(_09526_),
    .B1(net4683),
    .B2(net5099),
    .A2(net4598),
    .A1(net5110));
 sg13g2_a21o_1 _15285_ (.A2(_09526_),
    .A1(_08827_),
    .B1(net4691),
    .X(_09527_));
 sg13g2_o21ai_1 _15286_ (.B1(_09272_),
    .Y(_09528_),
    .A1(net5099),
    .A2(_09371_));
 sg13g2_nand3_1 _15287_ (.B(_09527_),
    .C(_09528_),
    .A(_09525_),
    .Y(_09529_));
 sg13g2_mux2_1 _15288_ (.A0(net1441),
    .A1(_09529_),
    .S(net4031),
    .X(_09530_));
 sg13g2_a22oi_1 _15289_ (.Y(_09531_),
    .B1(net3723),
    .B2(_09530_),
    .A2(net2749),
    .A1(net4930));
 sg13g2_inv_1 _15290_ (.Y(_00943_),
    .A(_09531_));
 sg13g2_nand2_1 _15291_ (.Y(_09532_),
    .A(net4929),
    .B(net2077));
 sg13g2_a21oi_1 _15292_ (.A1(net5089),
    .A2(net4683),
    .Y(_09533_),
    .B1(_09504_));
 sg13g2_nor3_1 _15293_ (.A(net5109),
    .B(net4601),
    .C(net4595),
    .Y(_09534_));
 sg13g2_nor2_1 _15294_ (.A(_09413_),
    .B(_09534_),
    .Y(_09535_));
 sg13g2_a21oi_1 _15295_ (.A1(net5097),
    .A2(net4684),
    .Y(_09536_),
    .B1(_09535_));
 sg13g2_a21o_1 _15296_ (.A2(_09536_),
    .A1(_09533_),
    .B1(_09500_),
    .X(_09537_));
 sg13g2_o21ai_1 _15297_ (.B1(_09272_),
    .Y(_09538_),
    .A1(net5097),
    .A2(_09371_));
 sg13g2_a21oi_1 _15298_ (.A1(_09537_),
    .A2(_09538_),
    .Y(_09539_),
    .B1(net4032));
 sg13g2_a21oi_1 _15299_ (.A1(net452),
    .A2(net4034),
    .Y(_09540_),
    .B1(_09539_));
 sg13g2_o21ai_1 _15300_ (.B1(_09532_),
    .Y(_00944_),
    .A1(net3721),
    .A2(_09540_));
 sg13g2_nand2_1 _15301_ (.Y(_09541_),
    .A(net4943),
    .B(net2325));
 sg13g2_o21ai_1 _15302_ (.B1(_09533_),
    .Y(_09542_),
    .A1(_08801_),
    .A2(_09386_));
 sg13g2_a21oi_1 _15303_ (.A1(net5095),
    .A2(net4684),
    .Y(_09543_),
    .B1(_09542_));
 sg13g2_o21ai_1 _15304_ (.B1(_09272_),
    .Y(_09544_),
    .A1(net5095),
    .A2(_09371_));
 sg13g2_o21ai_1 _15305_ (.B1(_09544_),
    .Y(_09545_),
    .A1(_09500_),
    .A2(_09543_));
 sg13g2_nor2_1 _15306_ (.A(net4033),
    .B(_09545_),
    .Y(_09546_));
 sg13g2_o21ai_1 _15307_ (.B1(net3729),
    .Y(_09547_),
    .A1(net1136),
    .A2(net4030));
 sg13g2_o21ai_1 _15308_ (.B1(_09541_),
    .Y(_00945_),
    .A1(_09546_),
    .A2(_09547_));
 sg13g2_nand2_1 _15309_ (.Y(_09548_),
    .A(net4929),
    .B(net2122));
 sg13g2_a21oi_1 _15310_ (.A1(net5093),
    .A2(_08794_),
    .Y(_09549_),
    .B1(_09355_));
 sg13g2_a21oi_1 _15311_ (.A1(net5100),
    .A2(net4684),
    .Y(_09550_),
    .B1(_09549_));
 sg13g2_nor2b_1 _15312_ (.A(_09542_),
    .B_N(_09550_),
    .Y(_09551_));
 sg13g2_o21ai_1 _15313_ (.B1(net4026),
    .Y(_09552_),
    .A1(_09500_),
    .A2(_09551_));
 sg13g2_o21ai_1 _15314_ (.B1(_09552_),
    .Y(_09553_),
    .A1(net321),
    .A2(net4024));
 sg13g2_o21ai_1 _15315_ (.B1(_09548_),
    .Y(_00946_),
    .A1(net3721),
    .A2(_09553_));
 sg13g2_nand2_1 _15316_ (.Y(_09554_),
    .A(net4892),
    .B(net2720));
 sg13g2_a21oi_1 _15317_ (.A1(net5089),
    .A2(net4684),
    .Y(_09555_),
    .B1(_09542_));
 sg13g2_o21ai_1 _15318_ (.B1(net4026),
    .Y(_09556_),
    .A1(_09500_),
    .A2(_09555_));
 sg13g2_o21ai_1 _15319_ (.B1(_09556_),
    .Y(_09557_),
    .A1(net319),
    .A2(net4024));
 sg13g2_o21ai_1 _15320_ (.B1(_09554_),
    .Y(_00947_),
    .A1(net3721),
    .A2(_09557_));
 sg13g2_a22oi_1 _15321_ (.Y(_00948_),
    .B1(net3727),
    .B2(_05435_),
    .A2(_05520_),
    .A1(net4985));
 sg13g2_a22oi_1 _15322_ (.Y(_00949_),
    .B1(net3726),
    .B2(_05436_),
    .A2(_05519_),
    .A1(net4985));
 sg13g2_a22oi_1 _15323_ (.Y(_00950_),
    .B1(net3726),
    .B2(_05437_),
    .A2(_05522_),
    .A1(net4985));
 sg13g2_a22oi_1 _15324_ (.Y(_00951_),
    .B1(net3726),
    .B2(_05438_),
    .A2(_05521_),
    .A1(net4982));
 sg13g2_a22oi_1 _15325_ (.Y(_00952_),
    .B1(net3726),
    .B2(_05440_),
    .A2(_05523_),
    .A1(net4973));
 sg13g2_a22oi_1 _15326_ (.Y(_00953_),
    .B1(net3726),
    .B2(_05442_),
    .A2(_05524_),
    .A1(net4982));
 sg13g2_a22oi_1 _15327_ (.Y(_00954_),
    .B1(net3727),
    .B2(_05444_),
    .A2(_05525_),
    .A1(net4973));
 sg13g2_a22oi_1 _15328_ (.Y(_00955_),
    .B1(net3727),
    .B2(_05445_),
    .A2(_05526_),
    .A1(net4982));
 sg13g2_a22oi_1 _15329_ (.Y(_00956_),
    .B1(net3726),
    .B2(_05446_),
    .A2(_05527_),
    .A1(net4965));
 sg13g2_a22oi_1 _15330_ (.Y(_00957_),
    .B1(net3726),
    .B2(_05448_),
    .A2(_05528_),
    .A1(net4965));
 sg13g2_a22oi_1 _15331_ (.Y(_00958_),
    .B1(net3726),
    .B2(_05450_),
    .A2(_05529_),
    .A1(net4961));
 sg13g2_a22oi_1 _15332_ (.Y(_00959_),
    .B1(net3725),
    .B2(_05452_),
    .A2(_05530_),
    .A1(net4961));
 sg13g2_a22oi_1 _15333_ (.Y(_00960_),
    .B1(net3725),
    .B2(_05453_),
    .A2(_05531_),
    .A1(net4961));
 sg13g2_a22oi_1 _15334_ (.Y(_00961_),
    .B1(net3728),
    .B2(_05454_),
    .A2(_05532_),
    .A1(net4964));
 sg13g2_a22oi_1 _15335_ (.Y(_00962_),
    .B1(net3725),
    .B2(_05455_),
    .A2(_05533_),
    .A1(net4961));
 sg13g2_a22oi_1 _15336_ (.Y(_00963_),
    .B1(net3725),
    .B2(_05456_),
    .A2(_05534_),
    .A1(net4963));
 sg13g2_a22oi_1 _15337_ (.Y(_00964_),
    .B1(net3724),
    .B2(_05457_),
    .A2(_05535_),
    .A1(net4914));
 sg13g2_a22oi_1 _15338_ (.Y(_00965_),
    .B1(net3724),
    .B2(_05458_),
    .A2(_05536_),
    .A1(net4915));
 sg13g2_a22oi_1 _15339_ (.Y(_00966_),
    .B1(net3724),
    .B2(_05459_),
    .A2(_05537_),
    .A1(net4914));
 sg13g2_a22oi_1 _15340_ (.Y(_00967_),
    .B1(net3724),
    .B2(_05460_),
    .A2(_05538_),
    .A1(net4914));
 sg13g2_a22oi_1 _15341_ (.Y(_00968_),
    .B1(net3724),
    .B2(_05461_),
    .A2(_05539_),
    .A1(net4952));
 sg13g2_a22oi_1 _15342_ (.Y(_00969_),
    .B1(net3724),
    .B2(_05462_),
    .A2(_05540_),
    .A1(net4953));
 sg13g2_a22oi_1 _15343_ (.Y(_00970_),
    .B1(net3724),
    .B2(_05464_),
    .A2(_05541_),
    .A1(net4954));
 sg13g2_a22oi_1 _15344_ (.Y(_00971_),
    .B1(net3724),
    .B2(_05465_),
    .A2(_05542_),
    .A1(net4953));
 sg13g2_nor2_1 _15345_ (.A(net2029),
    .B(net3723),
    .Y(_09558_));
 sg13g2_a21oi_1 _15346_ (.A1(net4034),
    .A2(net3722),
    .Y(_00972_),
    .B1(_09558_));
 sg13g2_mux2_1 _15347_ (.A0(net1213),
    .A1(net1339),
    .S(net4981),
    .X(_00973_));
 sg13g2_mux2_1 _15348_ (.A0(net808),
    .A1(\soc_inst.cpu_core.mem_rs1_data[1] ),
    .S(net4907),
    .X(_00974_));
 sg13g2_mux2_1 _15349_ (.A0(net801),
    .A1(net959),
    .S(net4981),
    .X(_00975_));
 sg13g2_mux2_1 _15350_ (.A0(\soc_inst.cpu_core.ex_rs1_data[3] ),
    .A1(net774),
    .S(net4981),
    .X(_00976_));
 sg13g2_mux2_1 _15351_ (.A0(net257),
    .A1(net660),
    .S(net4941),
    .X(_00977_));
 sg13g2_mux2_1 _15352_ (.A0(net305),
    .A1(net812),
    .S(net4945),
    .X(_00978_));
 sg13g2_mux2_1 _15353_ (.A0(net352),
    .A1(net1355),
    .S(net4943),
    .X(_00979_));
 sg13g2_mux2_1 _15354_ (.A0(net271),
    .A1(net457),
    .S(net4943),
    .X(_00980_));
 sg13g2_mux2_1 _15355_ (.A0(net1144),
    .A1(net1494),
    .S(net4939),
    .X(_00981_));
 sg13g2_mux2_1 _15356_ (.A0(net2589),
    .A1(net2600),
    .S(net4984),
    .X(_00982_));
 sg13g2_mux2_1 _15357_ (.A0(net2456),
    .A1(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .S(net4994),
    .X(_00983_));
 sg13g2_mux2_1 _15358_ (.A0(net637),
    .A1(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .S(net4924),
    .X(_00984_));
 sg13g2_mux2_1 _15359_ (.A0(net2107),
    .A1(net2201),
    .S(net4922),
    .X(_00985_));
 sg13g2_mux2_1 _15360_ (.A0(net780),
    .A1(net928),
    .S(net4918),
    .X(_00986_));
 sg13g2_mux2_1 _15361_ (.A0(net835),
    .A1(net2328),
    .S(net4961),
    .X(_00987_));
 sg13g2_mux2_1 _15362_ (.A0(net444),
    .A1(net932),
    .S(net4922),
    .X(_00988_));
 sg13g2_mux2_1 _15363_ (.A0(net1137),
    .A1(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .S(net4957),
    .X(_00989_));
 sg13g2_mux2_1 _15364_ (.A0(net2223),
    .A1(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .S(net4953),
    .X(_00990_));
 sg13g2_mux2_1 _15365_ (.A0(net873),
    .A1(net2128),
    .S(net4957),
    .X(_00991_));
 sg13g2_mux2_1 _15366_ (.A0(net737),
    .A1(net2381),
    .S(net4967),
    .X(_00992_));
 sg13g2_mux2_1 _15367_ (.A0(net1314),
    .A1(net1576),
    .S(net4954),
    .X(_00993_));
 sg13g2_mux2_1 _15368_ (.A0(net730),
    .A1(net2253),
    .S(net4967),
    .X(_00994_));
 sg13g2_mux2_1 _15369_ (.A0(net647),
    .A1(net2367),
    .S(net4967),
    .X(_00995_));
 sg13g2_mux2_1 _15370_ (.A0(net755),
    .A1(net2324),
    .S(net4957),
    .X(_00996_));
 sg13g2_mux2_1 _15371_ (.A0(net1256),
    .A1(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .S(net4992),
    .X(_00997_));
 sg13g2_mux2_1 _15372_ (.A0(net877),
    .A1(net1005),
    .S(net4991),
    .X(_00998_));
 sg13g2_mux2_1 _15373_ (.A0(net2264),
    .A1(net2640),
    .S(net4988),
    .X(_00999_));
 sg13g2_mux2_1 _15374_ (.A0(net934),
    .A1(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .S(net4988),
    .X(_01000_));
 sg13g2_mux2_1 _15375_ (.A0(net916),
    .A1(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .S(net4989),
    .X(_01001_));
 sg13g2_mux2_1 _15376_ (.A0(net847),
    .A1(net1095),
    .S(net4990),
    .X(_01002_));
 sg13g2_mux2_1 _15377_ (.A0(net2092),
    .A1(net2695),
    .S(net4987),
    .X(_01003_));
 sg13g2_mux2_1 _15378_ (.A0(net2633),
    .A1(net4879),
    .S(net4988),
    .X(_01004_));
 sg13g2_a22oi_1 _15379_ (.Y(_09559_),
    .B1(net4131),
    .B2(net1676),
    .A2(net4945),
    .A1(_00267_));
 sg13g2_inv_1 _15380_ (.Y(_01005_),
    .A(net1677));
 sg13g2_a22oi_1 _15381_ (.Y(_09560_),
    .B1(net4131),
    .B2(net1426),
    .A2(net4945),
    .A1(_00268_));
 sg13g2_inv_1 _15382_ (.Y(_01006_),
    .A(net1427));
 sg13g2_a22oi_1 _15383_ (.Y(_09561_),
    .B1(net2580),
    .B2(net4131),
    .A2(\soc_inst.cpu_core.id_instr[2] ),
    .A1(net4936));
 sg13g2_inv_1 _15384_ (.Y(_01007_),
    .A(net2581));
 sg13g2_a22oi_1 _15385_ (.Y(_09562_),
    .B1(net2798),
    .B2(net4131),
    .A2(\soc_inst.cpu_core.id_instr[3] ),
    .A1(net4945));
 sg13g2_inv_1 _15386_ (.Y(_01008_),
    .A(net2799));
 sg13g2_a22oi_1 _15387_ (.Y(_09563_),
    .B1(net4131),
    .B2(net2170),
    .A2(net4944),
    .A1(_00269_));
 sg13g2_inv_1 _15388_ (.Y(_01009_),
    .A(net2171));
 sg13g2_a22oi_1 _15389_ (.Y(_09564_),
    .B1(net2608),
    .B2(net4132),
    .A2(net541),
    .A1(net4940));
 sg13g2_inv_1 _15390_ (.Y(_01010_),
    .A(_09564_));
 sg13g2_a22oi_1 _15391_ (.Y(_09565_),
    .B1(net5016),
    .B2(net4132),
    .A2(net4878),
    .A1(net4937));
 sg13g2_inv_1 _15392_ (.Y(_01011_),
    .A(net2943));
 sg13g2_a22oi_1 _15393_ (.Y(_09566_),
    .B1(net4130),
    .B2(net905),
    .A2(\soc_inst.cpu_core.id_instr[7] ),
    .A1(net4927));
 sg13g2_inv_1 _15394_ (.Y(_01012_),
    .A(net906));
 sg13g2_a22oi_1 _15395_ (.Y(_09567_),
    .B1(net4130),
    .B2(net568),
    .A2(\soc_inst.cpu_core.id_instr[8] ),
    .A1(net4931));
 sg13g2_inv_1 _15396_ (.Y(_01013_),
    .A(net569));
 sg13g2_a22oi_1 _15397_ (.Y(_09568_),
    .B1(net4130),
    .B2(net1457),
    .A2(\soc_inst.cpu_core.id_instr[9] ),
    .A1(net4930));
 sg13g2_inv_1 _15398_ (.Y(_01014_),
    .A(net1458));
 sg13g2_a22oi_1 _15399_ (.Y(_09569_),
    .B1(net4130),
    .B2(net667),
    .A2(net841),
    .A1(net4931));
 sg13g2_inv_1 _15400_ (.Y(_01015_),
    .A(_09569_));
 sg13g2_a22oi_1 _15401_ (.Y(_09570_),
    .B1(net4130),
    .B2(net706),
    .A2(net1253),
    .A1(net4930));
 sg13g2_inv_1 _15402_ (.Y(_01016_),
    .A(_09570_));
 sg13g2_a22oi_1 _15403_ (.Y(_09571_),
    .B1(net1986),
    .B2(net4131),
    .A2(\soc_inst.cpu_core.id_funct3[0] ),
    .A1(net4908));
 sg13g2_inv_1 _15404_ (.Y(_01017_),
    .A(net1987));
 sg13g2_a22oi_1 _15405_ (.Y(_09572_),
    .B1(net2276),
    .B2(net4128),
    .A2(net2498),
    .A1(net4907));
 sg13g2_inv_1 _15406_ (.Y(_01018_),
    .A(_09572_));
 sg13g2_a22oi_1 _15407_ (.Y(_09573_),
    .B1(net2222),
    .B2(net4128),
    .A2(net2386),
    .A1(net4907));
 sg13g2_inv_1 _15408_ (.Y(_01019_),
    .A(_09573_));
 sg13g2_a22oi_1 _15409_ (.Y(_09574_),
    .B1(net4132),
    .B2(net1126),
    .A2(net1048),
    .A1(net4937));
 sg13g2_inv_1 _15410_ (.Y(_01020_),
    .A(_09574_));
 sg13g2_a22oi_1 _15411_ (.Y(_09575_),
    .B1(net4127),
    .B2(net2366),
    .A2(net2151),
    .A1(net4898));
 sg13g2_inv_1 _15412_ (.Y(_01021_),
    .A(_09575_));
 sg13g2_a22oi_1 _15413_ (.Y(_09576_),
    .B1(net4127),
    .B2(net5008),
    .A2(net1003),
    .A1(net4899));
 sg13g2_inv_1 _15414_ (.Y(_01022_),
    .A(_09576_));
 sg13g2_a22oi_1 _15415_ (.Y(_09577_),
    .B1(net4128),
    .B2(\soc_inst.cpu_core.if_instr[18] ),
    .A2(net1064),
    .A1(net4901));
 sg13g2_inv_1 _15416_ (.Y(_01023_),
    .A(net1065));
 sg13g2_a22oi_1 _15417_ (.Y(_09578_),
    .B1(net4127),
    .B2(net1587),
    .A2(net1242),
    .A1(net4901));
 sg13g2_inv_1 _15418_ (.Y(_01024_),
    .A(_09578_));
 sg13g2_a22oi_1 _15419_ (.Y(_09579_),
    .B1(net5006),
    .B2(net4127),
    .A2(net2702),
    .A1(net4898));
 sg13g2_inv_1 _15420_ (.Y(_01025_),
    .A(_09579_));
 sg13g2_a22oi_1 _15421_ (.Y(_09580_),
    .B1(net5004),
    .B2(net4127),
    .A2(net2631),
    .A1(net4898));
 sg13g2_inv_1 _15422_ (.Y(_01026_),
    .A(net2632));
 sg13g2_a22oi_1 _15423_ (.Y(_09581_),
    .B1(net5002),
    .B2(net4128),
    .A2(net2330),
    .A1(net4912));
 sg13g2_inv_1 _15424_ (.Y(_01027_),
    .A(_09581_));
 sg13g2_a22oi_1 _15425_ (.Y(_09582_),
    .B1(net5000),
    .B2(net4127),
    .A2(net2585),
    .A1(net4901));
 sg13g2_inv_1 _15426_ (.Y(_01028_),
    .A(net2586));
 sg13g2_a22oi_1 _15427_ (.Y(_09583_),
    .B1(\soc_inst.cpu_core.if_imm12[4] ),
    .B2(net4128),
    .A2(net2354),
    .A1(net4905));
 sg13g2_inv_1 _15428_ (.Y(_01029_),
    .A(net2355));
 sg13g2_a22oi_1 _15429_ (.Y(_09584_),
    .B1(net2251),
    .B2(net4128),
    .A2(net720),
    .A1(net4918));
 sg13g2_inv_1 _15430_ (.Y(_01030_),
    .A(_09584_));
 sg13g2_a22oi_1 _15431_ (.Y(_09585_),
    .B1(net1597),
    .B2(net4128),
    .A2(net2139),
    .A1(net4902));
 sg13g2_inv_1 _15432_ (.Y(_01031_),
    .A(_09585_));
 sg13g2_a22oi_1 _15433_ (.Y(_09586_),
    .B1(\soc_inst.cpu_core.if_funct7[2] ),
    .B2(net4129),
    .A2(net2358),
    .A1(net4905));
 sg13g2_inv_1 _15434_ (.Y(_01032_),
    .A(net2359));
 sg13g2_a22oi_1 _15435_ (.Y(_09587_),
    .B1(net2077),
    .B2(net4127),
    .A2(net2307),
    .A1(net4904));
 sg13g2_inv_1 _15436_ (.Y(_01033_),
    .A(_09587_));
 sg13g2_a22oi_1 _15437_ (.Y(_09588_),
    .B1(net2325),
    .B2(net4129),
    .A2(net567),
    .A1(net4919));
 sg13g2_inv_1 _15438_ (.Y(_01034_),
    .A(_09588_));
 sg13g2_nand2_1 _15439_ (.Y(_09589_),
    .A(net2122),
    .B(net4125));
 sg13g2_a22oi_1 _15440_ (.Y(_09590_),
    .B1(net2122),
    .B2(net4129),
    .A2(net583),
    .A1(net4923));
 sg13g2_inv_1 _15441_ (.Y(_01035_),
    .A(_09590_));
 sg13g2_a22oi_1 _15442_ (.Y(_09591_),
    .B1(\soc_inst.cpu_core.if_funct7[6] ),
    .B2(net4129),
    .A2(net2505),
    .A1(net4924));
 sg13g2_inv_1 _15443_ (.Y(_01036_),
    .A(net2506));
 sg13g2_nor3_2 _15444_ (.A(net5009),
    .B(net5008),
    .C(net5007),
    .Y(_09592_));
 sg13g2_or3_1 _15445_ (.A(net5009),
    .B(net5008),
    .C(net5007),
    .X(_09593_));
 sg13g2_o21ai_1 _15446_ (.B1(net4133),
    .Y(_09594_),
    .A1(net5010),
    .A2(_09593_));
 sg13g2_nand2_2 _15447_ (.Y(_09595_),
    .A(net5008),
    .B(net5007));
 sg13g2_nand2b_1 _15448_ (.Y(_09596_),
    .B(net5010),
    .A_N(net5009));
 sg13g2_nor2_1 _15449_ (.A(_09595_),
    .B(_09596_),
    .Y(_09597_));
 sg13g2_nand2b_2 _15450_ (.Y(_09598_),
    .B(net5008),
    .A_N(net5007));
 sg13g2_nor3_1 _15451_ (.A(net5010),
    .B(net5009),
    .C(_09598_),
    .Y(_09599_));
 sg13g2_nor2_1 _15452_ (.A(_09596_),
    .B(_09598_),
    .Y(_09600_));
 sg13g2_nand2b_2 _15453_ (.Y(_09601_),
    .B(net5007),
    .A_N(net5008));
 sg13g2_nor2_1 _15454_ (.A(_09596_),
    .B(_09601_),
    .Y(_09602_));
 sg13g2_nand2b_2 _15455_ (.Y(_09603_),
    .B(net5009),
    .A_N(net5010));
 sg13g2_nor2_1 _15456_ (.A(_09595_),
    .B(_09603_),
    .Y(_09604_));
 sg13g2_a22oi_1 _15457_ (.Y(_09605_),
    .B1(net4571),
    .B2(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][0] ));
 sg13g2_nand2_1 _15458_ (.Y(_09606_),
    .A(net5010),
    .B(net5009));
 sg13g2_nor3_1 _15459_ (.A(net5008),
    .B(net5007),
    .C(_09606_),
    .Y(_09607_));
 sg13g2_nor2_1 _15460_ (.A(_09598_),
    .B(_09606_),
    .Y(_09608_));
 sg13g2_a22oi_1 _15461_ (.Y(_09609_),
    .B1(net4561),
    .B2(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .A2(net4566),
    .A1(\soc_inst.cpu_core.register_file.registers[3][0] ));
 sg13g2_nor3_1 _15462_ (.A(net5010),
    .B(net5009),
    .C(_09595_),
    .Y(_09610_));
 sg13g2_nor2_1 _15463_ (.A(_09598_),
    .B(_09603_),
    .Y(_09611_));
 sg13g2_nor3_1 _15464_ (.A(net5008),
    .B(net5007),
    .C(_09603_),
    .Y(_09612_));
 sg13g2_nor2_1 _15465_ (.A(_09595_),
    .B(_09606_),
    .Y(_09613_));
 sg13g2_nor2_1 _15466_ (.A(_09601_),
    .B(_09603_),
    .Y(_09614_));
 sg13g2_nor2_1 _15467_ (.A(_09601_),
    .B(_09606_),
    .Y(_09615_));
 sg13g2_nor3_1 _15468_ (.A(net5010),
    .B(net5009),
    .C(_09601_),
    .Y(_09616_));
 sg13g2_a22oi_1 _15469_ (.Y(_09617_),
    .B1(net4551),
    .B2(\soc_inst.cpu_core.register_file.registers[6][0] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][0] ));
 sg13g2_a22oi_1 _15470_ (.Y(_09618_),
    .B1(net4556),
    .B2(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .A2(net4581),
    .A1(\soc_inst.cpu_core.register_file.registers[5][0] ));
 sg13g2_nand3_1 _15471_ (.B(_09617_),
    .C(_09618_),
    .A(_09605_),
    .Y(_09619_));
 sg13g2_a221oi_1 _15472_ (.B2(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .C1(_09619_),
    .B1(net4531),
    .A1(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .Y(_09620_),
    .A2(net4541));
 sg13g2_a22oi_1 _15473_ (.Y(_09621_),
    .B1(net4546),
    .B2(\soc_inst.cpu_core.register_file.registers[2][0] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][0] ));
 sg13g2_a22oi_1 _15474_ (.Y(_09622_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][0] ),
    .A2(net4536),
    .A1(\soc_inst.cpu_core.register_file.registers[10][0] ));
 sg13g2_nand4_1 _15475_ (.B(_09620_),
    .C(_09621_),
    .A(_09609_),
    .Y(_09623_),
    .D(_09622_));
 sg13g2_a21oi_1 _15476_ (.A1(net872),
    .A2(net4678),
    .Y(_09624_),
    .B1(_09623_));
 sg13g2_nor2_2 _15477_ (.A(net4082),
    .B(_09624_),
    .Y(_09625_));
 sg13g2_a21o_1 _15478_ (.A2(net2920),
    .A1(net4889),
    .B1(_09625_),
    .X(_01037_));
 sg13g2_a22oi_1 _15479_ (.Y(_09626_),
    .B1(net4571),
    .B2(\soc_inst.cpu_core.register_file.registers[14][1] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][1] ));
 sg13g2_a22oi_1 _15480_ (.Y(_09627_),
    .B1(net4551),
    .B2(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .A2(net4582),
    .A1(\soc_inst.cpu_core.register_file.registers[5][1] ));
 sg13g2_a22oi_1 _15481_ (.Y(_09628_),
    .B1(net4556),
    .B2(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .A2(net4561),
    .A1(\soc_inst.cpu_core.register_file.registers[7][1] ));
 sg13g2_a22oi_1 _15482_ (.Y(_09629_),
    .B1(net4547),
    .B2(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .A2(net4567),
    .A1(\soc_inst.cpu_core.register_file.registers[3][1] ));
 sg13g2_nand3_1 _15483_ (.B(_09628_),
    .C(_09629_),
    .A(_09627_),
    .Y(_09630_));
 sg13g2_a221oi_1 _15484_ (.B2(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .C1(_09630_),
    .B1(net4536),
    .A1(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .Y(_09631_),
    .A2(net4541));
 sg13g2_a22oi_1 _15485_ (.Y(_09632_),
    .B1(net4531),
    .B2(\soc_inst.cpu_core.register_file.registers[11][1] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][1] ));
 sg13g2_a22oi_1 _15486_ (.Y(_09633_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][1] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][1] ));
 sg13g2_nand4_1 _15487_ (.B(_09631_),
    .C(_09632_),
    .A(_09626_),
    .Y(_09634_),
    .D(_09633_));
 sg13g2_a21oi_1 _15488_ (.A1(net986),
    .A2(net4678),
    .Y(_09635_),
    .B1(_09634_));
 sg13g2_nor2_2 _15489_ (.A(net4082),
    .B(_09635_),
    .Y(_09636_));
 sg13g2_a21o_1 _15490_ (.A2(net1250),
    .A1(net4889),
    .B1(_09636_),
    .X(_01038_));
 sg13g2_a22oi_1 _15491_ (.Y(_09637_),
    .B1(net4531),
    .B2(\soc_inst.cpu_core.register_file.registers[11][2] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][2] ));
 sg13g2_a22oi_1 _15492_ (.Y(_09638_),
    .B1(net4566),
    .B2(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .A2(net4571),
    .A1(\soc_inst.cpu_core.register_file.registers[14][2] ));
 sg13g2_a22oi_1 _15493_ (.Y(_09639_),
    .B1(net4556),
    .B2(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .A2(net4581),
    .A1(\soc_inst.cpu_core.register_file.registers[5][2] ));
 sg13g2_a22oi_1 _15494_ (.Y(_09640_),
    .B1(net4536),
    .B2(\soc_inst.cpu_core.register_file.registers[10][2] ),
    .A2(net4551),
    .A1(\soc_inst.cpu_core.register_file.registers[6][2] ));
 sg13g2_nand3_1 _15495_ (.B(_09639_),
    .C(_09640_),
    .A(_09638_),
    .Y(_09641_));
 sg13g2_a221oi_1 _15496_ (.B2(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .C1(_09641_),
    .B1(net4561),
    .A1(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .Y(_09642_),
    .A2(net4576));
 sg13g2_a22oi_1 _15497_ (.Y(_09643_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][2] ),
    .A2(net4546),
    .A1(\soc_inst.cpu_core.register_file.registers[2][2] ));
 sg13g2_a22oi_1 _15498_ (.Y(_09644_),
    .B1(net4541),
    .B2(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][2] ));
 sg13g2_nand4_1 _15499_ (.B(_09642_),
    .C(_09643_),
    .A(_09637_),
    .Y(_09645_),
    .D(_09644_));
 sg13g2_a21oi_1 _15500_ (.A1(net673),
    .A2(net4680),
    .Y(_09646_),
    .B1(_09645_));
 sg13g2_nor2_2 _15501_ (.A(net4082),
    .B(_09646_),
    .Y(_09647_));
 sg13g2_a21o_1 _15502_ (.A2(net2918),
    .A1(net4894),
    .B1(_09647_),
    .X(_01039_));
 sg13g2_a22oi_1 _15503_ (.Y(_09648_),
    .B1(net4531),
    .B2(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .A2(net4546),
    .A1(\soc_inst.cpu_core.register_file.registers[2][3] ));
 sg13g2_a22oi_1 _15504_ (.Y(_09649_),
    .B1(net4551),
    .B2(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][3] ));
 sg13g2_a22oi_1 _15505_ (.Y(_09650_),
    .B1(net4571),
    .B2(\soc_inst.cpu_core.register_file.registers[14][3] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][3] ));
 sg13g2_nand3_1 _15506_ (.B(_09649_),
    .C(_09650_),
    .A(_09648_),
    .Y(_09651_));
 sg13g2_a221oi_1 _15507_ (.B2(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .C1(_09651_),
    .B1(net4541),
    .A1(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .Y(_09652_),
    .A2(net4556));
 sg13g2_a22oi_1 _15508_ (.Y(_09653_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][3] ),
    .A2(net4566),
    .A1(\soc_inst.cpu_core.register_file.registers[3][3] ));
 sg13g2_a22oi_1 _15509_ (.Y(_09654_),
    .B1(net4561),
    .B2(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .A2(net4581),
    .A1(\soc_inst.cpu_core.register_file.registers[5][3] ));
 sg13g2_a22oi_1 _15510_ (.Y(_09655_),
    .B1(net4536),
    .B2(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][3] ));
 sg13g2_nand4_1 _15511_ (.B(_09653_),
    .C(_09654_),
    .A(_09652_),
    .Y(_09656_),
    .D(_09655_));
 sg13g2_a21oi_1 _15512_ (.A1(net732),
    .A2(net4678),
    .Y(_09657_),
    .B1(_09656_));
 sg13g2_nor2_2 _15513_ (.A(net4082),
    .B(_09657_),
    .Y(_09658_));
 sg13g2_a21o_1 _15514_ (.A2(net2905),
    .A1(net4895),
    .B1(_09658_),
    .X(_01040_));
 sg13g2_nand2_1 _15515_ (.Y(_09659_),
    .A(\soc_inst.cpu_core.register_file.registers[9][4] ),
    .B(net4577));
 sg13g2_a22oi_1 _15516_ (.Y(_09660_),
    .B1(net4562),
    .B2(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .A2(net4592),
    .A1(\soc_inst.cpu_core.register_file.registers[13][4] ));
 sg13g2_a21oi_1 _15517_ (.A1(\soc_inst.cpu_core.register_file.registers[14][4] ),
    .A2(net4572),
    .Y(_09661_),
    .B1(net4679));
 sg13g2_a22oi_1 _15518_ (.Y(_09662_),
    .B1(net4547),
    .B2(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .A2(net4552),
    .A1(\soc_inst.cpu_core.register_file.registers[6][4] ));
 sg13g2_a22oi_1 _15519_ (.Y(_09663_),
    .B1(net4532),
    .B2(\soc_inst.cpu_core.register_file.registers[11][4] ),
    .A2(net4542),
    .A1(\soc_inst.cpu_core.register_file.registers[15][4] ));
 sg13g2_nand3_1 _15520_ (.B(_09662_),
    .C(_09663_),
    .A(_09661_),
    .Y(_09664_));
 sg13g2_a221oi_1 _15521_ (.B2(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .C1(_09664_),
    .B1(net4537),
    .A1(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .Y(_09665_),
    .A2(net4557));
 sg13g2_a22oi_1 _15522_ (.Y(_09666_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][4] ));
 sg13g2_nand3_1 _15523_ (.B(_09660_),
    .C(_09666_),
    .A(_09659_),
    .Y(_09667_));
 sg13g2_a221oi_1 _15524_ (.B2(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .C1(_09667_),
    .B1(net4567),
    .A1(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .Y(_09668_),
    .A2(net4582));
 sg13g2_a221oi_1 _15525_ (.B2(_09668_),
    .C1(net4083),
    .B1(_09665_),
    .A1(_05723_),
    .Y(_09669_),
    .A2(net4680));
 sg13g2_a21o_1 _15526_ (.A2(net2829),
    .A1(net4891),
    .B1(_09669_),
    .X(_01041_));
 sg13g2_nand2_1 _15527_ (.Y(_09670_),
    .A(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .B(net4537));
 sg13g2_a22oi_1 _15528_ (.Y(_09671_),
    .B1(net4581),
    .B2(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][5] ));
 sg13g2_a21oi_1 _15529_ (.A1(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .A2(net4562),
    .Y(_09672_),
    .B1(net4680));
 sg13g2_a22oi_1 _15530_ (.Y(_09673_),
    .B1(net4566),
    .B2(\soc_inst.cpu_core.register_file.registers[3][5] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][5] ));
 sg13g2_a22oi_1 _15531_ (.Y(_09674_),
    .B1(net4546),
    .B2(\soc_inst.cpu_core.register_file.registers[2][5] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][5] ));
 sg13g2_nand4_1 _15532_ (.B(_09672_),
    .C(_09673_),
    .A(_09671_),
    .Y(_09675_),
    .D(_09674_));
 sg13g2_a22oi_1 _15533_ (.Y(_09676_),
    .B1(net4552),
    .B2(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .A2(net4572),
    .A1(\soc_inst.cpu_core.register_file.registers[14][5] ));
 sg13g2_a22oi_1 _15534_ (.Y(_09677_),
    .B1(net4542),
    .B2(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .A2(net4557),
    .A1(\soc_inst.cpu_core.register_file.registers[12][5] ));
 sg13g2_a22oi_1 _15535_ (.Y(_09678_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .A2(net4532),
    .A1(\soc_inst.cpu_core.register_file.registers[11][5] ));
 sg13g2_nand4_1 _15536_ (.B(_09676_),
    .C(_09677_),
    .A(_09670_),
    .Y(_09679_),
    .D(_09678_));
 sg13g2_nor2_2 _15537_ (.A(_09675_),
    .B(_09679_),
    .Y(_09680_));
 sg13g2_nor2_1 _15538_ (.A(net879),
    .B(_09593_),
    .Y(_09681_));
 sg13g2_nor3_2 _15539_ (.A(net4083),
    .B(_09680_),
    .C(_09681_),
    .Y(_09682_));
 sg13g2_a21o_1 _15540_ (.A2(net2914),
    .A1(net4889),
    .B1(_09682_),
    .X(_01042_));
 sg13g2_nand2_1 _15541_ (.Y(_09683_),
    .A(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .B(net4542));
 sg13g2_a22oi_1 _15542_ (.Y(_09684_),
    .B1(net4552),
    .B2(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .A2(net4557),
    .A1(\soc_inst.cpu_core.register_file.registers[12][6] ));
 sg13g2_a21oi_1 _15543_ (.A1(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .A2(net4582),
    .Y(_09685_),
    .B1(net4680));
 sg13g2_a22oi_1 _15544_ (.Y(_09686_),
    .B1(net4547),
    .B2(\soc_inst.cpu_core.register_file.registers[2][6] ),
    .A2(net4592),
    .A1(\soc_inst.cpu_core.register_file.registers[13][6] ));
 sg13g2_a22oi_1 _15545_ (.Y(_09687_),
    .B1(net4537),
    .B2(\soc_inst.cpu_core.register_file.registers[10][6] ),
    .A2(net4562),
    .A1(\soc_inst.cpu_core.register_file.registers[7][6] ));
 sg13g2_a22oi_1 _15546_ (.Y(_09688_),
    .B1(net4567),
    .B2(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .A2(net4577),
    .A1(\soc_inst.cpu_core.register_file.registers[9][6] ));
 sg13g2_nand4_1 _15547_ (.B(_09686_),
    .C(_09687_),
    .A(_09685_),
    .Y(_09689_),
    .D(_09688_));
 sg13g2_a22oi_1 _15548_ (.Y(_09690_),
    .B1(net4532),
    .B2(\soc_inst.cpu_core.register_file.registers[11][6] ),
    .A2(net4572),
    .A1(\soc_inst.cpu_core.register_file.registers[14][6] ));
 sg13g2_a22oi_1 _15549_ (.Y(_09691_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][6] ));
 sg13g2_nand4_1 _15550_ (.B(_09684_),
    .C(_09690_),
    .A(_09683_),
    .Y(_09692_),
    .D(_09691_));
 sg13g2_nor2_2 _15551_ (.A(_09689_),
    .B(_09692_),
    .Y(_09693_));
 sg13g2_nor2_1 _15552_ (.A(net1267),
    .B(_09593_),
    .Y(_09694_));
 sg13g2_nor3_2 _15553_ (.A(net4083),
    .B(_09693_),
    .C(_09694_),
    .Y(_09695_));
 sg13g2_a21o_1 _15554_ (.A2(net2734),
    .A1(net4891),
    .B1(_09695_),
    .X(_01043_));
 sg13g2_a22oi_1 _15555_ (.Y(_09696_),
    .B1(net4561),
    .B2(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][7] ));
 sg13g2_a22oi_1 _15556_ (.Y(_09697_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][7] ),
    .A2(net4551),
    .A1(\soc_inst.cpu_core.register_file.registers[6][7] ));
 sg13g2_a22oi_1 _15557_ (.Y(_09698_),
    .B1(net4546),
    .B2(\soc_inst.cpu_core.register_file.registers[2][7] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][7] ));
 sg13g2_nand3_1 _15558_ (.B(_09697_),
    .C(_09698_),
    .A(_09696_),
    .Y(_09699_));
 sg13g2_a221oi_1 _15559_ (.B2(\soc_inst.cpu_core.register_file.registers[10][7] ),
    .C1(_09699_),
    .B1(net4536),
    .A1(\soc_inst.cpu_core.register_file.registers[12][7] ),
    .Y(_09700_),
    .A2(net4556));
 sg13g2_a22oi_1 _15560_ (.Y(_09701_),
    .B1(net4541),
    .B2(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .A2(net4566),
    .A1(\soc_inst.cpu_core.register_file.registers[3][7] ));
 sg13g2_a22oi_1 _15561_ (.Y(_09702_),
    .B1(net4571),
    .B2(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .A2(net4581),
    .A1(\soc_inst.cpu_core.register_file.registers[5][7] ));
 sg13g2_a22oi_1 _15562_ (.Y(_09703_),
    .B1(net4531),
    .B2(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][7] ));
 sg13g2_nand4_1 _15563_ (.B(_09701_),
    .C(_09702_),
    .A(_09700_),
    .Y(_09704_),
    .D(_09703_));
 sg13g2_a21oi_2 _15564_ (.B1(_09704_),
    .Y(_09705_),
    .A2(net4678),
    .A1(net2016));
 sg13g2_nor2_2 _15565_ (.A(net4084),
    .B(_09705_),
    .Y(_09706_));
 sg13g2_a21o_1 _15566_ (.A2(net2866),
    .A1(net4889),
    .B1(_09706_),
    .X(_01044_));
 sg13g2_a22oi_1 _15567_ (.Y(_09707_),
    .B1(net4529),
    .B2(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .A2(net4554),
    .A1(\soc_inst.cpu_core.register_file.registers[12][8] ));
 sg13g2_a22oi_1 _15568_ (.Y(_09708_),
    .B1(net4569),
    .B2(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][8] ));
 sg13g2_a22oi_1 _15569_ (.Y(_09709_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .A2(net4559),
    .A1(\soc_inst.cpu_core.register_file.registers[7][8] ));
 sg13g2_nand3_1 _15570_ (.B(_09708_),
    .C(_09709_),
    .A(_09707_),
    .Y(_09710_));
 sg13g2_a221oi_1 _15571_ (.B2(\soc_inst.cpu_core.register_file.registers[10][8] ),
    .C1(_09710_),
    .B1(net4534),
    .A1(\soc_inst.cpu_core.register_file.registers[4][8] ),
    .Y(_09711_),
    .A2(net4584));
 sg13g2_a22oi_1 _15572_ (.Y(_09712_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][8] ));
 sg13g2_a22oi_1 _15573_ (.Y(_09713_),
    .B1(net4549),
    .B2(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .A2(net4574),
    .A1(\soc_inst.cpu_core.register_file.registers[9][8] ));
 sg13g2_a22oi_1 _15574_ (.Y(_09714_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][8] ),
    .A2(net4589),
    .A1(\soc_inst.cpu_core.register_file.registers[13][8] ));
 sg13g2_nand4_1 _15575_ (.B(_09712_),
    .C(_09713_),
    .A(_09711_),
    .Y(_09715_),
    .D(_09714_));
 sg13g2_a21oi_1 _15576_ (.A1(net1594),
    .A2(net4677),
    .Y(_09716_),
    .B1(_09715_));
 sg13g2_nor2_2 _15577_ (.A(net4082),
    .B(_09716_),
    .Y(_09717_));
 sg13g2_a21o_1 _15578_ (.A2(net2850),
    .A1(net4892),
    .B1(_09717_),
    .X(_01045_));
 sg13g2_a22oi_1 _15579_ (.Y(_09718_),
    .B1(net4532),
    .B2(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][9] ));
 sg13g2_nand2_1 _15580_ (.Y(_09719_),
    .A(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .B(net4567));
 sg13g2_a22oi_1 _15581_ (.Y(_09720_),
    .B1(net4542),
    .B2(\soc_inst.cpu_core.register_file.registers[15][9] ),
    .A2(net4592),
    .A1(\soc_inst.cpu_core.register_file.registers[13][9] ));
 sg13g2_a21oi_1 _15582_ (.A1(\soc_inst.cpu_core.register_file.registers[5][9] ),
    .A2(net4582),
    .Y(_09721_),
    .B1(net4679));
 sg13g2_a22oi_1 _15583_ (.Y(_09722_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .A2(net4537),
    .A1(\soc_inst.cpu_core.register_file.registers[10][9] ));
 sg13g2_nand3_1 _15584_ (.B(_09721_),
    .C(_09722_),
    .A(_09718_),
    .Y(_09723_));
 sg13g2_a221oi_1 _15585_ (.B2(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .C1(_09723_),
    .B1(net4547),
    .A1(\soc_inst.cpu_core.register_file.registers[12][9] ),
    .Y(_09724_),
    .A2(net4557));
 sg13g2_a22oi_1 _15586_ (.Y(_09725_),
    .B1(net4552),
    .B2(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .A2(net4562),
    .A1(\soc_inst.cpu_core.register_file.registers[7][9] ));
 sg13g2_nand3_1 _15587_ (.B(_09720_),
    .C(_09725_),
    .A(_09719_),
    .Y(_09726_));
 sg13g2_a221oi_1 _15588_ (.B2(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .C1(_09726_),
    .B1(net4572),
    .A1(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .Y(_09727_),
    .A2(net4577));
 sg13g2_a221oi_1 _15589_ (.B2(_09727_),
    .C1(net4083),
    .B1(_09724_),
    .A1(_05724_),
    .Y(_09728_),
    .A2(net4679));
 sg13g2_a21o_1 _15590_ (.A2(net2822),
    .A1(net4892),
    .B1(_09728_),
    .X(_01046_));
 sg13g2_a22oi_1 _15591_ (.Y(_09729_),
    .B1(net4561),
    .B2(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][10] ));
 sg13g2_a22oi_1 _15592_ (.Y(_09730_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][10] ));
 sg13g2_a22oi_1 _15593_ (.Y(_09731_),
    .B1(net4541),
    .B2(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .A2(net4556),
    .A1(\soc_inst.cpu_core.register_file.registers[12][10] ));
 sg13g2_a22oi_1 _15594_ (.Y(_09732_),
    .B1(net4536),
    .B2(\soc_inst.cpu_core.register_file.registers[10][10] ),
    .A2(net4551),
    .A1(\soc_inst.cpu_core.register_file.registers[6][10] ));
 sg13g2_nand3_1 _15595_ (.B(_09731_),
    .C(_09732_),
    .A(_09730_),
    .Y(_09733_));
 sg13g2_a221oi_1 _15596_ (.B2(\soc_inst.cpu_core.register_file.registers[11][10] ),
    .C1(_09733_),
    .B1(net4531),
    .A1(\soc_inst.cpu_core.register_file.registers[2][10] ),
    .Y(_09734_),
    .A2(net4546));
 sg13g2_a22oi_1 _15597_ (.Y(_09735_),
    .B1(net4571),
    .B2(\soc_inst.cpu_core.register_file.registers[14][10] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][10] ));
 sg13g2_a22oi_1 _15598_ (.Y(_09736_),
    .B1(net4566),
    .B2(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .A2(net4581),
    .A1(\soc_inst.cpu_core.register_file.registers[5][10] ));
 sg13g2_nand4_1 _15599_ (.B(_09734_),
    .C(_09735_),
    .A(_09729_),
    .Y(_09737_),
    .D(_09736_));
 sg13g2_a21oi_1 _15600_ (.A1(net1171),
    .A2(net4678),
    .Y(_09738_),
    .B1(_09737_));
 sg13g2_nor2_2 _15601_ (.A(net4082),
    .B(_09738_),
    .Y(_09739_));
 sg13g2_a21o_1 _15602_ (.A2(net2550),
    .A1(net4892),
    .B1(_09739_),
    .X(_01047_));
 sg13g2_a22oi_1 _15603_ (.Y(_09740_),
    .B1(net4536),
    .B2(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .A2(net4571),
    .A1(\soc_inst.cpu_core.register_file.registers[14][11] ));
 sg13g2_a22oi_1 _15604_ (.Y(_09741_),
    .B1(net4541),
    .B2(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .A2(net4556),
    .A1(\soc_inst.cpu_core.register_file.registers[12][11] ));
 sg13g2_a22oi_1 _15605_ (.Y(_09742_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][11] ),
    .A2(net4592),
    .A1(\soc_inst.cpu_core.register_file.registers[13][11] ));
 sg13g2_nand3_1 _15606_ (.B(_09741_),
    .C(_09742_),
    .A(_09740_),
    .Y(_09743_));
 sg13g2_a221oi_1 _15607_ (.B2(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .C1(_09743_),
    .B1(net4561),
    .A1(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .Y(_09744_),
    .A2(net4581));
 sg13g2_a22oi_1 _15608_ (.Y(_09745_),
    .B1(net4546),
    .B2(\soc_inst.cpu_core.register_file.registers[2][11] ),
    .A2(net4586),
    .A1(\soc_inst.cpu_core.register_file.registers[4][11] ));
 sg13g2_a22oi_1 _15609_ (.Y(_09746_),
    .B1(net4531),
    .B2(\soc_inst.cpu_core.register_file.registers[11][11] ),
    .A2(net4566),
    .A1(\soc_inst.cpu_core.register_file.registers[3][11] ));
 sg13g2_a22oi_1 _15610_ (.Y(_09747_),
    .B1(net4551),
    .B2(\soc_inst.cpu_core.register_file.registers[6][11] ),
    .A2(net4577),
    .A1(\soc_inst.cpu_core.register_file.registers[9][11] ));
 sg13g2_nand4_1 _15611_ (.B(_09745_),
    .C(_09746_),
    .A(_09744_),
    .Y(_09748_),
    .D(_09747_));
 sg13g2_a21oi_2 _15612_ (.B1(_09748_),
    .Y(_09749_),
    .A2(net4680),
    .A1(net1845));
 sg13g2_nor2_2 _15613_ (.A(net4084),
    .B(_09749_),
    .Y(_09750_));
 sg13g2_a21o_1 _15614_ (.A2(net764),
    .A1(net4891),
    .B1(_09750_),
    .X(_01048_));
 sg13g2_a22oi_1 _15615_ (.Y(_09751_),
    .B1(net4542),
    .B2(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .A2(net4557),
    .A1(\soc_inst.cpu_core.register_file.registers[12][12] ));
 sg13g2_a22oi_1 _15616_ (.Y(_09752_),
    .B1(net4547),
    .B2(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .A2(net4552),
    .A1(\soc_inst.cpu_core.register_file.registers[6][12] ));
 sg13g2_a22oi_1 _15617_ (.Y(_09753_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .A2(net4592),
    .A1(\soc_inst.cpu_core.register_file.registers[13][12] ));
 sg13g2_nand3_1 _15618_ (.B(_09752_),
    .C(_09753_),
    .A(_09751_),
    .Y(_09754_));
 sg13g2_a221oi_1 _15619_ (.B2(\soc_inst.cpu_core.register_file.registers[11][12] ),
    .C1(_09754_),
    .B1(net4532),
    .A1(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .Y(_09755_),
    .A2(net4562));
 sg13g2_a22oi_1 _15620_ (.Y(_09756_),
    .B1(net4572),
    .B2(\soc_inst.cpu_core.register_file.registers[14][12] ),
    .A2(net4582),
    .A1(\soc_inst.cpu_core.register_file.registers[5][12] ));
 sg13g2_a22oi_1 _15621_ (.Y(_09757_),
    .B1(net4567),
    .B2(\soc_inst.cpu_core.register_file.registers[3][12] ),
    .A2(net4577),
    .A1(\soc_inst.cpu_core.register_file.registers[9][12] ));
 sg13g2_a22oi_1 _15622_ (.Y(_09758_),
    .B1(net4537),
    .B2(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][12] ));
 sg13g2_nand4_1 _15623_ (.B(_09756_),
    .C(_09757_),
    .A(_09755_),
    .Y(_09759_),
    .D(_09758_));
 sg13g2_a21oi_1 _15624_ (.A1(net1335),
    .A2(net4680),
    .Y(_09760_),
    .B1(_09759_));
 sg13g2_nor2_2 _15625_ (.A(net4083),
    .B(_09760_),
    .Y(_09761_));
 sg13g2_a21o_1 _15626_ (.A2(net2876),
    .A1(net4891),
    .B1(_09761_),
    .X(_01049_));
 sg13g2_a22oi_1 _15627_ (.Y(_09762_),
    .B1(net4529),
    .B2(\soc_inst.cpu_core.register_file.registers[11][13] ),
    .A2(net4559),
    .A1(\soc_inst.cpu_core.register_file.registers[7][13] ));
 sg13g2_a22oi_1 _15628_ (.Y(_09763_),
    .B1(net4574),
    .B2(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .A2(net4584),
    .A1(\soc_inst.cpu_core.register_file.registers[4][13] ));
 sg13g2_a22oi_1 _15629_ (.Y(_09764_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .A2(net4539),
    .A1(\soc_inst.cpu_core.register_file.registers[15][13] ));
 sg13g2_a22oi_1 _15630_ (.Y(_09765_),
    .B1(net4534),
    .B2(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][13] ));
 sg13g2_nand3_1 _15631_ (.B(_09764_),
    .C(_09765_),
    .A(_09763_),
    .Y(_09766_));
 sg13g2_a221oi_1 _15632_ (.B2(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .C1(_09766_),
    .B1(net4569),
    .A1(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .Y(_09767_),
    .A2(net4589));
 sg13g2_a22oi_1 _15633_ (.Y(_09768_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .A2(net4554),
    .A1(\soc_inst.cpu_core.register_file.registers[12][13] ));
 sg13g2_a22oi_1 _15634_ (.Y(_09769_),
    .B1(net4549),
    .B2(\soc_inst.cpu_core.register_file.registers[6][13] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][13] ));
 sg13g2_nand4_1 _15635_ (.B(_09767_),
    .C(_09768_),
    .A(_09762_),
    .Y(_09770_),
    .D(_09769_));
 sg13g2_a21oi_1 _15636_ (.A1(net715),
    .A2(net4677),
    .Y(_09771_),
    .B1(_09770_));
 sg13g2_nor2_2 _15637_ (.A(net4080),
    .B(_09771_),
    .Y(_09772_));
 sg13g2_a21o_1 _15638_ (.A2(net2915),
    .A1(net4880),
    .B1(_09772_),
    .X(_01050_));
 sg13g2_nand2_1 _15639_ (.Y(_09773_),
    .A(\soc_inst.cpu_core.register_file.registers[3][14] ),
    .B(net4567));
 sg13g2_a21oi_1 _15640_ (.A1(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .A2(net4562),
    .Y(_09774_),
    .B1(net4679));
 sg13g2_a22oi_1 _15641_ (.Y(_09775_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][14] ));
 sg13g2_a22oi_1 _15642_ (.Y(_09776_),
    .B1(net4547),
    .B2(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .A2(net4577),
    .A1(\soc_inst.cpu_core.register_file.registers[9][14] ));
 sg13g2_nand3_1 _15643_ (.B(_09775_),
    .C(_09776_),
    .A(_09774_),
    .Y(_09777_));
 sg13g2_a221oi_1 _15644_ (.B2(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .C1(_09777_),
    .B1(net4582),
    .A1(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .Y(_09778_),
    .A2(net4592));
 sg13g2_a22oi_1 _15645_ (.Y(_09779_),
    .B1(net4537),
    .B2(\soc_inst.cpu_core.register_file.registers[10][14] ),
    .A2(net4572),
    .A1(\soc_inst.cpu_core.register_file.registers[14][14] ));
 sg13g2_a22oi_1 _15646_ (.Y(_09780_),
    .B1(net4532),
    .B2(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .A2(net4557),
    .A1(\soc_inst.cpu_core.register_file.registers[12][14] ));
 sg13g2_nand3_1 _15647_ (.B(_09779_),
    .C(_09780_),
    .A(_09773_),
    .Y(_09781_));
 sg13g2_a221oi_1 _15648_ (.B2(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .C1(_09781_),
    .B1(net4542),
    .A1(\soc_inst.cpu_core.register_file.registers[6][14] ),
    .Y(_09782_),
    .A2(net4552));
 sg13g2_a221oi_1 _15649_ (.B2(_09782_),
    .C1(net4084),
    .B1(_09778_),
    .A1(_05726_),
    .Y(_09783_),
    .A2(net4679));
 sg13g2_a21o_1 _15650_ (.A2(net2551),
    .A1(net4902),
    .B1(_09783_),
    .X(_01051_));
 sg13g2_nand2_1 _15651_ (.Y(_09784_),
    .A(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .B(net4525));
 sg13g2_a21oi_1 _15652_ (.A1(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .A2(net4560),
    .Y(_09785_),
    .B1(net4676));
 sg13g2_a22oi_1 _15653_ (.Y(_09786_),
    .B1(net4530),
    .B2(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .A2(net4545),
    .A1(\soc_inst.cpu_core.register_file.registers[2][15] ));
 sg13g2_a22oi_1 _15654_ (.Y(_09787_),
    .B1(net4535),
    .B2(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][15] ));
 sg13g2_nand3_1 _15655_ (.B(_09786_),
    .C(_09787_),
    .A(_09785_),
    .Y(_09788_));
 sg13g2_a221oi_1 _15656_ (.B2(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .C1(_09788_),
    .B1(net4550),
    .A1(\soc_inst.cpu_core.register_file.registers[12][15] ),
    .Y(_09789_),
    .A2(net4555));
 sg13g2_a22oi_1 _15657_ (.Y(_09790_),
    .B1(net4565),
    .B2(\soc_inst.cpu_core.register_file.registers[3][15] ),
    .A2(net4590),
    .A1(\soc_inst.cpu_core.register_file.registers[13][15] ));
 sg13g2_a22oi_1 _15658_ (.Y(_09791_),
    .B1(net4540),
    .B2(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .A2(net4570),
    .A1(\soc_inst.cpu_core.register_file.registers[14][15] ));
 sg13g2_nand3_1 _15659_ (.B(_09790_),
    .C(_09791_),
    .A(_09784_),
    .Y(_09792_));
 sg13g2_a221oi_1 _15660_ (.B2(\soc_inst.cpu_core.register_file.registers[5][15] ),
    .C1(_09792_),
    .B1(net4580),
    .A1(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .Y(_09793_),
    .A2(net4585));
 sg13g2_a221oi_1 _15661_ (.B2(_09793_),
    .C1(net4080),
    .B1(_09789_),
    .A1(_05727_),
    .Y(_09794_),
    .A2(net4676));
 sg13g2_a21o_1 _15662_ (.A2(net2865),
    .A1(net4902),
    .B1(_09794_),
    .X(_01052_));
 sg13g2_a22oi_1 _15663_ (.Y(_09795_),
    .B1(net4574),
    .B2(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][16] ));
 sg13g2_a22oi_1 _15664_ (.Y(_09796_),
    .B1(net4534),
    .B2(\soc_inst.cpu_core.register_file.registers[10][16] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][16] ));
 sg13g2_a22oi_1 _15665_ (.Y(_09797_),
    .B1(net4559),
    .B2(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .A2(net4569),
    .A1(\soc_inst.cpu_core.register_file.registers[14][16] ));
 sg13g2_a22oi_1 _15666_ (.Y(_09798_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .A2(net4584),
    .A1(\soc_inst.cpu_core.register_file.registers[4][16] ));
 sg13g2_nand3_1 _15667_ (.B(_09797_),
    .C(_09798_),
    .A(_09796_),
    .Y(_09799_));
 sg13g2_a221oi_1 _15668_ (.B2(\soc_inst.cpu_core.register_file.registers[11][16] ),
    .C1(_09799_),
    .B1(net4529),
    .A1(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .Y(_09800_),
    .A2(net4589));
 sg13g2_a22oi_1 _15669_ (.Y(_09801_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][16] ),
    .A2(net4549),
    .A1(\soc_inst.cpu_core.register_file.registers[6][16] ));
 sg13g2_a22oi_1 _15670_ (.Y(_09802_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][16] ),
    .A2(net4554),
    .A1(\soc_inst.cpu_core.register_file.registers[12][16] ));
 sg13g2_nand4_1 _15671_ (.B(_09800_),
    .C(_09801_),
    .A(_09795_),
    .Y(_09803_),
    .D(_09802_));
 sg13g2_a21oi_1 _15672_ (.A1(net1027),
    .A2(net4675),
    .Y(_09804_),
    .B1(_09803_));
 sg13g2_nor2_2 _15673_ (.A(net4080),
    .B(_09804_),
    .Y(_09805_));
 sg13g2_a21o_1 _15674_ (.A2(net1516),
    .A1(net4883),
    .B1(_09805_),
    .X(_01053_));
 sg13g2_nand2_1 _15675_ (.Y(_09806_),
    .A(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .B(net4540));
 sg13g2_a22oi_1 _15676_ (.Y(_09807_),
    .B1(net4535),
    .B2(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .A2(net4545),
    .A1(\soc_inst.cpu_core.register_file.registers[2][17] ));
 sg13g2_a21oi_1 _15677_ (.A1(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .A2(net4560),
    .Y(_09808_),
    .B1(net4676));
 sg13g2_a22oi_1 _15678_ (.Y(_09809_),
    .B1(net4525),
    .B2(\soc_inst.cpu_core.register_file.registers[8][17] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][17] ));
 sg13g2_nand3_1 _15679_ (.B(_09808_),
    .C(_09809_),
    .A(_09807_),
    .Y(_09810_));
 sg13g2_a221oi_1 _15680_ (.B2(\soc_inst.cpu_core.register_file.registers[5][17] ),
    .C1(_09810_),
    .B1(net4580),
    .A1(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .Y(_09811_),
    .A2(net4590));
 sg13g2_a22oi_1 _15681_ (.Y(_09812_),
    .B1(net4550),
    .B2(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .A2(net4585),
    .A1(\soc_inst.cpu_core.register_file.registers[4][17] ));
 sg13g2_a22oi_1 _15682_ (.Y(_09813_),
    .B1(net4555),
    .B2(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .A2(net4565),
    .A1(\soc_inst.cpu_core.register_file.registers[3][17] ));
 sg13g2_nand3_1 _15683_ (.B(_09812_),
    .C(_09813_),
    .A(_09806_),
    .Y(_09814_));
 sg13g2_a221oi_1 _15684_ (.B2(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .C1(_09814_),
    .B1(net4530),
    .A1(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .Y(_09815_),
    .A2(net4570));
 sg13g2_a221oi_1 _15685_ (.B2(_09815_),
    .C1(net4081),
    .B1(_09811_),
    .A1(_05728_),
    .Y(_09816_),
    .A2(net4676));
 sg13g2_a21o_1 _15686_ (.A2(net2339),
    .A1(net4900),
    .B1(_09816_),
    .X(_01054_));
 sg13g2_a22oi_1 _15687_ (.Y(_09817_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .A2(net4529),
    .A1(\soc_inst.cpu_core.register_file.registers[11][18] ));
 sg13g2_a22oi_1 _15688_ (.Y(_09818_),
    .B1(net4549),
    .B2(\soc_inst.cpu_core.register_file.registers[6][18] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][18] ));
 sg13g2_a22oi_1 _15689_ (.Y(_09819_),
    .B1(net4534),
    .B2(\soc_inst.cpu_core.register_file.registers[10][18] ),
    .A2(net4584),
    .A1(\soc_inst.cpu_core.register_file.registers[4][18] ));
 sg13g2_nand3_1 _15690_ (.B(_09818_),
    .C(_09819_),
    .A(_09817_),
    .Y(_09820_));
 sg13g2_a221oi_1 _15691_ (.B2(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .C1(_09820_),
    .B1(net4559),
    .A1(\soc_inst.cpu_core.register_file.registers[9][18] ),
    .Y(_09821_),
    .A2(net4574));
 sg13g2_a22oi_1 _15692_ (.Y(_09822_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .A2(net4589),
    .A1(\soc_inst.cpu_core.register_file.registers[13][18] ));
 sg13g2_a22oi_1 _15693_ (.Y(_09823_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .A2(net4569),
    .A1(\soc_inst.cpu_core.register_file.registers[14][18] ));
 sg13g2_a22oi_1 _15694_ (.Y(_09824_),
    .B1(net4554),
    .B2(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][18] ));
 sg13g2_nand4_1 _15695_ (.B(_09822_),
    .C(_09823_),
    .A(_09821_),
    .Y(_09825_),
    .D(_09824_));
 sg13g2_a21oi_1 _15696_ (.A1(net723),
    .A2(net4675),
    .Y(_09826_),
    .B1(_09825_));
 sg13g2_nor2_2 _15697_ (.A(net4080),
    .B(_09826_),
    .Y(_09827_));
 sg13g2_a21o_1 _15698_ (.A2(net2797),
    .A1(net4882),
    .B1(_09827_),
    .X(_01055_));
 sg13g2_nand2_1 _15699_ (.Y(_09828_),
    .A(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .B(net4540));
 sg13g2_a22oi_1 _15700_ (.Y(_09829_),
    .B1(net4550),
    .B2(\soc_inst.cpu_core.register_file.registers[6][19] ),
    .A2(net4590),
    .A1(\soc_inst.cpu_core.register_file.registers[13][19] ));
 sg13g2_a21oi_1 _15701_ (.A1(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .A2(net4580),
    .Y(_09830_),
    .B1(net4675));
 sg13g2_a22oi_1 _15702_ (.Y(_09831_),
    .B1(net4535),
    .B2(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][19] ));
 sg13g2_a22oi_1 _15703_ (.Y(_09832_),
    .B1(net4555),
    .B2(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .A2(net4565),
    .A1(\soc_inst.cpu_core.register_file.registers[3][19] ));
 sg13g2_nand4_1 _15704_ (.B(_09830_),
    .C(_09831_),
    .A(_09829_),
    .Y(_09833_),
    .D(_09832_));
 sg13g2_a22oi_1 _15705_ (.Y(_09834_),
    .B1(net4525),
    .B2(\soc_inst.cpu_core.register_file.registers[8][19] ),
    .A2(net4585),
    .A1(\soc_inst.cpu_core.register_file.registers[4][19] ));
 sg13g2_a22oi_1 _15706_ (.Y(_09835_),
    .B1(net4545),
    .B2(\soc_inst.cpu_core.register_file.registers[2][19] ),
    .A2(net4560),
    .A1(\soc_inst.cpu_core.register_file.registers[7][19] ));
 sg13g2_a22oi_1 _15707_ (.Y(_09836_),
    .B1(net4530),
    .B2(\soc_inst.cpu_core.register_file.registers[11][19] ),
    .A2(net4570),
    .A1(\soc_inst.cpu_core.register_file.registers[14][19] ));
 sg13g2_nand4_1 _15708_ (.B(_09834_),
    .C(_09835_),
    .A(_09828_),
    .Y(_09837_),
    .D(_09836_));
 sg13g2_nor2_1 _15709_ (.A(_09833_),
    .B(_09837_),
    .Y(_09838_));
 sg13g2_nor2_1 _15710_ (.A(net768),
    .B(_09593_),
    .Y(_09839_));
 sg13g2_nor3_2 _15711_ (.A(net4080),
    .B(_09838_),
    .C(_09839_),
    .Y(_09840_));
 sg13g2_a21o_1 _15712_ (.A2(net2646),
    .A1(net4884),
    .B1(_09840_),
    .X(_01056_));
 sg13g2_a22oi_1 _15713_ (.Y(_09841_),
    .B1(net4559),
    .B2(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .A2(net4589),
    .A1(\soc_inst.cpu_core.register_file.registers[13][20] ));
 sg13g2_a22oi_1 _15714_ (.Y(_09842_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][20] ));
 sg13g2_a22oi_1 _15715_ (.Y(_09843_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][20] ));
 sg13g2_a22oi_1 _15716_ (.Y(_09844_),
    .B1(net4574),
    .B2(\soc_inst.cpu_core.register_file.registers[9][20] ),
    .A2(net4584),
    .A1(\soc_inst.cpu_core.register_file.registers[4][20] ));
 sg13g2_a22oi_1 _15717_ (.Y(_09845_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .A2(net4554),
    .A1(\soc_inst.cpu_core.register_file.registers[12][20] ));
 sg13g2_nand3_1 _15718_ (.B(_09844_),
    .C(_09845_),
    .A(_09843_),
    .Y(_09846_));
 sg13g2_a221oi_1 _15719_ (.B2(\soc_inst.cpu_core.register_file.registers[11][20] ),
    .C1(_09846_),
    .B1(net4529),
    .A1(\soc_inst.cpu_core.register_file.registers[14][20] ),
    .Y(_09847_),
    .A2(net4569));
 sg13g2_a22oi_1 _15720_ (.Y(_09848_),
    .B1(net4534),
    .B2(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .A2(net4549),
    .A1(\soc_inst.cpu_core.register_file.registers[6][20] ));
 sg13g2_nand4_1 _15721_ (.B(_09842_),
    .C(_09847_),
    .A(_09841_),
    .Y(_09849_),
    .D(_09848_));
 sg13g2_a21oi_1 _15722_ (.A1(net1278),
    .A2(net4675),
    .Y(_09850_),
    .B1(_09849_));
 sg13g2_nor2_2 _15723_ (.A(net4080),
    .B(_09850_),
    .Y(_09851_));
 sg13g2_a21o_1 _15724_ (.A2(net2823),
    .A1(net4884),
    .B1(_09851_),
    .X(_01057_));
 sg13g2_a22oi_1 _15725_ (.Y(_09852_),
    .B1(net4535),
    .B2(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .A2(net4545),
    .A1(\soc_inst.cpu_core.register_file.registers[2][21] ));
 sg13g2_nand2_1 _15726_ (.Y(_09853_),
    .A(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .B(net4565));
 sg13g2_a21oi_1 _15727_ (.A1(\soc_inst.cpu_core.register_file.registers[4][21] ),
    .A2(net4585),
    .Y(_09854_),
    .B1(net4676));
 sg13g2_a22oi_1 _15728_ (.Y(_09855_),
    .B1(net4570),
    .B2(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][21] ));
 sg13g2_a22oi_1 _15729_ (.Y(_09856_),
    .B1(net4560),
    .B2(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .A2(net4580),
    .A1(\soc_inst.cpu_core.register_file.registers[5][21] ));
 sg13g2_nand3_1 _15730_ (.B(_09855_),
    .C(_09856_),
    .A(_09854_),
    .Y(_09857_));
 sg13g2_a221oi_1 _15731_ (.B2(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .C1(_09857_),
    .B1(net4525),
    .A1(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .Y(_09858_),
    .A2(net4550));
 sg13g2_a22oi_1 _15732_ (.Y(_09859_),
    .B1(net4530),
    .B2(\soc_inst.cpu_core.register_file.registers[11][21] ),
    .A2(net4555),
    .A1(\soc_inst.cpu_core.register_file.registers[12][21] ));
 sg13g2_nand3_1 _15733_ (.B(_09853_),
    .C(_09859_),
    .A(_09852_),
    .Y(_09860_));
 sg13g2_a221oi_1 _15734_ (.B2(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .C1(_09860_),
    .B1(net4540),
    .A1(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .Y(_09861_),
    .A2(net4590));
 sg13g2_a221oi_1 _15735_ (.B2(_09861_),
    .C1(net4081),
    .B1(_09858_),
    .A1(_05729_),
    .Y(_09862_),
    .A2(net4676));
 sg13g2_a21o_1 _15736_ (.A2(net2639),
    .A1(net4883),
    .B1(_09862_),
    .X(_01058_));
 sg13g2_nand2_1 _15737_ (.Y(_09863_),
    .A(\soc_inst.cpu_core.register_file.registers[13][22] ),
    .B(net4590));
 sg13g2_a22oi_1 _15738_ (.Y(_09864_),
    .B1(net4550),
    .B2(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][22] ));
 sg13g2_a21oi_1 _15739_ (.A1(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .A2(net4535),
    .Y(_09865_),
    .B1(net4675));
 sg13g2_a22oi_1 _15740_ (.Y(_09866_),
    .B1(net4545),
    .B2(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .A2(net4555),
    .A1(\soc_inst.cpu_core.register_file.registers[12][22] ));
 sg13g2_a22oi_1 _15741_ (.Y(_09867_),
    .B1(net4560),
    .B2(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .A2(net4580),
    .A1(\soc_inst.cpu_core.register_file.registers[5][22] ));
 sg13g2_nand4_1 _15742_ (.B(_09865_),
    .C(_09866_),
    .A(_09864_),
    .Y(_09868_),
    .D(_09867_));
 sg13g2_a22oi_1 _15743_ (.Y(_09869_),
    .B1(net4540),
    .B2(\soc_inst.cpu_core.register_file.registers[15][22] ),
    .A2(net4570),
    .A1(\soc_inst.cpu_core.register_file.registers[14][22] ));
 sg13g2_a22oi_1 _15744_ (.Y(_09870_),
    .B1(net4530),
    .B2(\soc_inst.cpu_core.register_file.registers[11][22] ),
    .A2(net4565),
    .A1(\soc_inst.cpu_core.register_file.registers[3][22] ));
 sg13g2_a22oi_1 _15745_ (.Y(_09871_),
    .B1(net4525),
    .B2(\soc_inst.cpu_core.register_file.registers[8][22] ),
    .A2(net4585),
    .A1(\soc_inst.cpu_core.register_file.registers[4][22] ));
 sg13g2_nand4_1 _15746_ (.B(_09869_),
    .C(_09870_),
    .A(_09863_),
    .Y(_09872_),
    .D(_09871_));
 sg13g2_nor2_1 _15747_ (.A(_09868_),
    .B(_09872_),
    .Y(_09873_));
 sg13g2_nor2_1 _15748_ (.A(net769),
    .B(_09593_),
    .Y(_09874_));
 sg13g2_nor3_2 _15749_ (.A(net4081),
    .B(_09873_),
    .C(_09874_),
    .Y(_09875_));
 sg13g2_a21o_1 _15750_ (.A2(net2824),
    .A1(net4882),
    .B1(_09875_),
    .X(_01059_));
 sg13g2_a22oi_1 _15751_ (.Y(_09876_),
    .B1(net4569),
    .B2(\soc_inst.cpu_core.register_file.registers[14][23] ),
    .A2(net4584),
    .A1(\soc_inst.cpu_core.register_file.registers[4][23] ));
 sg13g2_a22oi_1 _15752_ (.Y(_09877_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .A2(net4589),
    .A1(\soc_inst.cpu_core.register_file.registers[13][23] ));
 sg13g2_a22oi_1 _15753_ (.Y(_09878_),
    .B1(net4549),
    .B2(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .A2(net4554),
    .A1(\soc_inst.cpu_core.register_file.registers[12][23] ));
 sg13g2_a22oi_1 _15754_ (.Y(_09879_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][23] ),
    .A2(net4574),
    .A1(\soc_inst.cpu_core.register_file.registers[9][23] ));
 sg13g2_nand3_1 _15755_ (.B(_09878_),
    .C(_09879_),
    .A(_09877_),
    .Y(_09880_));
 sg13g2_a221oi_1 _15756_ (.B2(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .C1(_09880_),
    .B1(net4559),
    .A1(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .Y(_09881_),
    .A2(net4579));
 sg13g2_a22oi_1 _15757_ (.Y(_09882_),
    .B1(net4529),
    .B2(\soc_inst.cpu_core.register_file.registers[11][23] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][23] ));
 sg13g2_a22oi_1 _15758_ (.Y(_09883_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][23] ),
    .A2(net4534),
    .A1(\soc_inst.cpu_core.register_file.registers[10][23] ));
 sg13g2_nand4_1 _15759_ (.B(_09881_),
    .C(_09882_),
    .A(_09876_),
    .Y(_09884_),
    .D(_09883_));
 sg13g2_a21oi_1 _15760_ (.A1(net739),
    .A2(net4675),
    .Y(_09885_),
    .B1(_09884_));
 sg13g2_nor2_2 _15761_ (.A(net4080),
    .B(_09885_),
    .Y(_09886_));
 sg13g2_a21o_1 _15762_ (.A2(net2753),
    .A1(net4882),
    .B1(_09886_),
    .X(_01060_));
 sg13g2_nand2_1 _15763_ (.Y(_09887_),
    .A(\soc_inst.cpu_core.register_file.registers[5][24] ),
    .B(net4583));
 sg13g2_a21oi_1 _15764_ (.A1(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .A2(net4530),
    .Y(_09888_),
    .B1(net4678));
 sg13g2_a22oi_1 _15765_ (.Y(_09889_),
    .B1(net4545),
    .B2(\soc_inst.cpu_core.register_file.registers[2][24] ),
    .A2(net4560),
    .A1(\soc_inst.cpu_core.register_file.registers[7][24] ));
 sg13g2_a22oi_1 _15766_ (.Y(_09890_),
    .B1(net4525),
    .B2(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .A2(net4535),
    .A1(\soc_inst.cpu_core.register_file.registers[10][24] ));
 sg13g2_nand3_1 _15767_ (.B(_09889_),
    .C(_09890_),
    .A(_09888_),
    .Y(_09891_));
 sg13g2_a221oi_1 _15768_ (.B2(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .C1(_09891_),
    .B1(net4550),
    .A1(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .Y(_09892_),
    .A2(net4590));
 sg13g2_a22oi_1 _15769_ (.Y(_09893_),
    .B1(net4570),
    .B2(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .A2(net4585),
    .A1(\soc_inst.cpu_core.register_file.registers[4][24] ));
 sg13g2_a22oi_1 _15770_ (.Y(_09894_),
    .B1(net4555),
    .B2(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][24] ));
 sg13g2_nand3_1 _15771_ (.B(_09893_),
    .C(_09894_),
    .A(_09887_),
    .Y(_09895_));
 sg13g2_a221oi_1 _15772_ (.B2(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .C1(_09895_),
    .B1(net4540),
    .A1(\soc_inst.cpu_core.register_file.registers[3][24] ),
    .Y(_09896_),
    .A2(net4565));
 sg13g2_a221oi_1 _15773_ (.B2(_09896_),
    .C1(net4082),
    .B1(_09892_),
    .A1(_05730_),
    .Y(_09897_),
    .A2(net4679));
 sg13g2_a21o_1 _15774_ (.A2(net1393),
    .A1(net4903),
    .B1(_09897_),
    .X(_01061_));
 sg13g2_a22oi_1 _15775_ (.Y(_09898_),
    .B1(net4577),
    .B2(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .A2(net4593),
    .A1(\soc_inst.cpu_core.register_file.registers[13][25] ));
 sg13g2_nand2_1 _15776_ (.Y(_09899_),
    .A(\soc_inst.cpu_core.register_file.registers[10][25] ),
    .B(net4537));
 sg13g2_a21oi_1 _15777_ (.A1(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .A2(net4527),
    .Y(_09900_),
    .B1(net4679));
 sg13g2_a22oi_1 _15778_ (.Y(_09901_),
    .B1(net4542),
    .B2(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][25] ));
 sg13g2_a22oi_1 _15779_ (.Y(_09902_),
    .B1(net4557),
    .B2(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .A2(net4562),
    .A1(\soc_inst.cpu_core.register_file.registers[7][25] ));
 sg13g2_and4_1 _15780_ (.A(_09898_),
    .B(_09900_),
    .C(_09901_),
    .D(_09902_),
    .X(_09903_));
 sg13g2_a22oi_1 _15781_ (.Y(_09904_),
    .B1(net4567),
    .B2(\soc_inst.cpu_core.register_file.registers[3][25] ),
    .A2(net4572),
    .A1(\soc_inst.cpu_core.register_file.registers[14][25] ));
 sg13g2_a22oi_1 _15782_ (.Y(_09905_),
    .B1(net4547),
    .B2(\soc_inst.cpu_core.register_file.registers[2][25] ),
    .A2(net4582),
    .A1(\soc_inst.cpu_core.register_file.registers[5][25] ));
 sg13g2_nand3_1 _15783_ (.B(_09904_),
    .C(_09905_),
    .A(_09899_),
    .Y(_09906_));
 sg13g2_a221oi_1 _15784_ (.B2(\soc_inst.cpu_core.register_file.registers[11][25] ),
    .C1(_09906_),
    .B1(net4532),
    .A1(\soc_inst.cpu_core.register_file.registers[6][25] ),
    .Y(_09907_),
    .A2(net4552));
 sg13g2_a221oi_1 _15785_ (.B2(_09907_),
    .C1(net4083),
    .B1(_09903_),
    .A1(_05731_),
    .Y(_09908_),
    .A2(net4679));
 sg13g2_a21o_1 _15786_ (.A2(net2970),
    .A1(net4891),
    .B1(_09908_),
    .X(_01062_));
 sg13g2_a22oi_1 _15787_ (.Y(_09909_),
    .B1(net4566),
    .B2(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .A2(net4581),
    .A1(\soc_inst.cpu_core.register_file.registers[5][26] ));
 sg13g2_a22oi_1 _15788_ (.Y(_09910_),
    .B1(net4526),
    .B2(\soc_inst.cpu_core.register_file.registers[8][26] ),
    .A2(net4536),
    .A1(\soc_inst.cpu_core.register_file.registers[10][26] ));
 sg13g2_a22oi_1 _15789_ (.Y(_09911_),
    .B1(net4531),
    .B2(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .A2(net4591),
    .A1(\soc_inst.cpu_core.register_file.registers[13][26] ));
 sg13g2_a22oi_1 _15790_ (.Y(_09912_),
    .B1(net4556),
    .B2(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .A2(net4576),
    .A1(\soc_inst.cpu_core.register_file.registers[9][26] ));
 sg13g2_nand3_1 _15791_ (.B(_09911_),
    .C(_09912_),
    .A(_09910_),
    .Y(_09913_));
 sg13g2_a221oi_1 _15792_ (.B2(\soc_inst.cpu_core.register_file.registers[2][26] ),
    .C1(_09913_),
    .B1(net4546),
    .A1(\soc_inst.cpu_core.register_file.registers[4][26] ),
    .Y(_09914_),
    .A2(net4586));
 sg13g2_a22oi_1 _15793_ (.Y(_09915_),
    .B1(net4551),
    .B2(\soc_inst.cpu_core.register_file.registers[6][26] ),
    .A2(net4571),
    .A1(\soc_inst.cpu_core.register_file.registers[14][26] ));
 sg13g2_a22oi_1 _15794_ (.Y(_09916_),
    .B1(net4541),
    .B2(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .A2(net4561),
    .A1(\soc_inst.cpu_core.register_file.registers[7][26] ));
 sg13g2_nand4_1 _15795_ (.B(_09914_),
    .C(_09915_),
    .A(_09909_),
    .Y(_09917_),
    .D(_09916_));
 sg13g2_a21oi_1 _15796_ (.A1(net719),
    .A2(net4678),
    .Y(_09918_),
    .B1(_09917_));
 sg13g2_nor2_2 _15797_ (.A(net4082),
    .B(_09918_),
    .Y(_09919_));
 sg13g2_a21o_1 _15798_ (.A2(net2932),
    .A1(net4889),
    .B1(_09919_),
    .X(_01063_));
 sg13g2_a22oi_1 _15799_ (.Y(_09920_),
    .B1(net4535),
    .B2(\soc_inst.cpu_core.register_file.registers[10][27] ),
    .A2(net4580),
    .A1(\soc_inst.cpu_core.register_file.registers[5][27] ));
 sg13g2_a22oi_1 _15800_ (.Y(_09921_),
    .B1(net4525),
    .B2(\soc_inst.cpu_core.register_file.registers[8][27] ),
    .A2(net4545),
    .A1(\soc_inst.cpu_core.register_file.registers[2][27] ));
 sg13g2_a22oi_1 _15801_ (.Y(_09922_),
    .B1(net4575),
    .B2(\soc_inst.cpu_core.register_file.registers[9][27] ),
    .A2(net4585),
    .A1(\soc_inst.cpu_core.register_file.registers[4][27] ));
 sg13g2_nand3_1 _15802_ (.B(_09921_),
    .C(_09922_),
    .A(_09920_),
    .Y(_09923_));
 sg13g2_a221oi_1 _15803_ (.B2(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .C1(_09923_),
    .B1(net4540),
    .A1(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .Y(_09924_),
    .A2(net4550));
 sg13g2_a22oi_1 _15804_ (.Y(_09925_),
    .B1(net4530),
    .B2(\soc_inst.cpu_core.register_file.registers[11][27] ),
    .A2(net4565),
    .A1(\soc_inst.cpu_core.register_file.registers[3][27] ));
 sg13g2_a22oi_1 _15805_ (.Y(_09926_),
    .B1(net4570),
    .B2(\soc_inst.cpu_core.register_file.registers[14][27] ),
    .A2(net4590),
    .A1(\soc_inst.cpu_core.register_file.registers[13][27] ));
 sg13g2_a22oi_1 _15806_ (.Y(_09927_),
    .B1(net4555),
    .B2(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .A2(net4560),
    .A1(\soc_inst.cpu_core.register_file.registers[7][27] ));
 sg13g2_nand4_1 _15807_ (.B(_09925_),
    .C(_09926_),
    .A(_09924_),
    .Y(_09928_),
    .D(_09927_));
 sg13g2_a21oi_1 _15808_ (.A1(net1834),
    .A2(net4676),
    .Y(_09929_),
    .B1(_09928_));
 sg13g2_nor2_1 _15809_ (.A(net4083),
    .B(_09929_),
    .Y(_09930_));
 sg13g2_a21o_1 _15810_ (.A2(net942),
    .A1(net4880),
    .B1(_09930_),
    .X(_01064_));
 sg13g2_a22oi_1 _15811_ (.Y(_09931_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][28] ),
    .A2(net4589),
    .A1(\soc_inst.cpu_core.register_file.registers[13][28] ));
 sg13g2_a22oi_1 _15812_ (.Y(_09932_),
    .B1(net4559),
    .B2(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .A2(net4564),
    .A1(\soc_inst.cpu_core.register_file.registers[3][28] ));
 sg13g2_a22oi_1 _15813_ (.Y(_09933_),
    .B1(net4529),
    .B2(\soc_inst.cpu_core.register_file.registers[11][28] ),
    .A2(net4574),
    .A1(\soc_inst.cpu_core.register_file.registers[9][28] ));
 sg13g2_a22oi_1 _15814_ (.Y(_09934_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .A2(net4554),
    .A1(\soc_inst.cpu_core.register_file.registers[12][28] ));
 sg13g2_nand3_1 _15815_ (.B(_09933_),
    .C(_09934_),
    .A(_09932_),
    .Y(_09935_));
 sg13g2_a221oi_1 _15816_ (.B2(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .C1(_09935_),
    .B1(net4569),
    .A1(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .Y(_09936_),
    .A2(net4584));
 sg13g2_a22oi_1 _15817_ (.Y(_09937_),
    .B1(net4534),
    .B2(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][28] ));
 sg13g2_a22oi_1 _15818_ (.Y(_09938_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][28] ),
    .A2(net4549),
    .A1(\soc_inst.cpu_core.register_file.registers[6][28] ));
 sg13g2_nand4_1 _15819_ (.B(_09936_),
    .C(_09937_),
    .A(_09931_),
    .Y(_09939_),
    .D(_09938_));
 sg13g2_a21oi_1 _15820_ (.A1(net654),
    .A2(net4675),
    .Y(_09940_),
    .B1(_09939_));
 sg13g2_nor2_2 _15821_ (.A(net4080),
    .B(_09940_),
    .Y(_09941_));
 sg13g2_a21o_1 _15822_ (.A2(net1030),
    .A1(net4897),
    .B1(_09941_),
    .X(_01065_));
 sg13g2_nand2_1 _15823_ (.Y(_09942_),
    .A(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .B(net4570));
 sg13g2_a21oi_1 _15824_ (.A1(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .A2(net4565),
    .Y(_09943_),
    .B1(net4677));
 sg13g2_a22oi_1 _15825_ (.Y(_09944_),
    .B1(net4535),
    .B2(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .A2(net4590),
    .A1(\soc_inst.cpu_core.register_file.registers[13][29] ));
 sg13g2_a22oi_1 _15826_ (.Y(_09945_),
    .B1(net4540),
    .B2(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .A2(net4550),
    .A1(\soc_inst.cpu_core.register_file.registers[6][29] ));
 sg13g2_nand3_1 _15827_ (.B(_09944_),
    .C(_09945_),
    .A(_09943_),
    .Y(_09946_));
 sg13g2_a221oi_1 _15828_ (.B2(\soc_inst.cpu_core.register_file.registers[8][29] ),
    .C1(_09946_),
    .B1(net4525),
    .A1(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .Y(_09947_),
    .A2(net4585));
 sg13g2_a22oi_1 _15829_ (.Y(_09948_),
    .B1(net4555),
    .B2(\soc_inst.cpu_core.register_file.registers[12][29] ),
    .A2(net4580),
    .A1(\soc_inst.cpu_core.register_file.registers[5][29] ));
 sg13g2_a22oi_1 _15830_ (.Y(_09949_),
    .B1(net4530),
    .B2(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .A2(net4560),
    .A1(\soc_inst.cpu_core.register_file.registers[7][29] ));
 sg13g2_a22oi_1 _15831_ (.Y(_09950_),
    .B1(net4545),
    .B2(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .A2(net4575),
    .A1(\soc_inst.cpu_core.register_file.registers[9][29] ));
 sg13g2_and4_1 _15832_ (.A(_09942_),
    .B(_09948_),
    .C(_09949_),
    .D(_09950_),
    .X(_09951_));
 sg13g2_a221oi_1 _15833_ (.B2(_09951_),
    .C1(net4081),
    .B1(_09947_),
    .A1(_05732_),
    .Y(_09952_),
    .A2(net4676));
 sg13g2_a21o_1 _15834_ (.A2(net2962),
    .A1(net4881),
    .B1(_09952_),
    .X(_01066_));
 sg13g2_a22oi_1 _15835_ (.Y(_09953_),
    .B1(net4542),
    .B2(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .A2(net4592),
    .A1(\soc_inst.cpu_core.register_file.registers[13][30] ));
 sg13g2_a22oi_1 _15836_ (.Y(_09954_),
    .B1(net4568),
    .B2(\soc_inst.cpu_core.register_file.registers[3][30] ),
    .A2(net4587),
    .A1(\soc_inst.cpu_core.register_file.registers[4][30] ));
 sg13g2_a22oi_1 _15837_ (.Y(_09955_),
    .B1(net4548),
    .B2(\soc_inst.cpu_core.register_file.registers[2][30] ),
    .A2(net4552),
    .A1(\soc_inst.cpu_core.register_file.registers[6][30] ));
 sg13g2_a22oi_1 _15838_ (.Y(_09956_),
    .B1(net4557),
    .B2(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .A2(net4562),
    .A1(\soc_inst.cpu_core.register_file.registers[7][30] ));
 sg13g2_nand3_1 _15839_ (.B(_09955_),
    .C(_09956_),
    .A(_09954_),
    .Y(_09957_));
 sg13g2_a221oi_1 _15840_ (.B2(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .C1(_09957_),
    .B1(net4572),
    .A1(\soc_inst.cpu_core.register_file.registers[9][30] ),
    .Y(_09958_),
    .A2(net4578));
 sg13g2_a22oi_1 _15841_ (.Y(_09959_),
    .B1(net4537),
    .B2(\soc_inst.cpu_core.register_file.registers[10][30] ),
    .A2(net4583),
    .A1(\soc_inst.cpu_core.register_file.registers[5][30] ));
 sg13g2_a22oi_1 _15842_ (.Y(_09960_),
    .B1(net4527),
    .B2(\soc_inst.cpu_core.register_file.registers[8][30] ),
    .A2(net4532),
    .A1(\soc_inst.cpu_core.register_file.registers[11][30] ));
 sg13g2_nand4_1 _15843_ (.B(_09958_),
    .C(_09959_),
    .A(_09953_),
    .Y(_09961_),
    .D(_09960_));
 sg13g2_a21oi_1 _15844_ (.A1(net2385),
    .A2(net4678),
    .Y(_09962_),
    .B1(_09961_));
 sg13g2_nor2_2 _15845_ (.A(net4084),
    .B(_09962_),
    .Y(_09963_));
 sg13g2_a21o_1 _15846_ (.A2(net2800),
    .A1(net4892),
    .B1(_09963_),
    .X(_01067_));
 sg13g2_nand2_1 _15847_ (.Y(_09964_),
    .A(\soc_inst.cpu_core.register_file.registers[12][31] ),
    .B(net4554));
 sg13g2_a22oi_1 _15848_ (.Y(_09965_),
    .B1(net4539),
    .B2(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .A2(net4559),
    .A1(\soc_inst.cpu_core.register_file.registers[7][31] ));
 sg13g2_a22oi_1 _15849_ (.Y(_09966_),
    .B1(net4544),
    .B2(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .A2(net4549),
    .A1(\soc_inst.cpu_core.register_file.registers[6][31] ));
 sg13g2_a21oi_1 _15850_ (.A1(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .A2(net4529),
    .Y(_09967_),
    .B1(net4675));
 sg13g2_a22oi_1 _15851_ (.Y(_09968_),
    .B1(net4534),
    .B2(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .A2(net4574),
    .A1(\soc_inst.cpu_core.register_file.registers[9][31] ));
 sg13g2_a22oi_1 _15852_ (.Y(_09969_),
    .B1(net4569),
    .B2(\soc_inst.cpu_core.register_file.registers[14][31] ),
    .A2(net4579),
    .A1(\soc_inst.cpu_core.register_file.registers[5][31] ));
 sg13g2_nand4_1 _15853_ (.B(_09967_),
    .C(_09968_),
    .A(_09966_),
    .Y(_09970_),
    .D(_09969_));
 sg13g2_a22oi_1 _15854_ (.Y(_09971_),
    .B1(net4524),
    .B2(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .A2(net4584),
    .A1(\soc_inst.cpu_core.register_file.registers[4][31] ));
 sg13g2_a22oi_1 _15855_ (.Y(_09972_),
    .B1(net4564),
    .B2(\soc_inst.cpu_core.register_file.registers[3][31] ),
    .A2(net4589),
    .A1(\soc_inst.cpu_core.register_file.registers[13][31] ));
 sg13g2_nand4_1 _15856_ (.B(_09965_),
    .C(_09971_),
    .A(_09964_),
    .Y(_09973_),
    .D(_09972_));
 sg13g2_nor2_2 _15857_ (.A(_09970_),
    .B(_09973_),
    .Y(_09974_));
 sg13g2_nor2_1 _15858_ (.A(net1193),
    .B(_09593_),
    .Y(_09975_));
 sg13g2_nor3_2 _15859_ (.A(net4083),
    .B(_09974_),
    .C(_09975_),
    .Y(_09976_));
 sg13g2_a21o_1 _15860_ (.A2(net2896),
    .A1(net4892),
    .B1(_09976_),
    .X(_01068_));
 sg13g2_mux2_1 _15861_ (.A0(_00273_),
    .A1(net849),
    .S(net4975),
    .X(_01069_));
 sg13g2_mux2_1 _15862_ (.A0(_00274_),
    .A1(net1285),
    .S(net4981),
    .X(_01070_));
 sg13g2_nand2_1 _15863_ (.Y(_09977_),
    .A(net196),
    .B(net4974));
 sg13g2_o21ai_1 _15864_ (.B1(_09977_),
    .Y(_01071_),
    .A1(_05475_),
    .A2(net4974));
 sg13g2_mux2_1 _15865_ (.A0(\soc_inst.cpu_core.ex_instr[3] ),
    .A1(net821),
    .S(net4975),
    .X(_01072_));
 sg13g2_nor2_1 _15866_ (.A(_00275_),
    .B(net4981),
    .Y(_09978_));
 sg13g2_a21oi_1 _15867_ (.A1(_05403_),
    .A2(net4985),
    .Y(_01073_),
    .B1(_09978_));
 sg13g2_nand2_1 _15868_ (.Y(_09979_),
    .A(net586),
    .B(net4984));
 sg13g2_o21ai_1 _15869_ (.B1(_09979_),
    .Y(_01074_),
    .A1(_05476_),
    .A2(net4982));
 sg13g2_mux2_1 _15870_ (.A0(\soc_inst.cpu_core.ex_instr[6] ),
    .A1(net2187),
    .S(net4985),
    .X(_01075_));
 sg13g2_mux2_1 _15871_ (.A0(net2086),
    .A1(net2655),
    .S(net4928),
    .X(_01076_));
 sg13g2_mux2_1 _15872_ (.A0(net2609),
    .A1(net4876),
    .S(net4969),
    .X(_01077_));
 sg13g2_nor2_1 _15873_ (.A(net2252),
    .B(net4969),
    .Y(_09980_));
 sg13g2_a21oi_1 _15874_ (.A1(net4756),
    .A2(net4969),
    .Y(_01078_),
    .B1(_09980_));
 sg13g2_nor2_1 _15875_ (.A(net1870),
    .B(net4965),
    .Y(_09981_));
 sg13g2_a21oi_1 _15876_ (.A1(net4753),
    .A2(net4965),
    .Y(_01079_),
    .B1(_09981_));
 sg13g2_mux2_1 _15877_ (.A0(\soc_inst.cpu_core.ex_instr[15] ),
    .A1(net810),
    .S(net4973),
    .X(_01080_));
 sg13g2_mux2_1 _15878_ (.A0(\soc_inst.cpu_core.ex_instr[16] ),
    .A1(net2130),
    .S(net4955),
    .X(_01081_));
 sg13g2_mux2_1 _15879_ (.A0(\soc_inst.cpu_core.ex_instr[17] ),
    .A1(net1882),
    .S(net4958),
    .X(_01082_));
 sg13g2_mux2_1 _15880_ (.A0(net1529),
    .A1(net2043),
    .S(net4958),
    .X(_01083_));
 sg13g2_mux2_1 _15881_ (.A0(\soc_inst.cpu_core.ex_instr[19] ),
    .A1(net1074),
    .S(net4971),
    .X(_01084_));
 sg13g2_nor2_1 _15882_ (.A(net4968),
    .B(net2041),
    .Y(_09982_));
 sg13g2_a21oi_1 _15883_ (.A1(_05414_),
    .A2(net4987),
    .Y(_01085_),
    .B1(_09982_));
 sg13g2_mux2_1 _15884_ (.A0(net2535),
    .A1(net2563),
    .S(net4987),
    .X(_01086_));
 sg13g2_mux2_1 _15885_ (.A0(\soc_inst.cpu_core.ex_instr[22] ),
    .A1(net1809),
    .S(net4987),
    .X(_01087_));
 sg13g2_nand2_1 _15886_ (.Y(_09983_),
    .A(net855),
    .B(net4967));
 sg13g2_o21ai_1 _15887_ (.B1(_09983_),
    .Y(_01088_),
    .A1(net4958),
    .A2(_05773_));
 sg13g2_mux2_1 _15888_ (.A0(net2362),
    .A1(net2364),
    .S(net4968),
    .X(_01089_));
 sg13g2_nand2_1 _15889_ (.Y(_09984_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .B(net4958));
 sg13g2_o21ai_1 _15890_ (.B1(_09984_),
    .Y(_01090_),
    .A1(net4955),
    .A2(_05775_));
 sg13g2_mux2_1 _15891_ (.A0(net2067),
    .A1(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .S(net4922),
    .X(_01091_));
 sg13g2_mux2_1 _15892_ (.A0(net2078),
    .A1(net2214),
    .S(net4922),
    .X(_01092_));
 sg13g2_mux2_1 _15893_ (.A0(net2082),
    .A1(net2207),
    .S(net4967),
    .X(_01093_));
 sg13g2_nand2_1 _15894_ (.Y(_09985_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .B(net4964));
 sg13g2_o21ai_1 _15895_ (.B1(_09985_),
    .Y(_01094_),
    .A1(net4958),
    .A2(_05778_));
 sg13g2_nand2_1 _15896_ (.Y(_09986_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .B(net4964));
 sg13g2_o21ai_1 _15897_ (.B1(_09986_),
    .Y(_01095_),
    .A1(net4964),
    .A2(_05781_));
 sg13g2_mux2_1 _15898_ (.A0(\soc_inst.cpu_core.ex_funct7[6] ),
    .A1(net2045),
    .S(net4964),
    .X(_01096_));
 sg13g2_nor4_1 _15899_ (.A(net5001),
    .B(net4999),
    .C(net5005),
    .D(net5003),
    .Y(_09987_));
 sg13g2_nand2b_1 _15900_ (.Y(_09988_),
    .B(net4126),
    .A_N(_09987_));
 sg13g2_nor3_1 _15901_ (.A(net5001),
    .B(net4999),
    .C(net5003),
    .Y(_09989_));
 sg13g2_or3_1 _15902_ (.A(net5001),
    .B(net4999),
    .C(net5004),
    .X(_09990_));
 sg13g2_nor2_1 _15903_ (.A(net872),
    .B(net4665),
    .Y(_09991_));
 sg13g2_nand2b_2 _15904_ (.Y(_09992_),
    .B(net5001),
    .A_N(net4999));
 sg13g2_nand2b_1 _15905_ (.Y(_09993_),
    .B(net5005),
    .A_N(net5003));
 sg13g2_nor2_1 _15906_ (.A(_09992_),
    .B(_09993_),
    .Y(_09994_));
 sg13g2_nand2_1 _15907_ (.Y(_09995_),
    .A(net5001),
    .B(net4999));
 sg13g2_nor2_1 _15908_ (.A(_09993_),
    .B(_09995_),
    .Y(_09996_));
 sg13g2_a22oi_1 _15909_ (.Y(_09997_),
    .B1(net4516),
    .B2(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][0] ));
 sg13g2_nand2b_2 _15910_ (.Y(_09998_),
    .B(net4999),
    .A_N(net5001));
 sg13g2_nand2b_2 _15911_ (.Y(_09999_),
    .B(net5003),
    .A_N(net5005));
 sg13g2_nor2_1 _15912_ (.A(_09998_),
    .B(_09999_),
    .Y(_10000_));
 sg13g2_nand2_1 _15913_ (.Y(_10001_),
    .A(net5005),
    .B(net5003));
 sg13g2_nor3_1 _15914_ (.A(net5001),
    .B(net4999),
    .C(_10001_),
    .Y(_10002_));
 sg13g2_nor2_1 _15915_ (.A(_09992_),
    .B(_09999_),
    .Y(_10003_));
 sg13g2_nor2_1 _15916_ (.A(_09998_),
    .B(_10001_),
    .Y(_10004_));
 sg13g2_a22oi_1 _15917_ (.Y(_10005_),
    .B1(net4496),
    .B2(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .A2(net4501),
    .A1(\soc_inst.cpu_core.register_file.registers[6][0] ));
 sg13g2_nor2_1 _15918_ (.A(_09993_),
    .B(_09998_),
    .Y(_10006_));
 sg13g2_nand2_1 _15919_ (.Y(_10007_),
    .A(\soc_inst.cpu_core.register_file.registers[9][0] ),
    .B(net4491));
 sg13g2_nor3_1 _15920_ (.A(net5005),
    .B(net5003),
    .C(_09992_),
    .Y(_10008_));
 sg13g2_nor3_1 _15921_ (.A(net5005),
    .B(net5003),
    .C(_09998_),
    .Y(_10009_));
 sg13g2_nor3_1 _15922_ (.A(net5001),
    .B(net4999),
    .C(_09999_),
    .Y(_10010_));
 sg13g2_nor3_1 _15923_ (.A(net5005),
    .B(net5003),
    .C(_09995_),
    .Y(_10011_));
 sg13g2_nor2_1 _15924_ (.A(_09995_),
    .B(_10001_),
    .Y(_10012_));
 sg13g2_nor2_1 _15925_ (.A(_09995_),
    .B(_09999_),
    .Y(_10013_));
 sg13g2_nor2_1 _15926_ (.A(_09992_),
    .B(_10001_),
    .Y(_10014_));
 sg13g2_a22oi_1 _15927_ (.Y(_10015_),
    .B1(net4471),
    .B2(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .A2(net4481),
    .A1(\soc_inst.cpu_core.register_file.registers[8][0] ));
 sg13g2_a21oi_1 _15928_ (.A1(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .A2(net4461),
    .Y(_10016_),
    .B1(net4673));
 sg13g2_a22oi_1 _15929_ (.Y(_10017_),
    .B1(net4466),
    .B2(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .A2(net4476),
    .A1(\soc_inst.cpu_core.register_file.registers[2][0] ));
 sg13g2_nand4_1 _15930_ (.B(_10015_),
    .C(_10016_),
    .A(_10005_),
    .Y(_10018_),
    .D(_10017_));
 sg13g2_a22oi_1 _15931_ (.Y(_10019_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .A2(net4511),
    .A1(\soc_inst.cpu_core.register_file.registers[10][0] ));
 sg13g2_a22oi_1 _15932_ (.Y(_10020_),
    .B1(net4486),
    .B2(\soc_inst.cpu_core.register_file.registers[4][0] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][0] ));
 sg13g2_nand4_1 _15933_ (.B(_10007_),
    .C(_10019_),
    .A(_09997_),
    .Y(_10021_),
    .D(_10020_));
 sg13g2_nor2_1 _15934_ (.A(_10018_),
    .B(_10021_),
    .Y(_10022_));
 sg13g2_nor3_2 _15935_ (.A(net4078),
    .B(_09991_),
    .C(_10022_),
    .Y(_10023_));
 sg13g2_a21o_1 _15936_ (.A2(net2256),
    .A1(net4932),
    .B1(_10023_),
    .X(_01097_));
 sg13g2_nand2_1 _15937_ (.Y(_10024_),
    .A(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .B(net4466));
 sg13g2_a22oi_1 _15938_ (.Y(_10025_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .A2(net4486),
    .A1(\soc_inst.cpu_core.register_file.registers[4][1] ));
 sg13g2_a21oi_1 _15939_ (.A1(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .A2(net4511),
    .Y(_10026_),
    .B1(net4673));
 sg13g2_a22oi_1 _15940_ (.Y(_10027_),
    .B1(net4461),
    .B2(\soc_inst.cpu_core.register_file.registers[14][1] ),
    .A2(net4496),
    .A1(\soc_inst.cpu_core.register_file.registers[11][1] ));
 sg13g2_a22oi_1 _15941_ (.Y(_10028_),
    .B1(net4471),
    .B2(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .A2(net4501),
    .A1(\soc_inst.cpu_core.register_file.registers[6][1] ));
 sg13g2_nand4_1 _15942_ (.B(_10026_),
    .C(_10027_),
    .A(_10025_),
    .Y(_10029_),
    .D(_10028_));
 sg13g2_a22oi_1 _15943_ (.Y(_10030_),
    .B1(net4491),
    .B2(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][1] ));
 sg13g2_a22oi_1 _15944_ (.Y(_10031_),
    .B1(net4476),
    .B2(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .A2(net4481),
    .A1(\soc_inst.cpu_core.register_file.registers[8][1] ));
 sg13g2_a22oi_1 _15945_ (.Y(_10032_),
    .B1(net4516),
    .B2(\soc_inst.cpu_core.register_file.registers[13][1] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][1] ));
 sg13g2_nand4_1 _15946_ (.B(_10030_),
    .C(_10031_),
    .A(_10024_),
    .Y(_10033_),
    .D(_10032_));
 sg13g2_nor2_1 _15947_ (.A(_10029_),
    .B(_10033_),
    .Y(_10034_));
 sg13g2_nor2_1 _15948_ (.A(net986),
    .B(net4665),
    .Y(_10035_));
 sg13g2_nor3_2 _15949_ (.A(net4077),
    .B(_10034_),
    .C(_10035_),
    .Y(_10036_));
 sg13g2_a21o_1 _15950_ (.A2(net1057),
    .A1(net4890),
    .B1(_10036_),
    .X(_01098_));
 sg13g2_nand2_1 _15951_ (.Y(_10037_),
    .A(\soc_inst.cpu_core.register_file.registers[8][2] ),
    .B(net4481));
 sg13g2_a22oi_1 _15952_ (.Y(_10038_),
    .B1(net4466),
    .B2(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .A2(net4501),
    .A1(\soc_inst.cpu_core.register_file.registers[6][2] ));
 sg13g2_a22oi_1 _15953_ (.Y(_10039_),
    .B1(net4476),
    .B2(\soc_inst.cpu_core.register_file.registers[2][2] ),
    .A2(net4491),
    .A1(\soc_inst.cpu_core.register_file.registers[9][2] ));
 sg13g2_a22oi_1 _15954_ (.Y(_10040_),
    .B1(net4487),
    .B2(\soc_inst.cpu_core.register_file.registers[4][2] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][2] ));
 sg13g2_a22oi_1 _15955_ (.Y(_10041_),
    .B1(net4516),
    .B2(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][2] ));
 sg13g2_a21oi_1 _15956_ (.A1(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .A2(net4456),
    .Y(_10042_),
    .B1(net4673));
 sg13g2_nand4_1 _15957_ (.B(_10040_),
    .C(_10041_),
    .A(_10039_),
    .Y(_10043_),
    .D(_10042_));
 sg13g2_a22oi_1 _15958_ (.Y(_10044_),
    .B1(net4461),
    .B2(\soc_inst.cpu_core.register_file.registers[14][2] ),
    .A2(net4511),
    .A1(\soc_inst.cpu_core.register_file.registers[10][2] ));
 sg13g2_a22oi_1 _15959_ (.Y(_10045_),
    .B1(net4471),
    .B2(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .A2(net4496),
    .A1(\soc_inst.cpu_core.register_file.registers[11][2] ));
 sg13g2_nand4_1 _15960_ (.B(_10038_),
    .C(_10044_),
    .A(_10037_),
    .Y(_10046_),
    .D(_10045_));
 sg13g2_nor2_1 _15961_ (.A(_10043_),
    .B(_10046_),
    .Y(_10047_));
 sg13g2_nor2_1 _15962_ (.A(net673),
    .B(net4665),
    .Y(_10048_));
 sg13g2_nor3_2 _15963_ (.A(net4078),
    .B(_10047_),
    .C(_10048_),
    .Y(_10049_));
 sg13g2_a21o_1 _15964_ (.A2(net1404),
    .A1(net4934),
    .B1(_10049_),
    .X(_01099_));
 sg13g2_nor2_1 _15965_ (.A(net732),
    .B(net4666),
    .Y(_10050_));
 sg13g2_nand2_1 _15966_ (.Y(_10051_),
    .A(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .B(net4501));
 sg13g2_a22oi_1 _15967_ (.Y(_10052_),
    .B1(net4486),
    .B2(\soc_inst.cpu_core.register_file.registers[4][3] ),
    .A2(net4511),
    .A1(\soc_inst.cpu_core.register_file.registers[10][3] ));
 sg13g2_a22oi_1 _15968_ (.Y(_10053_),
    .B1(net4471),
    .B2(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .A2(net4481),
    .A1(\soc_inst.cpu_core.register_file.registers[8][3] ));
 sg13g2_a21oi_1 _15969_ (.A1(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .A2(net4466),
    .Y(_10054_),
    .B1(net4673));
 sg13g2_a22oi_1 _15970_ (.Y(_10055_),
    .B1(net4496),
    .B2(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][3] ));
 sg13g2_a22oi_1 _15971_ (.Y(_10056_),
    .B1(net4491),
    .B2(\soc_inst.cpu_core.register_file.registers[9][3] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][3] ));
 sg13g2_nand4_1 _15972_ (.B(_10054_),
    .C(_10055_),
    .A(_10053_),
    .Y(_10057_),
    .D(_10056_));
 sg13g2_a22oi_1 _15973_ (.Y(_10058_),
    .B1(net4476),
    .B2(\soc_inst.cpu_core.register_file.registers[2][3] ),
    .A2(net4516),
    .A1(\soc_inst.cpu_core.register_file.registers[13][3] ));
 sg13g2_a22oi_1 _15974_ (.Y(_10059_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .A2(net4461),
    .A1(\soc_inst.cpu_core.register_file.registers[14][3] ));
 sg13g2_nand4_1 _15975_ (.B(_10052_),
    .C(_10058_),
    .A(_10051_),
    .Y(_10060_),
    .D(_10059_));
 sg13g2_nor2_2 _15976_ (.A(_10057_),
    .B(_10060_),
    .Y(_10061_));
 sg13g2_nor3_2 _15977_ (.A(net4077),
    .B(_10050_),
    .C(_10061_),
    .Y(_10062_));
 sg13g2_a21o_1 _15978_ (.A2(net875),
    .A1(net4896),
    .B1(_10062_),
    .X(_01100_));
 sg13g2_nand2_1 _15979_ (.Y(_10063_),
    .A(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .B(net4482));
 sg13g2_a22oi_1 _15980_ (.Y(_10064_),
    .B1(net4487),
    .B2(\soc_inst.cpu_core.register_file.registers[4][4] ),
    .A2(net4492),
    .A1(\soc_inst.cpu_core.register_file.registers[9][4] ));
 sg13g2_a22oi_1 _15981_ (.Y(_10065_),
    .B1(net4477),
    .B2(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .A2(net4507),
    .A1(\soc_inst.cpu_core.register_file.registers[3][4] ));
 sg13g2_a21oi_1 _15982_ (.A1(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .A2(net4457),
    .Y(_10066_),
    .B1(net4671));
 sg13g2_nand3_1 _15983_ (.B(_10065_),
    .C(_10066_),
    .A(_10064_),
    .Y(_10067_));
 sg13g2_a221oi_1 _15984_ (.B2(\soc_inst.cpu_core.register_file.registers[14][4] ),
    .C1(_10067_),
    .B1(net4462),
    .A1(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .Y(_10068_),
    .A2(net4521));
 sg13g2_a22oi_1 _15985_ (.Y(_10069_),
    .B1(net4512),
    .B2(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .A2(net4517),
    .A1(\soc_inst.cpu_core.register_file.registers[13][4] ));
 sg13g2_a22oi_1 _15986_ (.Y(_10070_),
    .B1(net4472),
    .B2(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .A2(net4497),
    .A1(\soc_inst.cpu_core.register_file.registers[11][4] ));
 sg13g2_nand3_1 _15987_ (.B(_10069_),
    .C(_10070_),
    .A(_10063_),
    .Y(_10071_));
 sg13g2_a221oi_1 _15988_ (.B2(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .C1(_10071_),
    .B1(net4467),
    .A1(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .Y(_10072_),
    .A2(net4502));
 sg13g2_a221oi_1 _15989_ (.B2(_10072_),
    .C1(net4079),
    .B1(_10068_),
    .A1(_05723_),
    .Y(_10073_),
    .A2(net4672));
 sg13g2_a21o_1 _15990_ (.A2(net2275),
    .A1(net4943),
    .B1(_10073_),
    .X(_01101_));
 sg13g2_a21oi_1 _15991_ (.A1(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .A2(net4502),
    .Y(_10074_),
    .B1(net4672));
 sg13g2_nand2_1 _15992_ (.Y(_10075_),
    .A(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .B(net4521));
 sg13g2_a22oi_1 _15993_ (.Y(_10076_),
    .B1(net4486),
    .B2(\soc_inst.cpu_core.register_file.registers[4][5] ),
    .A2(net4491),
    .A1(\soc_inst.cpu_core.register_file.registers[9][5] ));
 sg13g2_a22oi_1 _15994_ (.Y(_10077_),
    .B1(net4497),
    .B2(\soc_inst.cpu_core.register_file.registers[11][5] ),
    .A2(net4512),
    .A1(\soc_inst.cpu_core.register_file.registers[10][5] ));
 sg13g2_a22oi_1 _15995_ (.Y(_10078_),
    .B1(net4482),
    .B2(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .A2(net4507),
    .A1(\soc_inst.cpu_core.register_file.registers[3][5] ));
 sg13g2_nand4_1 _15996_ (.B(_10076_),
    .C(_10077_),
    .A(_10074_),
    .Y(_10079_),
    .D(_10078_));
 sg13g2_a22oi_1 _15997_ (.Y(_10080_),
    .B1(net4467),
    .B2(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .A2(net4517),
    .A1(\soc_inst.cpu_core.register_file.registers[13][5] ));
 sg13g2_a22oi_1 _15998_ (.Y(_10081_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .A2(net4472),
    .A1(\soc_inst.cpu_core.register_file.registers[12][5] ));
 sg13g2_a22oi_1 _15999_ (.Y(_10082_),
    .B1(net4462),
    .B2(\soc_inst.cpu_core.register_file.registers[14][5] ),
    .A2(net4477),
    .A1(\soc_inst.cpu_core.register_file.registers[2][5] ));
 sg13g2_nand4_1 _16000_ (.B(_10080_),
    .C(_10081_),
    .A(_10075_),
    .Y(_10083_),
    .D(_10082_));
 sg13g2_nor2_2 _16001_ (.A(_10079_),
    .B(_10083_),
    .Y(_10084_));
 sg13g2_nor2_1 _16002_ (.A(net879),
    .B(net4666),
    .Y(_10085_));
 sg13g2_nor3_2 _16003_ (.A(net4078),
    .B(_10084_),
    .C(_10085_),
    .Y(_10086_));
 sg13g2_a21o_1 _16004_ (.A2(net2299),
    .A1(net4943),
    .B1(_10086_),
    .X(_01102_));
 sg13g2_nor2_1 _16005_ (.A(net1267),
    .B(net4666),
    .Y(_10087_));
 sg13g2_nand2_1 _16006_ (.Y(_10088_),
    .A(\soc_inst.cpu_core.register_file.registers[9][6] ),
    .B(net4492));
 sg13g2_a22oi_1 _16007_ (.Y(_10089_),
    .B1(net4517),
    .B2(\soc_inst.cpu_core.register_file.registers[13][6] ),
    .A2(net4521),
    .A1(\soc_inst.cpu_core.register_file.registers[5][6] ));
 sg13g2_a21oi_1 _16008_ (.A1(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .A2(net4507),
    .Y(_10090_),
    .B1(net4671));
 sg13g2_a22oi_1 _16009_ (.Y(_10091_),
    .B1(net4472),
    .B2(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .A2(net4502),
    .A1(\soc_inst.cpu_core.register_file.registers[6][6] ));
 sg13g2_a22oi_1 _16010_ (.Y(_10092_),
    .B1(net4487),
    .B2(\soc_inst.cpu_core.register_file.registers[4][6] ),
    .A2(net4512),
    .A1(\soc_inst.cpu_core.register_file.registers[10][6] ));
 sg13g2_nand4_1 _16011_ (.B(_10090_),
    .C(_10091_),
    .A(_10089_),
    .Y(_10093_),
    .D(_10092_));
 sg13g2_a22oi_1 _16012_ (.Y(_10094_),
    .B1(net4462),
    .B2(\soc_inst.cpu_core.register_file.registers[14][6] ),
    .A2(net4477),
    .A1(\soc_inst.cpu_core.register_file.registers[2][6] ));
 sg13g2_a22oi_1 _16013_ (.Y(_10095_),
    .B1(net4482),
    .B2(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .A2(net4497),
    .A1(\soc_inst.cpu_core.register_file.registers[11][6] ));
 sg13g2_a22oi_1 _16014_ (.Y(_10096_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .A2(net4467),
    .A1(\soc_inst.cpu_core.register_file.registers[15][6] ));
 sg13g2_nand4_1 _16015_ (.B(_10094_),
    .C(_10095_),
    .A(_10088_),
    .Y(_10097_),
    .D(_10096_));
 sg13g2_nor2_2 _16016_ (.A(_10093_),
    .B(_10097_),
    .Y(_10098_));
 sg13g2_nor3_2 _16017_ (.A(net4078),
    .B(_10087_),
    .C(_10098_),
    .Y(_10099_));
 sg13g2_a21o_1 _16018_ (.A2(net1261),
    .A1(net4896),
    .B1(_10099_),
    .X(_01103_));
 sg13g2_nand2_1 _16019_ (.Y(_10100_),
    .A(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .B(net4516));
 sg13g2_a22oi_1 _16020_ (.Y(_10101_),
    .B1(net4486),
    .B2(\soc_inst.cpu_core.register_file.registers[4][7] ),
    .A2(net4491),
    .A1(\soc_inst.cpu_core.register_file.registers[9][7] ));
 sg13g2_a22oi_1 _16021_ (.Y(_10102_),
    .B1(net4461),
    .B2(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][7] ));
 sg13g2_a21oi_1 _16022_ (.A1(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .A2(net4501),
    .Y(_10103_),
    .B1(net4673));
 sg13g2_a22oi_1 _16023_ (.Y(_10104_),
    .B1(net4476),
    .B2(\soc_inst.cpu_core.register_file.registers[2][7] ),
    .A2(net4481),
    .A1(\soc_inst.cpu_core.register_file.registers[8][7] ));
 sg13g2_nand4_1 _16024_ (.B(_10102_),
    .C(_10103_),
    .A(_10101_),
    .Y(_10105_),
    .D(_10104_));
 sg13g2_a22oi_1 _16025_ (.Y(_10106_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .A2(net4511),
    .A1(\soc_inst.cpu_core.register_file.registers[10][7] ));
 sg13g2_a22oi_1 _16026_ (.Y(_10107_),
    .B1(net4466),
    .B2(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .A2(net4471),
    .A1(\soc_inst.cpu_core.register_file.registers[12][7] ));
 sg13g2_a22oi_1 _16027_ (.Y(_10108_),
    .B1(net4496),
    .B2(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][7] ));
 sg13g2_nand4_1 _16028_ (.B(_10106_),
    .C(_10107_),
    .A(_10100_),
    .Y(_10109_),
    .D(_10108_));
 sg13g2_nor2_1 _16029_ (.A(_10105_),
    .B(_10109_),
    .Y(_10110_));
 sg13g2_nor2_1 _16030_ (.A(net2016),
    .B(net4665),
    .Y(_10111_));
 sg13g2_nor3_2 _16031_ (.A(net4077),
    .B(_10110_),
    .C(_10111_),
    .Y(_10112_));
 sg13g2_a21o_1 _16032_ (.A2(net1606),
    .A1(net4896),
    .B1(_10112_),
    .X(_01104_));
 sg13g2_a22oi_1 _16033_ (.Y(_10113_),
    .B1(net4489),
    .B2(\soc_inst.cpu_core.register_file.registers[9][8] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][8] ));
 sg13g2_nand2_1 _16034_ (.Y(_10114_),
    .A(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .B(net4464));
 sg13g2_a22oi_1 _16035_ (.Y(_10115_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .A2(net4479),
    .A1(\soc_inst.cpu_core.register_file.registers[8][8] ));
 sg13g2_a21oi_1 _16036_ (.A1(\soc_inst.cpu_core.register_file.registers[4][8] ),
    .A2(net4484),
    .Y(_10116_),
    .B1(net4670));
 sg13g2_a22oi_1 _16037_ (.Y(_10117_),
    .B1(net4474),
    .B2(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .A2(net4499),
    .A1(\soc_inst.cpu_core.register_file.registers[6][8] ));
 sg13g2_nand4_1 _16038_ (.B(_10115_),
    .C(_10116_),
    .A(_10113_),
    .Y(_10118_),
    .D(_10117_));
 sg13g2_a22oi_1 _16039_ (.Y(_10119_),
    .B1(net4469),
    .B2(\soc_inst.cpu_core.register_file.registers[12][8] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][8] ));
 sg13g2_a22oi_1 _16040_ (.Y(_10120_),
    .B1(net4494),
    .B2(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .A2(net4514),
    .A1(\soc_inst.cpu_core.register_file.registers[13][8] ));
 sg13g2_a22oi_1 _16041_ (.Y(_10121_),
    .B1(net4454),
    .B2(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .A2(net4509),
    .A1(\soc_inst.cpu_core.register_file.registers[10][8] ));
 sg13g2_nand4_1 _16042_ (.B(_10119_),
    .C(_10120_),
    .A(_10114_),
    .Y(_10122_),
    .D(_10121_));
 sg13g2_nor2_1 _16043_ (.A(_10118_),
    .B(_10122_),
    .Y(_10123_));
 sg13g2_nor2_1 _16044_ (.A(net1594),
    .B(net4664),
    .Y(_10124_));
 sg13g2_nor3_2 _16045_ (.A(net4077),
    .B(_10123_),
    .C(_10124_),
    .Y(_10125_));
 sg13g2_a21o_1 _16046_ (.A2(net2377),
    .A1(net4907),
    .B1(_10125_),
    .X(_01105_));
 sg13g2_a22oi_1 _16047_ (.Y(_10126_),
    .B1(net4492),
    .B2(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .A2(net4507),
    .A1(\soc_inst.cpu_core.register_file.registers[3][9] ));
 sg13g2_nand2_1 _16048_ (.Y(_10127_),
    .A(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .B(net4512));
 sg13g2_a22oi_1 _16049_ (.Y(_10128_),
    .B1(net4482),
    .B2(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .A2(net4521),
    .A1(\soc_inst.cpu_core.register_file.registers[5][9] ));
 sg13g2_a21oi_1 _16050_ (.A1(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .A2(net4497),
    .Y(_10129_),
    .B1(net4671));
 sg13g2_a22oi_1 _16051_ (.Y(_10130_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .A2(net4472),
    .A1(\soc_inst.cpu_core.register_file.registers[12][9] ));
 sg13g2_a22oi_1 _16052_ (.Y(_10131_),
    .B1(net4477),
    .B2(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .A2(net4487),
    .A1(\soc_inst.cpu_core.register_file.registers[4][9] ));
 sg13g2_and4_1 _16053_ (.A(_10128_),
    .B(_10129_),
    .C(_10130_),
    .D(_10131_),
    .X(_10132_));
 sg13g2_a22oi_1 _16054_ (.Y(_10133_),
    .B1(net4502),
    .B2(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .A2(net4517),
    .A1(\soc_inst.cpu_core.register_file.registers[13][9] ));
 sg13g2_nand3_1 _16055_ (.B(_10127_),
    .C(_10133_),
    .A(_10126_),
    .Y(_10134_));
 sg13g2_a221oi_1 _16056_ (.B2(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .C1(_10134_),
    .B1(net4462),
    .A1(\soc_inst.cpu_core.register_file.registers[15][9] ),
    .Y(_10135_),
    .A2(net4467));
 sg13g2_a221oi_1 _16057_ (.B2(_10135_),
    .C1(net4079),
    .B1(_10132_),
    .A1(_05724_),
    .Y(_10136_),
    .A2(net4671));
 sg13g2_a21o_1 _16058_ (.A2(net2897),
    .A1(net4895),
    .B1(_10136_),
    .X(_01106_));
 sg13g2_nor2_1 _16059_ (.A(net1171),
    .B(net4665),
    .Y(_10137_));
 sg13g2_nand2_1 _16060_ (.Y(_10138_),
    .A(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .B(net4491));
 sg13g2_a22oi_1 _16061_ (.Y(_10139_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .A2(net4461),
    .A1(\soc_inst.cpu_core.register_file.registers[14][10] ));
 sg13g2_a22oi_1 _16062_ (.Y(_10140_),
    .B1(net4471),
    .B2(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .A2(net4516),
    .A1(\soc_inst.cpu_core.register_file.registers[13][10] ));
 sg13g2_a21oi_1 _16063_ (.A1(\soc_inst.cpu_core.register_file.registers[5][10] ),
    .A2(net4522),
    .Y(_10141_),
    .B1(net4673));
 sg13g2_a22oi_1 _16064_ (.Y(_10142_),
    .B1(net4501),
    .B2(\soc_inst.cpu_core.register_file.registers[6][10] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][10] ));
 sg13g2_a22oi_1 _16065_ (.Y(_10143_),
    .B1(net4486),
    .B2(\soc_inst.cpu_core.register_file.registers[4][10] ),
    .A2(net4511),
    .A1(\soc_inst.cpu_core.register_file.registers[10][10] ));
 sg13g2_nand4_1 _16066_ (.B(_10141_),
    .C(_10142_),
    .A(_10140_),
    .Y(_10144_),
    .D(_10143_));
 sg13g2_a22oi_1 _16067_ (.Y(_10145_),
    .B1(net4466),
    .B2(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .A2(net4476),
    .A1(\soc_inst.cpu_core.register_file.registers[2][10] ));
 sg13g2_a22oi_1 _16068_ (.Y(_10146_),
    .B1(net4481),
    .B2(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .A2(net4496),
    .A1(\soc_inst.cpu_core.register_file.registers[11][10] ));
 sg13g2_nand4_1 _16069_ (.B(_10139_),
    .C(_10145_),
    .A(_10138_),
    .Y(_10147_),
    .D(_10146_));
 sg13g2_nor2_1 _16070_ (.A(_10144_),
    .B(_10147_),
    .Y(_10148_));
 sg13g2_nor3_2 _16071_ (.A(net4077),
    .B(_10137_),
    .C(_10148_),
    .Y(_10149_));
 sg13g2_a21o_1 _16072_ (.A2(net2576),
    .A1(net4893),
    .B1(_10149_),
    .X(_01107_));
 sg13g2_a22oi_1 _16073_ (.Y(_10150_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .A2(net4461),
    .A1(\soc_inst.cpu_core.register_file.registers[14][11] ));
 sg13g2_nand2_1 _16074_ (.Y(_10151_),
    .A(\soc_inst.cpu_core.register_file.registers[4][11] ),
    .B(net4486));
 sg13g2_a22oi_1 _16075_ (.Y(_10152_),
    .B1(net4471),
    .B2(\soc_inst.cpu_core.register_file.registers[12][11] ),
    .A2(net4496),
    .A1(\soc_inst.cpu_core.register_file.registers[11][11] ));
 sg13g2_a22oi_1 _16076_ (.Y(_10153_),
    .B1(net4516),
    .B2(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][11] ));
 sg13g2_a21oi_1 _16077_ (.A1(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .A2(net4511),
    .Y(_10154_),
    .B1(net4673));
 sg13g2_a22oi_1 _16078_ (.Y(_10155_),
    .B1(net4481),
    .B2(\soc_inst.cpu_core.register_file.registers[8][11] ),
    .A2(net4501),
    .A1(\soc_inst.cpu_core.register_file.registers[6][11] ));
 sg13g2_nand4_1 _16079_ (.B(_10153_),
    .C(_10154_),
    .A(_10150_),
    .Y(_10156_),
    .D(_10155_));
 sg13g2_a22oi_1 _16080_ (.Y(_10157_),
    .B1(net4492),
    .B2(\soc_inst.cpu_core.register_file.registers[9][11] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][11] ));
 sg13g2_a22oi_1 _16081_ (.Y(_10158_),
    .B1(net4466),
    .B2(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .A2(net4476),
    .A1(\soc_inst.cpu_core.register_file.registers[2][11] ));
 sg13g2_nand4_1 _16082_ (.B(_10152_),
    .C(_10157_),
    .A(_10151_),
    .Y(_10159_),
    .D(_10158_));
 sg13g2_nor2_2 _16083_ (.A(_10156_),
    .B(_10159_),
    .Y(_10160_));
 sg13g2_nor2_1 _16084_ (.A(net1845),
    .B(net4665),
    .Y(_10161_));
 sg13g2_nor3_2 _16085_ (.A(net4077),
    .B(_10160_),
    .C(_10161_),
    .Y(_10162_));
 sg13g2_a21o_1 _16086_ (.A2(net2846),
    .A1(net4894),
    .B1(_10162_),
    .X(_01108_));
 sg13g2_nand2_1 _16087_ (.Y(_10163_),
    .A(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .B(net4482));
 sg13g2_a22oi_1 _16088_ (.Y(_10164_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .A2(net4467),
    .A1(\soc_inst.cpu_core.register_file.registers[15][12] ));
 sg13g2_a22oi_1 _16089_ (.Y(_10165_),
    .B1(net4487),
    .B2(\soc_inst.cpu_core.register_file.registers[4][12] ),
    .A2(net4492),
    .A1(\soc_inst.cpu_core.register_file.registers[9][12] ));
 sg13g2_a22oi_1 _16090_ (.Y(_10166_),
    .B1(net4477),
    .B2(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .A2(net4507),
    .A1(\soc_inst.cpu_core.register_file.registers[3][12] ));
 sg13g2_a22oi_1 _16091_ (.Y(_10167_),
    .B1(net4462),
    .B2(\soc_inst.cpu_core.register_file.registers[14][12] ),
    .A2(net4523),
    .A1(\soc_inst.cpu_core.register_file.registers[5][12] ));
 sg13g2_a21oi_1 _16092_ (.A1(\soc_inst.cpu_core.register_file.registers[6][12] ),
    .A2(net4502),
    .Y(_10168_),
    .B1(net4672));
 sg13g2_nand4_1 _16093_ (.B(_10166_),
    .C(_10167_),
    .A(_10165_),
    .Y(_10169_),
    .D(_10168_));
 sg13g2_a22oi_1 _16094_ (.Y(_10170_),
    .B1(net4512),
    .B2(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .A2(net4517),
    .A1(\soc_inst.cpu_core.register_file.registers[13][12] ));
 sg13g2_a22oi_1 _16095_ (.Y(_10171_),
    .B1(net4472),
    .B2(\soc_inst.cpu_core.register_file.registers[12][12] ),
    .A2(net4497),
    .A1(\soc_inst.cpu_core.register_file.registers[11][12] ));
 sg13g2_nand4_1 _16096_ (.B(_10164_),
    .C(_10170_),
    .A(_10163_),
    .Y(_10172_),
    .D(_10171_));
 sg13g2_nor2_1 _16097_ (.A(_10169_),
    .B(_10172_),
    .Y(_10173_));
 sg13g2_nor2_1 _16098_ (.A(net1335),
    .B(net4666),
    .Y(_10174_));
 sg13g2_nor3_2 _16099_ (.A(net4079),
    .B(_10173_),
    .C(_10174_),
    .Y(_10175_));
 sg13g2_a21o_1 _16100_ (.A2(net1373),
    .A1(net4893),
    .B1(_10175_),
    .X(_01109_));
 sg13g2_nor2_1 _16101_ (.A(net715),
    .B(net4664),
    .Y(_10176_));
 sg13g2_nand2_1 _16102_ (.Y(_10177_),
    .A(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .B(net4504));
 sg13g2_a22oi_1 _16103_ (.Y(_10178_),
    .B1(net4479),
    .B2(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .A2(net4484),
    .A1(\soc_inst.cpu_core.register_file.registers[4][13] ));
 sg13g2_a22oi_1 _16104_ (.Y(_10179_),
    .B1(net4464),
    .B2(\soc_inst.cpu_core.register_file.registers[15][13] ),
    .A2(net4494),
    .A1(\soc_inst.cpu_core.register_file.registers[11][13] ));
 sg13g2_a21oi_1 _16105_ (.A1(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .A2(net4474),
    .Y(_10180_),
    .B1(net4670));
 sg13g2_a22oi_1 _16106_ (.Y(_10181_),
    .B1(net4489),
    .B2(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .A2(net4499),
    .A1(\soc_inst.cpu_core.register_file.registers[6][13] ));
 sg13g2_nand4_1 _16107_ (.B(_10179_),
    .C(_10180_),
    .A(_10178_),
    .Y(_10182_),
    .D(_10181_));
 sg13g2_a22oi_1 _16108_ (.Y(_10183_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .A2(net4509),
    .A1(\soc_inst.cpu_core.register_file.registers[10][13] ));
 sg13g2_a22oi_1 _16109_ (.Y(_10184_),
    .B1(net4454),
    .B2(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][13] ));
 sg13g2_a22oi_1 _16110_ (.Y(_10185_),
    .B1(net4469),
    .B2(\soc_inst.cpu_core.register_file.registers[12][13] ),
    .A2(net4514),
    .A1(\soc_inst.cpu_core.register_file.registers[13][13] ));
 sg13g2_nand4_1 _16111_ (.B(_10183_),
    .C(_10184_),
    .A(_10177_),
    .Y(_10186_),
    .D(_10185_));
 sg13g2_nor2_1 _16112_ (.A(_10182_),
    .B(_10186_),
    .Y(_10187_));
 sg13g2_nor3_2 _16113_ (.A(net4075),
    .B(_10176_),
    .C(_10187_),
    .Y(_10188_));
 sg13g2_a21o_1 _16114_ (.A2(net2257),
    .A1(net4905),
    .B1(_10188_),
    .X(_01110_));
 sg13g2_nand2_1 _16115_ (.Y(_10189_),
    .A(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .B(net4517));
 sg13g2_a21oi_1 _16116_ (.A1(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .A2(net4482),
    .Y(_10190_),
    .B1(net4671));
 sg13g2_a22oi_1 _16117_ (.Y(_10191_),
    .B1(net4477),
    .B2(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .A2(net4492),
    .A1(\soc_inst.cpu_core.register_file.registers[9][14] ));
 sg13g2_a22oi_1 _16118_ (.Y(_10192_),
    .B1(net4467),
    .B2(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .A2(net4507),
    .A1(\soc_inst.cpu_core.register_file.registers[3][14] ));
 sg13g2_a22oi_1 _16119_ (.Y(_10193_),
    .B1(net4497),
    .B2(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .A2(net4502),
    .A1(\soc_inst.cpu_core.register_file.registers[6][14] ));
 sg13g2_and4_1 _16120_ (.A(_10190_),
    .B(_10191_),
    .C(_10192_),
    .D(_10193_),
    .X(_10194_));
 sg13g2_a22oi_1 _16121_ (.Y(_10195_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .A2(net4472),
    .A1(\soc_inst.cpu_core.register_file.registers[12][14] ));
 sg13g2_a22oi_1 _16122_ (.Y(_10196_),
    .B1(net4462),
    .B2(\soc_inst.cpu_core.register_file.registers[14][14] ),
    .A2(net4512),
    .A1(\soc_inst.cpu_core.register_file.registers[10][14] ));
 sg13g2_nand3_1 _16123_ (.B(_10195_),
    .C(_10196_),
    .A(_10189_),
    .Y(_10197_));
 sg13g2_a221oi_1 _16124_ (.B2(\soc_inst.cpu_core.register_file.registers[4][14] ),
    .C1(_10197_),
    .B1(net4487),
    .A1(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .Y(_10198_),
    .A2(net4521));
 sg13g2_a221oi_1 _16125_ (.B2(_10198_),
    .C1(net4078),
    .B1(_10194_),
    .A1(_05726_),
    .Y(_10199_),
    .A2(net4671));
 sg13g2_a21o_1 _16126_ (.A2(net1334),
    .A1(net4891),
    .B1(_10199_),
    .X(_01111_));
 sg13g2_nand2_1 _16127_ (.Y(_10200_),
    .A(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .B(net4515));
 sg13g2_a21oi_1 _16128_ (.A1(\soc_inst.cpu_core.register_file.registers[9][15] ),
    .A2(net4490),
    .Y(_10201_),
    .B1(net4668));
 sg13g2_a22oi_1 _16129_ (.Y(_10202_),
    .B1(net4460),
    .B2(\soc_inst.cpu_core.register_file.registers[14][15] ),
    .A2(net4500),
    .A1(\soc_inst.cpu_core.register_file.registers[6][15] ));
 sg13g2_a22oi_1 _16130_ (.Y(_10203_),
    .B1(net4485),
    .B2(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][15] ));
 sg13g2_nand3_1 _16131_ (.B(_10202_),
    .C(_10203_),
    .A(_10201_),
    .Y(_10204_));
 sg13g2_a221oi_1 _16132_ (.B2(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .C1(_10204_),
    .B1(net4465),
    .A1(\soc_inst.cpu_core.register_file.registers[2][15] ),
    .Y(_10205_),
    .A2(net4475));
 sg13g2_a22oi_1 _16133_ (.Y(_10206_),
    .B1(net4455),
    .B2(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .A2(net4470),
    .A1(\soc_inst.cpu_core.register_file.registers[12][15] ));
 sg13g2_a22oi_1 _16134_ (.Y(_10207_),
    .B1(net4495),
    .B2(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .A2(net4510),
    .A1(\soc_inst.cpu_core.register_file.registers[10][15] ));
 sg13g2_a22oi_1 _16135_ (.Y(_10208_),
    .B1(net4480),
    .B2(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .A2(net4505),
    .A1(\soc_inst.cpu_core.register_file.registers[3][15] ));
 sg13g2_and4_1 _16136_ (.A(_10200_),
    .B(_10206_),
    .C(_10207_),
    .D(_10208_),
    .X(_10209_));
 sg13g2_a221oi_1 _16137_ (.B2(_10209_),
    .C1(net4076),
    .B1(_10205_),
    .A1(_05727_),
    .Y(_10210_),
    .A2(net4669));
 sg13g2_a21o_1 _16138_ (.A2(net2636),
    .A1(net4881),
    .B1(_10210_),
    .X(_01112_));
 sg13g2_nand2_1 _16139_ (.Y(_10211_),
    .A(\soc_inst.cpu_core.register_file.registers[4][16] ),
    .B(net4484));
 sg13g2_a21oi_1 _16140_ (.A1(\soc_inst.cpu_core.register_file.registers[2][16] ),
    .A2(net4474),
    .Y(_10212_),
    .B1(net4670));
 sg13g2_a22oi_1 _16141_ (.Y(_10213_),
    .B1(net4464),
    .B2(\soc_inst.cpu_core.register_file.registers[15][16] ),
    .A2(net4469),
    .A1(\soc_inst.cpu_core.register_file.registers[12][16] ));
 sg13g2_a22oi_1 _16142_ (.Y(_10214_),
    .B1(net4489),
    .B2(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][16] ));
 sg13g2_a22oi_1 _16143_ (.Y(_02156_),
    .B1(net4454),
    .B2(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][16] ));
 sg13g2_nand4_1 _16144_ (.B(_10213_),
    .C(_10214_),
    .A(_10212_),
    .Y(_02157_),
    .D(_02156_));
 sg13g2_a22oi_1 _16145_ (.Y(_02158_),
    .B1(net4479),
    .B2(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .A2(net4509),
    .A1(\soc_inst.cpu_core.register_file.registers[10][16] ));
 sg13g2_a22oi_1 _16146_ (.Y(_02159_),
    .B1(net4499),
    .B2(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .A2(net4514),
    .A1(\soc_inst.cpu_core.register_file.registers[13][16] ));
 sg13g2_a22oi_1 _16147_ (.Y(_02160_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .A2(net4494),
    .A1(\soc_inst.cpu_core.register_file.registers[11][16] ));
 sg13g2_nand4_1 _16148_ (.B(_02158_),
    .C(_02159_),
    .A(_10211_),
    .Y(_02161_),
    .D(_02160_));
 sg13g2_nor2_1 _16149_ (.A(_02157_),
    .B(_02161_),
    .Y(_02162_));
 sg13g2_nor2_1 _16150_ (.A(net1027),
    .B(net4664),
    .Y(_02163_));
 sg13g2_nor3_2 _16151_ (.A(net4075),
    .B(_02162_),
    .C(_02163_),
    .Y(_02164_));
 sg13g2_a21o_1 _16152_ (.A2(net1283),
    .A1(net4899),
    .B1(_02164_),
    .X(_01113_));
 sg13g2_nand2_1 _16153_ (.Y(_02165_),
    .A(\soc_inst.cpu_core.register_file.registers[9][17] ),
    .B(net4490));
 sg13g2_a22oi_1 _16154_ (.Y(_02166_),
    .B1(net4495),
    .B2(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][17] ));
 sg13g2_a22oi_1 _16155_ (.Y(_02167_),
    .B1(net4470),
    .B2(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .A2(net4515),
    .A1(\soc_inst.cpu_core.register_file.registers[13][17] ));
 sg13g2_a21oi_1 _16156_ (.A1(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .A2(net4460),
    .Y(_02168_),
    .B1(net4668));
 sg13g2_a22oi_1 _16157_ (.Y(_02169_),
    .B1(net4465),
    .B2(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .A2(net4485),
    .A1(\soc_inst.cpu_core.register_file.registers[4][17] ));
 sg13g2_nand3_1 _16158_ (.B(_02168_),
    .C(_02169_),
    .A(_02167_),
    .Y(_02170_));
 sg13g2_a221oi_1 _16159_ (.B2(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .C1(_02170_),
    .B1(net4505),
    .A1(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .Y(_02171_),
    .A2(net4510));
 sg13g2_a22oi_1 _16160_ (.Y(_02172_),
    .B1(net4475),
    .B2(\soc_inst.cpu_core.register_file.registers[2][17] ),
    .A2(net4480),
    .A1(\soc_inst.cpu_core.register_file.registers[8][17] ));
 sg13g2_nand3_1 _16161_ (.B(_02166_),
    .C(_02172_),
    .A(_02165_),
    .Y(_02173_));
 sg13g2_a221oi_1 _16162_ (.B2(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .C1(_02173_),
    .B1(net4455),
    .A1(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .Y(_02174_),
    .A2(net4500));
 sg13g2_a221oi_1 _16163_ (.B2(_02174_),
    .C1(net4075),
    .B1(_02171_),
    .A1(_05728_),
    .Y(_02175_),
    .A2(net4668));
 sg13g2_a21o_1 _16164_ (.A2(net2444),
    .A1(net4897),
    .B1(_02175_),
    .X(_01114_));
 sg13g2_a22oi_1 _16165_ (.Y(_02176_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][18] ),
    .A2(net4509),
    .A1(\soc_inst.cpu_core.register_file.registers[10][18] ));
 sg13g2_nand2_1 _16166_ (.Y(_02177_),
    .A(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .B(net4479));
 sg13g2_a21oi_1 _16167_ (.A1(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .A2(net4454),
    .Y(_02178_),
    .B1(net4670));
 sg13g2_a22oi_1 _16168_ (.Y(_02179_),
    .B1(net4464),
    .B2(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .A2(net4499),
    .A1(\soc_inst.cpu_core.register_file.registers[6][18] ));
 sg13g2_a22oi_1 _16169_ (.Y(_02180_),
    .B1(net4474),
    .B2(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .A2(net4489),
    .A1(\soc_inst.cpu_core.register_file.registers[9][18] ));
 sg13g2_a22oi_1 _16170_ (.Y(_02181_),
    .B1(net4484),
    .B2(\soc_inst.cpu_core.register_file.registers[4][18] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][18] ));
 sg13g2_a22oi_1 _16171_ (.Y(_02182_),
    .B1(net4514),
    .B2(\soc_inst.cpu_core.register_file.registers[13][18] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][18] ));
 sg13g2_nand4_1 _16172_ (.B(_02180_),
    .C(_02181_),
    .A(_02178_),
    .Y(_02183_),
    .D(_02182_));
 sg13g2_a22oi_1 _16173_ (.Y(_02184_),
    .B1(net4469),
    .B2(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .A2(net4494),
    .A1(\soc_inst.cpu_core.register_file.registers[11][18] ));
 sg13g2_nand4_1 _16174_ (.B(_02177_),
    .C(_02179_),
    .A(_02176_),
    .Y(_02185_),
    .D(_02184_));
 sg13g2_nor2_1 _16175_ (.A(_02183_),
    .B(_02185_),
    .Y(_02186_));
 sg13g2_nor2_1 _16176_ (.A(net723),
    .B(net4664),
    .Y(_02187_));
 sg13g2_nor3_2 _16177_ (.A(net4075),
    .B(_02186_),
    .C(_02187_),
    .Y(_02188_));
 sg13g2_a21o_1 _16178_ (.A2(net2921),
    .A1(net4899),
    .B1(_02188_),
    .X(_01115_));
 sg13g2_a22oi_1 _16179_ (.Y(_02189_),
    .B1(net4490),
    .B2(\soc_inst.cpu_core.register_file.registers[9][19] ),
    .A2(net4515),
    .A1(\soc_inst.cpu_core.register_file.registers[13][19] ));
 sg13g2_nand2_1 _16180_ (.Y(_02190_),
    .A(\soc_inst.cpu_core.register_file.registers[14][19] ),
    .B(net4460));
 sg13g2_a22oi_1 _16181_ (.Y(_02191_),
    .B1(net4470),
    .B2(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .A2(net4505),
    .A1(\soc_inst.cpu_core.register_file.registers[3][19] ));
 sg13g2_a21oi_1 _16182_ (.A1(\soc_inst.cpu_core.register_file.registers[6][19] ),
    .A2(net4500),
    .Y(_02192_),
    .B1(net4668));
 sg13g2_a22oi_1 _16183_ (.Y(_02193_),
    .B1(net4465),
    .B2(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .A2(net4475),
    .A1(\soc_inst.cpu_core.register_file.registers[2][19] ));
 sg13g2_a22oi_1 _16184_ (.Y(_02194_),
    .B1(net4485),
    .B2(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .A2(net4495),
    .A1(\soc_inst.cpu_core.register_file.registers[11][19] ));
 sg13g2_nand4_1 _16185_ (.B(_02192_),
    .C(_02193_),
    .A(_02189_),
    .Y(_02195_),
    .D(_02194_));
 sg13g2_a22oi_1 _16186_ (.Y(_02196_),
    .B1(net4510),
    .B2(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][19] ));
 sg13g2_a22oi_1 _16187_ (.Y(_02197_),
    .B1(net4455),
    .B2(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .A2(net4480),
    .A1(\soc_inst.cpu_core.register_file.registers[8][19] ));
 sg13g2_nand4_1 _16188_ (.B(_02191_),
    .C(_02196_),
    .A(_02190_),
    .Y(_02198_),
    .D(_02197_));
 sg13g2_nor2_1 _16189_ (.A(_02195_),
    .B(_02198_),
    .Y(_02199_));
 sg13g2_nor2_1 _16190_ (.A(net768),
    .B(net4664),
    .Y(_02200_));
 sg13g2_nor3_2 _16191_ (.A(net4076),
    .B(_02199_),
    .C(_02200_),
    .Y(_02201_));
 sg13g2_a21o_1 _16192_ (.A2(net2836),
    .A1(net4897),
    .B1(_02201_),
    .X(_01116_));
 sg13g2_nand2_1 _16193_ (.Y(_02202_),
    .A(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .B(net4479));
 sg13g2_a22oi_1 _16194_ (.Y(_02203_),
    .B1(net4464),
    .B2(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .A2(net4499),
    .A1(\soc_inst.cpu_core.register_file.registers[6][20] ));
 sg13g2_a22oi_1 _16195_ (.Y(_02204_),
    .B1(net4484),
    .B2(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .A2(net4489),
    .A1(\soc_inst.cpu_core.register_file.registers[9][20] ));
 sg13g2_a22oi_1 _16196_ (.Y(_02205_),
    .B1(net4474),
    .B2(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][20] ));
 sg13g2_a22oi_1 _16197_ (.Y(_02206_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][20] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][20] ));
 sg13g2_a21oi_1 _16198_ (.A1(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .A2(net4454),
    .Y(_02207_),
    .B1(net4670));
 sg13g2_nand4_1 _16199_ (.B(_02205_),
    .C(_02206_),
    .A(_02204_),
    .Y(_02208_),
    .D(_02207_));
 sg13g2_a22oi_1 _16200_ (.Y(_02209_),
    .B1(net4509),
    .B2(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .A2(net4514),
    .A1(\soc_inst.cpu_core.register_file.registers[13][20] ));
 sg13g2_a22oi_1 _16201_ (.Y(_02210_),
    .B1(net4469),
    .B2(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .A2(net4494),
    .A1(\soc_inst.cpu_core.register_file.registers[11][20] ));
 sg13g2_nand4_1 _16202_ (.B(_02203_),
    .C(_02209_),
    .A(_02202_),
    .Y(_02211_),
    .D(_02210_));
 sg13g2_nor2_1 _16203_ (.A(_02208_),
    .B(_02211_),
    .Y(_02212_));
 sg13g2_nor2_1 _16204_ (.A(net1278),
    .B(net4664),
    .Y(_02213_));
 sg13g2_nor3_2 _16205_ (.A(net4075),
    .B(_02212_),
    .C(_02213_),
    .Y(_02214_));
 sg13g2_a21o_1 _16206_ (.A2(net1648),
    .A1(net4900),
    .B1(_02214_),
    .X(_01117_));
 sg13g2_nand2_1 _16207_ (.Y(_02215_),
    .A(\soc_inst.cpu_core.register_file.registers[4][21] ),
    .B(net4485));
 sg13g2_a21oi_1 _16208_ (.A1(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .A2(net4505),
    .Y(_02216_),
    .B1(net4668));
 sg13g2_a22oi_1 _16209_ (.Y(_02217_),
    .B1(net4455),
    .B2(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .A2(net4475),
    .A1(\soc_inst.cpu_core.register_file.registers[2][21] ));
 sg13g2_a22oi_1 _16210_ (.Y(_02218_),
    .B1(net4490),
    .B2(\soc_inst.cpu_core.register_file.registers[9][21] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][21] ));
 sg13g2_nand3_1 _16211_ (.B(_02217_),
    .C(_02218_),
    .A(_02216_),
    .Y(_02219_));
 sg13g2_a221oi_1 _16212_ (.B2(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .C1(_02219_),
    .B1(net4460),
    .A1(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .Y(_02220_),
    .A2(net4510));
 sg13g2_a22oi_1 _16213_ (.Y(_02221_),
    .B1(net4500),
    .B2(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .A2(net4515),
    .A1(\soc_inst.cpu_core.register_file.registers[13][21] ));
 sg13g2_a22oi_1 _16214_ (.Y(_02222_),
    .B1(net4465),
    .B2(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .A2(net4470),
    .A1(\soc_inst.cpu_core.register_file.registers[12][21] ));
 sg13g2_a22oi_1 _16215_ (.Y(_02223_),
    .B1(net4480),
    .B2(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .A2(net4495),
    .A1(\soc_inst.cpu_core.register_file.registers[11][21] ));
 sg13g2_and4_1 _16216_ (.A(_02215_),
    .B(_02221_),
    .C(_02222_),
    .D(_02223_),
    .X(_02224_));
 sg13g2_a221oi_1 _16217_ (.B2(_02224_),
    .C1(net4075),
    .B1(_02220_),
    .A1(_05729_),
    .Y(_02225_),
    .A2(net4668));
 sg13g2_a21o_1 _16218_ (.A2(net1282),
    .A1(net4900),
    .B1(_02225_),
    .X(_01118_));
 sg13g2_a22oi_1 _16219_ (.Y(_02226_),
    .B1(net4475),
    .B2(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .A2(net4480),
    .A1(\soc_inst.cpu_core.register_file.registers[8][22] ));
 sg13g2_nand2_1 _16220_ (.Y(_02227_),
    .A(\soc_inst.cpu_core.register_file.registers[3][22] ),
    .B(net4505));
 sg13g2_a22oi_1 _16221_ (.Y(_02228_),
    .B1(net4485),
    .B2(\soc_inst.cpu_core.register_file.registers[4][22] ),
    .A2(net4490),
    .A1(\soc_inst.cpu_core.register_file.registers[9][22] ));
 sg13g2_a21oi_1 _16222_ (.A1(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .A2(net4500),
    .Y(_02229_),
    .B1(net4668));
 sg13g2_a22oi_1 _16223_ (.Y(_02230_),
    .B1(net4460),
    .B2(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][22] ));
 sg13g2_nand4_1 _16224_ (.B(_02228_),
    .C(_02229_),
    .A(_02226_),
    .Y(_02231_),
    .D(_02230_));
 sg13g2_a22oi_1 _16225_ (.Y(_02232_),
    .B1(net4455),
    .B2(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .A2(net4465),
    .A1(\soc_inst.cpu_core.register_file.registers[15][22] ));
 sg13g2_a22oi_1 _16226_ (.Y(_02233_),
    .B1(net4510),
    .B2(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .A2(net4515),
    .A1(\soc_inst.cpu_core.register_file.registers[13][22] ));
 sg13g2_a22oi_1 _16227_ (.Y(_02234_),
    .B1(net4470),
    .B2(\soc_inst.cpu_core.register_file.registers[12][22] ),
    .A2(net4495),
    .A1(\soc_inst.cpu_core.register_file.registers[11][22] ));
 sg13g2_nand4_1 _16228_ (.B(_02232_),
    .C(_02233_),
    .A(_02227_),
    .Y(_02235_),
    .D(_02234_));
 sg13g2_nor2_1 _16229_ (.A(_02231_),
    .B(_02235_),
    .Y(_02236_));
 sg13g2_nor2_1 _16230_ (.A(net769),
    .B(net4667),
    .Y(_02237_));
 sg13g2_nor3_2 _16231_ (.A(net4076),
    .B(_02236_),
    .C(_02237_),
    .Y(_02238_));
 sg13g2_a21o_1 _16232_ (.A2(net2235),
    .A1(net4897),
    .B1(_02238_),
    .X(_01119_));
 sg13g2_nand2_1 _16233_ (.Y(_02239_),
    .A(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .B(net4519));
 sg13g2_a21oi_1 _16234_ (.A1(\soc_inst.cpu_core.register_file.registers[13][23] ),
    .A2(net4514),
    .Y(_02240_),
    .B1(net4670));
 sg13g2_a22oi_1 _16235_ (.Y(_02241_),
    .B1(net4454),
    .B2(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .A2(net4474),
    .A1(\soc_inst.cpu_core.register_file.registers[2][23] ));
 sg13g2_a22oi_1 _16236_ (.Y(_02242_),
    .B1(net4464),
    .B2(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .A2(net4494),
    .A1(\soc_inst.cpu_core.register_file.registers[11][23] ));
 sg13g2_a22oi_1 _16237_ (.Y(_02243_),
    .B1(net4469),
    .B2(\soc_inst.cpu_core.register_file.registers[12][23] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][23] ));
 sg13g2_nand4_1 _16238_ (.B(_02241_),
    .C(_02242_),
    .A(_02240_),
    .Y(_02244_),
    .D(_02243_));
 sg13g2_a22oi_1 _16239_ (.Y(_02245_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][23] ),
    .A2(net4499),
    .A1(\soc_inst.cpu_core.register_file.registers[6][23] ));
 sg13g2_a22oi_1 _16240_ (.Y(_02246_),
    .B1(net4489),
    .B2(\soc_inst.cpu_core.register_file.registers[9][23] ),
    .A2(net4509),
    .A1(\soc_inst.cpu_core.register_file.registers[10][23] ));
 sg13g2_a22oi_1 _16241_ (.Y(_02247_),
    .B1(net4479),
    .B2(\soc_inst.cpu_core.register_file.registers[8][23] ),
    .A2(net4484),
    .A1(\soc_inst.cpu_core.register_file.registers[4][23] ));
 sg13g2_nand4_1 _16242_ (.B(_02245_),
    .C(_02246_),
    .A(_02239_),
    .Y(_02248_),
    .D(_02247_));
 sg13g2_nor2_1 _16243_ (.A(_02244_),
    .B(_02248_),
    .Y(_02249_));
 sg13g2_nor2_1 _16244_ (.A(net739),
    .B(net4664),
    .Y(_02250_));
 sg13g2_nor3_2 _16245_ (.A(net4075),
    .B(_02249_),
    .C(_02250_),
    .Y(_02251_));
 sg13g2_a21o_1 _16246_ (.A2(net2435),
    .A1(net4899),
    .B1(_02251_),
    .X(_01120_));
 sg13g2_a22oi_1 _16247_ (.Y(_02252_),
    .B1(net4485),
    .B2(\soc_inst.cpu_core.register_file.registers[4][24] ),
    .A2(net4505),
    .A1(\soc_inst.cpu_core.register_file.registers[3][24] ));
 sg13g2_nand2_1 _16248_ (.Y(_02253_),
    .A(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .B(net4495));
 sg13g2_a21oi_1 _16249_ (.A1(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .A2(net4500),
    .Y(_02254_),
    .B1(net4669));
 sg13g2_a22oi_1 _16250_ (.Y(_02255_),
    .B1(net4455),
    .B2(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .A2(net4470),
    .A1(\soc_inst.cpu_core.register_file.registers[12][24] ));
 sg13g2_a22oi_1 _16251_ (.Y(_02256_),
    .B1(net4465),
    .B2(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .A2(net4521),
    .A1(\soc_inst.cpu_core.register_file.registers[5][24] ));
 sg13g2_nand3_1 _16252_ (.B(_02255_),
    .C(_02256_),
    .A(_02254_),
    .Y(_02257_));
 sg13g2_a221oi_1 _16253_ (.B2(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .C1(_02257_),
    .B1(net4480),
    .A1(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .Y(_02258_),
    .A2(net4515));
 sg13g2_a22oi_1 _16254_ (.Y(_02259_),
    .B1(net4475),
    .B2(\soc_inst.cpu_core.register_file.registers[2][24] ),
    .A2(net4490),
    .A1(\soc_inst.cpu_core.register_file.registers[9][24] ));
 sg13g2_nand3_1 _16255_ (.B(_02253_),
    .C(_02259_),
    .A(_02252_),
    .Y(_02260_));
 sg13g2_a221oi_1 _16256_ (.B2(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .C1(_02260_),
    .B1(net4460),
    .A1(\soc_inst.cpu_core.register_file.registers[10][24] ),
    .Y(_02261_),
    .A2(net4510));
 sg13g2_a221oi_1 _16257_ (.B2(_02261_),
    .C1(net4078),
    .B1(_02258_),
    .A1(_05730_),
    .Y(_02262_),
    .A2(net4669));
 sg13g2_a21o_1 _16258_ (.A2(net2501),
    .A1(net4902),
    .B1(_02262_),
    .X(_01121_));
 sg13g2_nand2_1 _16259_ (.Y(_02263_),
    .A(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .B(net4482));
 sg13g2_a22oi_1 _16260_ (.Y(_02264_),
    .B1(net4487),
    .B2(\soc_inst.cpu_core.register_file.registers[4][25] ),
    .A2(net4497),
    .A1(\soc_inst.cpu_core.register_file.registers[11][25] ));
 sg13g2_a22oi_1 _16261_ (.Y(_02265_),
    .B1(net4507),
    .B2(\soc_inst.cpu_core.register_file.registers[3][25] ),
    .A2(net4512),
    .A1(\soc_inst.cpu_core.register_file.registers[10][25] ));
 sg13g2_a21oi_1 _16262_ (.A1(\soc_inst.cpu_core.register_file.registers[5][25] ),
    .A2(net4521),
    .Y(_02266_),
    .B1(net4671));
 sg13g2_nand3_1 _16263_ (.B(_02265_),
    .C(_02266_),
    .A(_02264_),
    .Y(_02267_));
 sg13g2_a221oi_1 _16264_ (.B2(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .C1(_02267_),
    .B1(net4472),
    .A1(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .Y(_02268_),
    .A2(net4492));
 sg13g2_a22oi_1 _16265_ (.Y(_02269_),
    .B1(net4467),
    .B2(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .A2(net4517),
    .A1(\soc_inst.cpu_core.register_file.registers[13][25] ));
 sg13g2_a22oi_1 _16266_ (.Y(_02270_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .A2(net4502),
    .A1(\soc_inst.cpu_core.register_file.registers[6][25] ));
 sg13g2_nand3_1 _16267_ (.B(_02269_),
    .C(_02270_),
    .A(_02263_),
    .Y(_02271_));
 sg13g2_a221oi_1 _16268_ (.B2(\soc_inst.cpu_core.register_file.registers[14][25] ),
    .C1(_02271_),
    .B1(net4462),
    .A1(\soc_inst.cpu_core.register_file.registers[2][25] ),
    .Y(_02272_),
    .A2(net4477));
 sg13g2_a221oi_1 _16269_ (.B2(_02272_),
    .C1(net4078),
    .B1(_02268_),
    .A1(_05731_),
    .Y(_02273_),
    .A2(net4671));
 sg13g2_a21o_1 _16270_ (.A2(net1248),
    .A1(net4887),
    .B1(_02273_),
    .X(_01122_));
 sg13g2_nor2_1 _16271_ (.A(net719),
    .B(net4665),
    .Y(_02274_));
 sg13g2_nand2_1 _16272_ (.Y(_02275_),
    .A(\soc_inst.cpu_core.register_file.registers[10][26] ),
    .B(net4511));
 sg13g2_a21oi_1 _16273_ (.A1(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .A2(net4471),
    .Y(_02276_),
    .B1(net4673));
 sg13g2_a22oi_1 _16274_ (.Y(_02277_),
    .B1(net4456),
    .B2(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .A2(net4491),
    .A1(\soc_inst.cpu_core.register_file.registers[9][26] ));
 sg13g2_a22oi_1 _16275_ (.Y(_02278_),
    .B1(net4496),
    .B2(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .A2(net4516),
    .A1(\soc_inst.cpu_core.register_file.registers[13][26] ));
 sg13g2_a22oi_1 _16276_ (.Y(_02279_),
    .B1(net4476),
    .B2(\soc_inst.cpu_core.register_file.registers[2][26] ),
    .A2(net4506),
    .A1(\soc_inst.cpu_core.register_file.registers[3][26] ));
 sg13g2_nand4_1 _16277_ (.B(_02277_),
    .C(_02278_),
    .A(_02276_),
    .Y(_02280_),
    .D(_02279_));
 sg13g2_a22oi_1 _16278_ (.Y(_02281_),
    .B1(net4466),
    .B2(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .A2(net4522),
    .A1(\soc_inst.cpu_core.register_file.registers[5][26] ));
 sg13g2_a22oi_1 _16279_ (.Y(_02282_),
    .B1(net4461),
    .B2(\soc_inst.cpu_core.register_file.registers[14][26] ),
    .A2(net4481),
    .A1(\soc_inst.cpu_core.register_file.registers[8][26] ));
 sg13g2_a22oi_1 _16280_ (.Y(_02283_),
    .B1(net4486),
    .B2(\soc_inst.cpu_core.register_file.registers[4][26] ),
    .A2(net4501),
    .A1(\soc_inst.cpu_core.register_file.registers[6][26] ));
 sg13g2_nand4_1 _16281_ (.B(_02281_),
    .C(_02282_),
    .A(_02275_),
    .Y(_02284_),
    .D(_02283_));
 sg13g2_nor2_1 _16282_ (.A(_02280_),
    .B(_02284_),
    .Y(_02285_));
 sg13g2_nor3_2 _16283_ (.A(net4077),
    .B(_02274_),
    .C(_02285_),
    .Y(_02286_));
 sg13g2_a21o_1 _16284_ (.A2(net2787),
    .A1(net4903),
    .B1(_02286_),
    .X(_01123_));
 sg13g2_a22oi_1 _16285_ (.Y(_02287_),
    .B1(net4510),
    .B2(\soc_inst.cpu_core.register_file.registers[10][27] ),
    .A2(net4515),
    .A1(\soc_inst.cpu_core.register_file.registers[13][27] ));
 sg13g2_nand2_1 _16286_ (.Y(_02288_),
    .A(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .B(net4455));
 sg13g2_a22oi_1 _16287_ (.Y(_02289_),
    .B1(net4485),
    .B2(\soc_inst.cpu_core.register_file.registers[4][27] ),
    .A2(net4505),
    .A1(\soc_inst.cpu_core.register_file.registers[3][27] ));
 sg13g2_a22oi_1 _16288_ (.Y(_02290_),
    .B1(net4475),
    .B2(\soc_inst.cpu_core.register_file.registers[2][27] ),
    .A2(net4490),
    .A1(\soc_inst.cpu_core.register_file.registers[9][27] ));
 sg13g2_a22oi_1 _16289_ (.Y(_02291_),
    .B1(net4460),
    .B2(\soc_inst.cpu_core.register_file.registers[14][27] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][27] ));
 sg13g2_a21oi_1 _16290_ (.A1(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .A2(net4500),
    .Y(_02292_),
    .B1(net4669));
 sg13g2_nand4_1 _16291_ (.B(_02290_),
    .C(_02291_),
    .A(_02289_),
    .Y(_02293_),
    .D(_02292_));
 sg13g2_a22oi_1 _16292_ (.Y(_02294_),
    .B1(net4465),
    .B2(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .A2(net4470),
    .A1(\soc_inst.cpu_core.register_file.registers[12][27] ));
 sg13g2_a22oi_1 _16293_ (.Y(_02295_),
    .B1(net4480),
    .B2(\soc_inst.cpu_core.register_file.registers[8][27] ),
    .A2(net4495),
    .A1(\soc_inst.cpu_core.register_file.registers[11][27] ));
 sg13g2_nand4_1 _16294_ (.B(_02288_),
    .C(_02294_),
    .A(_02287_),
    .Y(_02296_),
    .D(_02295_));
 sg13g2_nor2_1 _16295_ (.A(_02293_),
    .B(_02296_),
    .Y(_02297_));
 sg13g2_nor2_1 _16296_ (.A(net1834),
    .B(net4667),
    .Y(_02298_));
 sg13g2_nor3_2 _16297_ (.A(net4076),
    .B(_02297_),
    .C(_02298_),
    .Y(_02299_));
 sg13g2_a21o_1 _16298_ (.A2(net2612),
    .A1(net4904),
    .B1(_02299_),
    .X(_01124_));
 sg13g2_nand2_1 _16299_ (.Y(_02300_),
    .A(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .B(net4479));
 sg13g2_a22oi_1 _16300_ (.Y(_02301_),
    .B1(net4484),
    .B2(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .A2(net4489),
    .A1(\soc_inst.cpu_core.register_file.registers[9][28] ));
 sg13g2_a22oi_1 _16301_ (.Y(_02302_),
    .B1(net4474),
    .B2(\soc_inst.cpu_core.register_file.registers[2][28] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][28] ));
 sg13g2_a22oi_1 _16302_ (.Y(_02303_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][28] ));
 sg13g2_a21oi_1 _16303_ (.A1(\soc_inst.cpu_core.register_file.registers[6][28] ),
    .A2(net4499),
    .Y(_02304_),
    .B1(net4670));
 sg13g2_nand4_1 _16304_ (.B(_02302_),
    .C(_02303_),
    .A(_02301_),
    .Y(_02305_),
    .D(_02304_));
 sg13g2_a22oi_1 _16305_ (.Y(_02306_),
    .B1(net4509),
    .B2(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .A2(net4514),
    .A1(\soc_inst.cpu_core.register_file.registers[13][28] ));
 sg13g2_a22oi_1 _16306_ (.Y(_02307_),
    .B1(net4454),
    .B2(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .A2(net4464),
    .A1(\soc_inst.cpu_core.register_file.registers[15][28] ));
 sg13g2_a22oi_1 _16307_ (.Y(_02308_),
    .B1(net4469),
    .B2(\soc_inst.cpu_core.register_file.registers[12][28] ),
    .A2(net4494),
    .A1(\soc_inst.cpu_core.register_file.registers[11][28] ));
 sg13g2_nand4_1 _16308_ (.B(_02306_),
    .C(_02307_),
    .A(_02300_),
    .Y(_02309_),
    .D(_02308_));
 sg13g2_nor2_1 _16309_ (.A(_02305_),
    .B(_02309_),
    .Y(_02310_));
 sg13g2_nor2_1 _16310_ (.A(net654),
    .B(net4664),
    .Y(_02311_));
 sg13g2_nor3_2 _16311_ (.A(net4075),
    .B(_02310_),
    .C(_02311_),
    .Y(_02312_));
 sg13g2_a21o_1 _16312_ (.A2(net2555),
    .A1(net4884),
    .B1(_02312_),
    .X(_01125_));
 sg13g2_nand2_1 _16313_ (.Y(_02313_),
    .A(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .B(net4505));
 sg13g2_a22oi_1 _16314_ (.Y(_02314_),
    .B1(net4485),
    .B2(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .A2(net4500),
    .A1(\soc_inst.cpu_core.register_file.registers[6][29] ));
 sg13g2_a21oi_1 _16315_ (.A1(\soc_inst.cpu_core.register_file.registers[9][29] ),
    .A2(net4490),
    .Y(_02315_),
    .B1(net4668));
 sg13g2_a22oi_1 _16316_ (.Y(_02316_),
    .B1(net4515),
    .B2(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .A2(net4520),
    .A1(\soc_inst.cpu_core.register_file.registers[5][29] ));
 sg13g2_a22oi_1 _16317_ (.Y(_02317_),
    .B1(net4460),
    .B2(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .A2(net4480),
    .A1(\soc_inst.cpu_core.register_file.registers[8][29] ));
 sg13g2_nand3_1 _16318_ (.B(_02316_),
    .C(_02317_),
    .A(_02315_),
    .Y(_02318_));
 sg13g2_a221oi_1 _16319_ (.B2(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .C1(_02318_),
    .B1(net4455),
    .A1(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .Y(_02319_),
    .A2(net4495));
 sg13g2_a22oi_1 _16320_ (.Y(_02320_),
    .B1(net4465),
    .B2(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .A2(net4470),
    .A1(\soc_inst.cpu_core.register_file.registers[12][29] ));
 sg13g2_nand3_1 _16321_ (.B(_02314_),
    .C(_02320_),
    .A(_02313_),
    .Y(_02321_));
 sg13g2_a221oi_1 _16322_ (.B2(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .C1(_02321_),
    .B1(net4475),
    .A1(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .Y(_02322_),
    .A2(net4510));
 sg13g2_a221oi_1 _16323_ (.B2(_02322_),
    .C1(net4076),
    .B1(_02319_),
    .A1(_05732_),
    .Y(_02323_),
    .A2(net4669));
 sg13g2_a21o_1 _16324_ (.A2(net1607),
    .A1(net4904),
    .B1(_02323_),
    .X(_01126_));
 sg13g2_nor2_1 _16325_ (.A(net2385),
    .B(net4665),
    .Y(_02324_));
 sg13g2_nand2_1 _16326_ (.Y(_02325_),
    .A(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .B(net4488));
 sg13g2_a22oi_1 _16327_ (.Y(_02326_),
    .B1(net4462),
    .B2(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .A2(net4512),
    .A1(\soc_inst.cpu_core.register_file.registers[10][30] ));
 sg13g2_a22oi_1 _16328_ (.Y(_02327_),
    .B1(net4517),
    .B2(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .A2(net4521),
    .A1(\soc_inst.cpu_core.register_file.registers[5][30] ));
 sg13g2_a21oi_1 _16329_ (.A1(\soc_inst.cpu_core.register_file.registers[6][30] ),
    .A2(net4502),
    .Y(_02328_),
    .B1(net4672));
 sg13g2_a22oi_1 _16330_ (.Y(_02329_),
    .B1(net4467),
    .B2(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .A2(net4493),
    .A1(\soc_inst.cpu_core.register_file.registers[9][30] ));
 sg13g2_nand4_1 _16331_ (.B(_02327_),
    .C(_02328_),
    .A(_02326_),
    .Y(_02330_),
    .D(_02329_));
 sg13g2_a22oi_1 _16332_ (.Y(_02331_),
    .B1(net4472),
    .B2(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .A2(net4482),
    .A1(\soc_inst.cpu_core.register_file.registers[8][30] ));
 sg13g2_a22oi_1 _16333_ (.Y(_02332_),
    .B1(net4477),
    .B2(\soc_inst.cpu_core.register_file.registers[2][30] ),
    .A2(net4507),
    .A1(\soc_inst.cpu_core.register_file.registers[3][30] ));
 sg13g2_a22oi_1 _16334_ (.Y(_02333_),
    .B1(net4457),
    .B2(\soc_inst.cpu_core.register_file.registers[7][30] ),
    .A2(net4497),
    .A1(\soc_inst.cpu_core.register_file.registers[11][30] ));
 sg13g2_nand4_1 _16335_ (.B(_02331_),
    .C(_02332_),
    .A(_02325_),
    .Y(_02334_),
    .D(_02333_));
 sg13g2_nor2_1 _16336_ (.A(_02330_),
    .B(_02334_),
    .Y(_02335_));
 sg13g2_nor3_2 _16337_ (.A(net4077),
    .B(_02324_),
    .C(_02335_),
    .Y(_02336_));
 sg13g2_a21o_1 _16338_ (.A2(net2756),
    .A1(net4903),
    .B1(_02336_),
    .X(_01127_));
 sg13g2_nand2_1 _16339_ (.Y(_02337_),
    .A(\soc_inst.cpu_core.register_file.registers[6][31] ),
    .B(net4499));
 sg13g2_a22oi_1 _16340_ (.Y(_02338_),
    .B1(net4494),
    .B2(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .A2(net4514),
    .A1(\soc_inst.cpu_core.register_file.registers[13][31] ));
 sg13g2_a22oi_1 _16341_ (.Y(_02339_),
    .B1(net4474),
    .B2(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .A2(net4489),
    .A1(\soc_inst.cpu_core.register_file.registers[9][31] ));
 sg13g2_a21oi_1 _16342_ (.A1(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .A2(net4509),
    .Y(_02340_),
    .B1(net4670));
 sg13g2_a22oi_1 _16343_ (.Y(_02341_),
    .B1(net4464),
    .B2(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .A2(net4504),
    .A1(\soc_inst.cpu_core.register_file.registers[3][31] ));
 sg13g2_nand4_1 _16344_ (.B(_02339_),
    .C(_02340_),
    .A(_02338_),
    .Y(_02342_),
    .D(_02341_));
 sg13g2_a22oi_1 _16345_ (.Y(_02343_),
    .B1(net4484),
    .B2(\soc_inst.cpu_core.register_file.registers[4][31] ),
    .A2(net4519),
    .A1(\soc_inst.cpu_core.register_file.registers[5][31] ));
 sg13g2_a22oi_1 _16346_ (.Y(_02344_),
    .B1(net4454),
    .B2(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .A2(net4469),
    .A1(\soc_inst.cpu_core.register_file.registers[12][31] ));
 sg13g2_a22oi_1 _16347_ (.Y(_02345_),
    .B1(net4459),
    .B2(\soc_inst.cpu_core.register_file.registers[14][31] ),
    .A2(net4479),
    .A1(\soc_inst.cpu_core.register_file.registers[8][31] ));
 sg13g2_nand4_1 _16348_ (.B(_02343_),
    .C(_02344_),
    .A(_02337_),
    .Y(_02346_),
    .D(_02345_));
 sg13g2_nor2_2 _16349_ (.A(_02342_),
    .B(_02346_),
    .Y(_02347_));
 sg13g2_nor2_1 _16350_ (.A(net1193),
    .B(net4666),
    .Y(_02348_));
 sg13g2_nor3_2 _16351_ (.A(net4076),
    .B(_02347_),
    .C(_02348_),
    .Y(_02349_));
 sg13g2_a21o_1 _16352_ (.A2(net2934),
    .A1(net4902),
    .B1(_02349_),
    .X(_01128_));
 sg13g2_nor2_1 _16353_ (.A(_00265_),
    .B(_00264_),
    .Y(_02350_));
 sg13g2_nor4_2 _16354_ (.A(net1426),
    .B(net1676),
    .C(\soc_inst.cpu_core.if_instr[3] ),
    .Y(_02351_),
    .D(net2801));
 sg13g2_nor2b_1 _16355_ (.A(net5015),
    .B_N(_02351_),
    .Y(_02352_));
 sg13g2_nand2b_2 _16356_ (.Y(_02353_),
    .B(_02351_),
    .A_N(net5015));
 sg13g2_nand2_2 _16357_ (.Y(_02354_),
    .A(\soc_inst.cpu_core.if_instr[2] ),
    .B(_02350_));
 sg13g2_inv_1 _16358_ (.Y(_02355_),
    .A(_02354_));
 sg13g2_and4_1 _16359_ (.A(net5017),
    .B(\soc_inst.cpu_core.if_instr[5] ),
    .C(net5014),
    .D(_02355_),
    .X(_02356_));
 sg13g2_nand4_1 _16360_ (.B(net2608),
    .C(net5013),
    .A(net5017),
    .Y(_02357_),
    .D(_02355_));
 sg13g2_nor2_1 _16361_ (.A(\soc_inst.cpu_core.if_instr[3] ),
    .B(_02357_),
    .Y(_02358_));
 sg13g2_a21oi_2 _16362_ (.B1(_02358_),
    .Y(_02359_),
    .A2(net4452),
    .A1(_05721_));
 sg13g2_nor2_1 _16363_ (.A(net5006),
    .B(_02359_),
    .Y(_02360_));
 sg13g2_nand2_1 _16364_ (.Y(_02361_),
    .A(net5017),
    .B(net4452));
 sg13g2_o21ai_1 _16365_ (.B1(_02359_),
    .Y(_02362_),
    .A1(_05722_),
    .A2(_02361_));
 sg13g2_nor2b_2 _16366_ (.A(_02360_),
    .B_N(_02362_),
    .Y(_02363_));
 sg13g2_a22oi_1 _16367_ (.Y(_02364_),
    .B1(net4131),
    .B2(_02363_),
    .A2(net2517),
    .A1(net4931));
 sg13g2_inv_1 _16368_ (.Y(_01129_),
    .A(_02364_));
 sg13g2_and2_1 _16369_ (.A(\soc_inst.cpu_core.if_instr[3] ),
    .B(_02356_),
    .X(_02365_));
 sg13g2_inv_2 _16370_ (.Y(_02366_),
    .A(net4073));
 sg13g2_nand2_2 _16371_ (.Y(_02367_),
    .A(_02359_),
    .B(_02366_));
 sg13g2_and3_2 _16372_ (.X(_02368_),
    .A(_00266_),
    .B(\soc_inst.cpu_core.if_instr[5] ),
    .C(_02351_));
 sg13g2_a22oi_1 _16373_ (.Y(_02369_),
    .B1(_02368_),
    .B2(net568),
    .A2(_02367_),
    .A1(net5004));
 sg13g2_nand2_1 _16374_ (.Y(_02370_),
    .A(net4931),
    .B(net1915));
 sg13g2_o21ai_1 _16375_ (.B1(_02370_),
    .Y(_01130_),
    .A1(net4122),
    .A2(_02369_));
 sg13g2_a22oi_1 _16376_ (.Y(_02371_),
    .B1(_02368_),
    .B2(net1457),
    .A2(_02367_),
    .A1(net5002));
 sg13g2_nand2_1 _16377_ (.Y(_02372_),
    .A(net4935),
    .B(net1592));
 sg13g2_o21ai_1 _16378_ (.B1(_02372_),
    .Y(_01131_),
    .A1(net4122),
    .A2(_02371_));
 sg13g2_a22oi_1 _16379_ (.Y(_02373_),
    .B1(_02368_),
    .B2(net667),
    .A2(_02367_),
    .A1(net5000));
 sg13g2_nand2_1 _16380_ (.Y(_02374_),
    .A(net4936),
    .B(net1959));
 sg13g2_o21ai_1 _16381_ (.B1(_02374_),
    .Y(_01132_),
    .A1(net4122),
    .A2(_02373_));
 sg13g2_a22oi_1 _16382_ (.Y(_02375_),
    .B1(_02368_),
    .B2(net706),
    .A2(_02367_),
    .A1(\soc_inst.cpu_core.if_imm12[4] ));
 sg13g2_nand2_1 _16383_ (.Y(_02376_),
    .A(net4933),
    .B(net2019));
 sg13g2_o21ai_1 _16384_ (.B1(_02376_),
    .Y(_01133_),
    .A1(net4123),
    .A2(_02375_));
 sg13g2_nand2_1 _16385_ (.Y(_02377_),
    .A(net4936),
    .B(net2238));
 sg13g2_or2_1 _16386_ (.X(_02378_),
    .B(_02368_),
    .A(_02367_));
 sg13g2_nand2_2 _16387_ (.Y(_02379_),
    .A(\soc_inst.cpu_core.if_funct7[0] ),
    .B(_02378_));
 sg13g2_o21ai_1 _16388_ (.B1(_02377_),
    .Y(_01134_),
    .A1(net4122),
    .A2(_02379_));
 sg13g2_nand2_1 _16389_ (.Y(_02380_),
    .A(net4933),
    .B(net2091));
 sg13g2_nand2_1 _16390_ (.Y(_02381_),
    .A(net1597),
    .B(_02378_));
 sg13g2_o21ai_1 _16391_ (.B1(_02380_),
    .Y(_01135_),
    .A1(net4122),
    .A2(_02381_));
 sg13g2_nand2_1 _16392_ (.Y(_02382_),
    .A(net4931),
    .B(net2036));
 sg13g2_nand2_1 _16393_ (.Y(_02383_),
    .A(\soc_inst.cpu_core.if_funct7[2] ),
    .B(_02378_));
 sg13g2_o21ai_1 _16394_ (.B1(_02382_),
    .Y(_01136_),
    .A1(net4122),
    .A2(_02383_));
 sg13g2_nand2_1 _16395_ (.Y(_02384_),
    .A(net4935),
    .B(net1490));
 sg13g2_nand2_2 _16396_ (.Y(_02385_),
    .A(net2077),
    .B(_02378_));
 sg13g2_o21ai_1 _16397_ (.B1(_02384_),
    .Y(_01137_),
    .A1(net4122),
    .A2(_02385_));
 sg13g2_nand2_1 _16398_ (.Y(_02386_),
    .A(net4933),
    .B(net1581));
 sg13g2_nand2_2 _16399_ (.Y(_02387_),
    .A(net2976),
    .B(_02378_));
 sg13g2_o21ai_1 _16400_ (.B1(_02386_),
    .Y(_01138_),
    .A1(net4122),
    .A2(_02387_));
 sg13g2_nand2_1 _16401_ (.Y(_02388_),
    .A(net4933),
    .B(net2166));
 sg13g2_nand2_1 _16402_ (.Y(_02389_),
    .A(net2122),
    .B(_02378_));
 sg13g2_o21ai_1 _16403_ (.B1(_02388_),
    .Y(_01139_),
    .A1(net4123),
    .A2(_02389_));
 sg13g2_nand4_1 _16404_ (.B(net905),
    .C(net4130),
    .A(net5014),
    .Y(_02390_),
    .D(_02368_));
 sg13g2_o21ai_1 _16405_ (.B1(_02361_),
    .Y(_02391_),
    .A1(\soc_inst.cpu_core.if_instr[5] ),
    .A2(_02353_));
 sg13g2_o21ai_1 _16406_ (.B1(\soc_inst.cpu_core.if_funct7[6] ),
    .Y(_02392_),
    .A1(_02358_),
    .A2(_02391_));
 sg13g2_nand2_1 _16407_ (.Y(_02393_),
    .A(net5005),
    .B(net4074));
 sg13g2_and2_1 _16408_ (.A(_02392_),
    .B(_02393_),
    .X(_02394_));
 sg13g2_nand2_1 _16409_ (.Y(_02395_),
    .A(_02392_),
    .B(_02393_));
 sg13g2_a22oi_1 _16410_ (.Y(_02396_),
    .B1(net4133),
    .B2(_02395_),
    .A2(net1061),
    .A1(net4927));
 sg13g2_nand2_1 _16411_ (.Y(_01140_),
    .A(_02390_),
    .B(net1062));
 sg13g2_nand2b_1 _16412_ (.Y(_02397_),
    .B(_02359_),
    .A_N(_02368_));
 sg13g2_and2_1 _16413_ (.A(\soc_inst.cpu_core.if_funct7[6] ),
    .B(_02397_),
    .X(_02398_));
 sg13g2_nand2_2 _16414_ (.Y(_02399_),
    .A(\soc_inst.cpu_core.if_funct7[6] ),
    .B(_02397_));
 sg13g2_or4_1 _16415_ (.A(net5017),
    .B(\soc_inst.cpu_core.if_instr[3] ),
    .C(net5014),
    .D(_02354_),
    .X(_02400_));
 sg13g2_inv_1 _16416_ (.Y(_02401_),
    .A(_02400_));
 sg13g2_nand2_1 _16417_ (.Y(_02402_),
    .A(_02366_),
    .B(_02400_));
 sg13g2_a21oi_1 _16418_ (.A1(net2982),
    .A2(net3970),
    .Y(_02403_),
    .B1(_02398_));
 sg13g2_nand2_1 _16419_ (.Y(_02404_),
    .A(net4908),
    .B(net1803));
 sg13g2_o21ai_1 _16420_ (.B1(_02404_),
    .Y(_01141_),
    .A1(net4123),
    .A2(_02403_));
 sg13g2_a21oi_1 _16421_ (.A1(net2276),
    .A2(net3970),
    .Y(_02405_),
    .B1(_02398_));
 sg13g2_nand2_1 _16422_ (.Y(_02406_),
    .A(net4902),
    .B(net2493));
 sg13g2_o21ai_1 _16423_ (.B1(_02406_),
    .Y(_01142_),
    .A1(net4124),
    .A2(_02405_));
 sg13g2_a21oi_1 _16424_ (.A1(net2222),
    .A2(net3970),
    .Y(_02407_),
    .B1(_02398_));
 sg13g2_nand2_1 _16425_ (.Y(_02408_),
    .A(net4903),
    .B(net2280));
 sg13g2_o21ai_1 _16426_ (.B1(_02408_),
    .Y(_01143_),
    .A1(net4123),
    .A2(_02407_));
 sg13g2_a21oi_1 _16427_ (.A1(net5010),
    .A2(_02402_),
    .Y(_02409_),
    .B1(_02398_));
 sg13g2_nand2_1 _16428_ (.Y(_02410_),
    .A(net4904),
    .B(net2332));
 sg13g2_o21ai_1 _16429_ (.B1(_02410_),
    .Y(_01144_),
    .A1(net4124),
    .A2(_02409_));
 sg13g2_a21oi_1 _16430_ (.A1(\soc_inst.cpu_core.if_instr[16] ),
    .A2(net3970),
    .Y(_02411_),
    .B1(_02398_));
 sg13g2_nand2_1 _16431_ (.Y(_02412_),
    .A(net4898),
    .B(net2189));
 sg13g2_o21ai_1 _16432_ (.B1(_02412_),
    .Y(_01145_),
    .A1(net4124),
    .A2(_02411_));
 sg13g2_a21oi_1 _16433_ (.A1(net1239),
    .A2(net3970),
    .Y(_02413_),
    .B1(_02398_));
 sg13g2_nand2_1 _16434_ (.Y(_02414_),
    .A(net4899),
    .B(net2172));
 sg13g2_o21ai_1 _16435_ (.B1(_02414_),
    .Y(_01146_),
    .A1(net4124),
    .A2(_02413_));
 sg13g2_a21oi_1 _16436_ (.A1(net5007),
    .A2(net3970),
    .Y(_02415_),
    .B1(_02398_));
 sg13g2_nand2_1 _16437_ (.Y(_02416_),
    .A(net4899),
    .B(net2089));
 sg13g2_o21ai_1 _16438_ (.B1(_02416_),
    .Y(_01147_),
    .A1(net4124),
    .A2(_02415_));
 sg13g2_a21oi_1 _16439_ (.A1(\soc_inst.cpu_core.if_instr[19] ),
    .A2(net3970),
    .Y(_02417_),
    .B1(_02398_));
 sg13g2_nand2_1 _16440_ (.Y(_02418_),
    .A(net4897),
    .B(net1251));
 sg13g2_o21ai_1 _16441_ (.B1(_02418_),
    .Y(_01148_),
    .A1(net4124),
    .A2(_02417_));
 sg13g2_o21ai_1 _16442_ (.B1(net3970),
    .Y(_02419_),
    .A1(\soc_inst.cpu_core.if_funct7[6] ),
    .A2(_02366_));
 sg13g2_nor2_1 _16443_ (.A(net5006),
    .B(net4073),
    .Y(_02420_));
 sg13g2_o21ai_1 _16444_ (.B1(net3881),
    .Y(_02421_),
    .A1(net3880),
    .A2(_02420_));
 sg13g2_inv_1 _16445_ (.Y(_02422_),
    .A(_02421_));
 sg13g2_a22oi_1 _16446_ (.Y(_02423_),
    .B1(net4127),
    .B2(_02421_),
    .A2(net2835),
    .A1(net4897));
 sg13g2_inv_1 _16447_ (.Y(_01149_),
    .A(_02423_));
 sg13g2_nor2_1 _16448_ (.A(net5004),
    .B(net4073),
    .Y(_02424_));
 sg13g2_o21ai_1 _16449_ (.B1(net3881),
    .Y(_02425_),
    .A1(net3880),
    .A2(_02424_));
 sg13g2_inv_1 _16450_ (.Y(_02426_),
    .A(_02425_));
 sg13g2_a22oi_1 _16451_ (.Y(_02427_),
    .B1(net4125),
    .B2(_02425_),
    .A2(net2731),
    .A1(net4884));
 sg13g2_inv_1 _16452_ (.Y(_01150_),
    .A(_02427_));
 sg13g2_nor2_1 _16453_ (.A(net5002),
    .B(net4073),
    .Y(_02428_));
 sg13g2_o21ai_1 _16454_ (.B1(net3881),
    .Y(_02429_),
    .A1(net3880),
    .A2(_02428_));
 sg13g2_inv_1 _16455_ (.Y(_02430_),
    .A(_02429_));
 sg13g2_a22oi_1 _16456_ (.Y(_02431_),
    .B1(net4125),
    .B2(_02429_),
    .A2(net2708),
    .A1(net4897));
 sg13g2_inv_1 _16457_ (.Y(_01151_),
    .A(_02431_));
 sg13g2_nor2_1 _16458_ (.A(net5000),
    .B(net4073),
    .Y(_02432_));
 sg13g2_o21ai_1 _16459_ (.B1(net3881),
    .Y(_02433_),
    .A1(net3880),
    .A2(_02432_));
 sg13g2_inv_1 _16460_ (.Y(_02434_),
    .A(_02433_));
 sg13g2_a22oi_1 _16461_ (.Y(_02435_),
    .B1(net4125),
    .B2(_02433_),
    .A2(net2703),
    .A1(net4898));
 sg13g2_inv_1 _16462_ (.Y(_01152_),
    .A(_02435_));
 sg13g2_nor2_1 _16463_ (.A(net2717),
    .B(net4073),
    .Y(_02436_));
 sg13g2_o21ai_1 _16464_ (.B1(net3881),
    .Y(_02437_),
    .A1(net3880),
    .A2(_02436_));
 sg13g2_inv_1 _16465_ (.Y(_02438_),
    .A(_02437_));
 sg13g2_a22oi_1 _16466_ (.Y(_02439_),
    .B1(net4125),
    .B2(_02437_),
    .A2(net2814),
    .A1(net4904));
 sg13g2_inv_1 _16467_ (.Y(_01153_),
    .A(_02439_));
 sg13g2_nor2_1 _16468_ (.A(net2251),
    .B(net4074),
    .Y(_02440_));
 sg13g2_o21ai_1 _16469_ (.B1(net3881),
    .Y(_02441_),
    .A1(net3880),
    .A2(_02440_));
 sg13g2_inv_1 _16470_ (.Y(_02442_),
    .A(_02441_));
 sg13g2_a22oi_1 _16471_ (.Y(_02443_),
    .B1(net4125),
    .B2(_02441_),
    .A2(net2623),
    .A1(net4885));
 sg13g2_inv_1 _16472_ (.Y(_01154_),
    .A(_02443_));
 sg13g2_nor2_1 _16473_ (.A(net1597),
    .B(net4074),
    .Y(_02444_));
 sg13g2_o21ai_1 _16474_ (.B1(net3881),
    .Y(_02445_),
    .A1(net3880),
    .A2(_02444_));
 sg13g2_inv_1 _16475_ (.Y(_02446_),
    .A(_02445_));
 sg13g2_a22oi_1 _16476_ (.Y(_02447_),
    .B1(net4126),
    .B2(_02445_),
    .A2(net2713),
    .A1(net4904));
 sg13g2_inv_1 _16477_ (.Y(_01155_),
    .A(_02447_));
 sg13g2_nor2_1 _16478_ (.A(\soc_inst.cpu_core.if_funct7[2] ),
    .B(net4074),
    .Y(_02448_));
 sg13g2_o21ai_1 _16479_ (.B1(_02399_),
    .Y(_02449_),
    .A1(_02419_),
    .A2(_02448_));
 sg13g2_inv_1 _16480_ (.Y(_02450_),
    .A(_02449_));
 sg13g2_a22oi_1 _16481_ (.Y(_02451_),
    .B1(net4126),
    .B2(_02449_),
    .A2(net2650),
    .A1(net4904));
 sg13g2_inv_1 _16482_ (.Y(_01156_),
    .A(net2651));
 sg13g2_nor2_1 _16483_ (.A(net2077),
    .B(net4073),
    .Y(_02452_));
 sg13g2_o21ai_1 _16484_ (.B1(net3881),
    .Y(_02453_),
    .A1(net3880),
    .A2(_02452_));
 sg13g2_inv_1 _16485_ (.Y(_02454_),
    .A(_02453_));
 sg13g2_a22oi_1 _16486_ (.Y(_02455_),
    .B1(net4125),
    .B2(_02453_),
    .A2(net2701),
    .A1(net4898));
 sg13g2_inv_1 _16487_ (.Y(_01157_),
    .A(_02455_));
 sg13g2_nor2_1 _16488_ (.A(\soc_inst.cpu_core.if_funct7[4] ),
    .B(net4073),
    .Y(_02456_));
 sg13g2_o21ai_1 _16489_ (.B1(_02399_),
    .Y(_02457_),
    .A1(_02419_),
    .A2(_02456_));
 sg13g2_inv_1 _16490_ (.Y(_02458_),
    .A(_02457_));
 sg13g2_a22oi_1 _16491_ (.Y(_02459_),
    .B1(net4126),
    .B2(_02457_),
    .A2(net2605),
    .A1(net4885));
 sg13g2_inv_1 _16492_ (.Y(_01158_),
    .A(net2606));
 sg13g2_nor2_1 _16493_ (.A(net2122),
    .B(net4074),
    .Y(_02460_));
 sg13g2_o21ai_1 _16494_ (.B1(_02399_),
    .Y(_02461_),
    .A1(_02419_),
    .A2(_02460_));
 sg13g2_inv_1 _16495_ (.Y(_02462_),
    .A(_02461_));
 sg13g2_a22oi_1 _16496_ (.Y(_02463_),
    .B1(net4129),
    .B2(_02461_),
    .A2(net2360),
    .A1(net4902));
 sg13g2_inv_1 _16497_ (.Y(_01159_),
    .A(net2361));
 sg13g2_nand2_1 _16498_ (.Y(_02464_),
    .A(net4902),
    .B(net993));
 sg13g2_o21ai_1 _16499_ (.B1(\soc_inst.cpu_core.if_funct7[6] ),
    .Y(_02465_),
    .A1(_02378_),
    .A2(_02401_));
 sg13g2_o21ai_1 _16500_ (.B1(_02464_),
    .Y(_01160_),
    .A1(net4123),
    .A2(_02465_));
 sg13g2_nor2_1 _16501_ (.A(net4970),
    .B(_05543_),
    .Y(_02466_));
 sg13g2_a22oi_1 _16502_ (.Y(_02467_),
    .B1(net3862),
    .B2(_02466_),
    .A2(net2764),
    .A1(net4970));
 sg13g2_inv_1 _16503_ (.Y(_01161_),
    .A(_02467_));
 sg13g2_nor2_1 _16504_ (.A(net5017),
    .B(_02353_),
    .Y(_02468_));
 sg13g2_nand4_1 _16505_ (.B(_02357_),
    .C(_02361_),
    .A(net4130),
    .Y(_02469_),
    .D(_02400_));
 sg13g2_a21oi_1 _16506_ (.A1(_05725_),
    .A2(_02468_),
    .Y(_02470_),
    .B1(_02469_));
 sg13g2_a21o_1 _16507_ (.A2(net2745),
    .A1(net4886),
    .B1(_02470_),
    .X(_01162_));
 sg13g2_nor3_1 _16508_ (.A(net5017),
    .B(net2276),
    .C(_02353_),
    .Y(_02471_));
 sg13g2_nand2_1 _16509_ (.Y(_02472_),
    .A(net4885),
    .B(net2349));
 sg13g2_o21ai_1 _16510_ (.B1(_02472_),
    .Y(_01163_),
    .A1(_02469_),
    .A2(_02471_));
 sg13g2_nor3_1 _16511_ (.A(net5017),
    .B(net2222),
    .C(_02353_),
    .Y(_02473_));
 sg13g2_nand2_1 _16512_ (.Y(_02474_),
    .A(net4885),
    .B(net2423));
 sg13g2_o21ai_1 _16513_ (.B1(_02474_),
    .Y(_01164_),
    .A1(_02469_),
    .A2(_02473_));
 sg13g2_nand3b_1 _16514_ (.B(net2222),
    .C(net2122),
    .Y(_02475_),
    .A_N(net2276));
 sg13g2_nand2_1 _16515_ (.Y(_02476_),
    .A(_02468_),
    .B(_02475_));
 sg13g2_nand2_1 _16516_ (.Y(_02477_),
    .A(\soc_inst.cpu_core.if_instr[5] ),
    .B(_02468_));
 sg13g2_a22oi_1 _16517_ (.Y(_02478_),
    .B1(_02470_),
    .B2(_02476_),
    .A2(net4865),
    .A1(net4885));
 sg13g2_o21ai_1 _16518_ (.B1(_02478_),
    .Y(_01165_),
    .A1(_09589_),
    .A2(net4114));
 sg13g2_a21oi_1 _16519_ (.A1(_05721_),
    .A2(_02401_),
    .Y(_02479_),
    .B1(_02356_));
 sg13g2_nor2_1 _16520_ (.A(_09209_),
    .B(_02479_),
    .Y(_02480_));
 sg13g2_nor2_2 _16521_ (.A(net4974),
    .B(_05520_),
    .Y(_02481_));
 sg13g2_a22oi_1 _16522_ (.Y(_02482_),
    .B1(net4020),
    .B2(_02481_),
    .A2(net4451),
    .A1(_09625_));
 sg13g2_o21ai_1 _16523_ (.B1(_02482_),
    .Y(_01166_),
    .A1(net4747),
    .A2(_05840_));
 sg13g2_nor2_2 _16524_ (.A(net4973),
    .B(_05519_),
    .Y(_02483_));
 sg13g2_a22oi_1 _16525_ (.Y(_02484_),
    .B1(net4020),
    .B2(_02483_),
    .A2(net4450),
    .A1(_09636_));
 sg13g2_o21ai_1 _16526_ (.B1(_02484_),
    .Y(_01167_),
    .A1(net4748),
    .A2(_05838_));
 sg13g2_nor2_2 _16527_ (.A(net4975),
    .B(_05522_),
    .Y(_02485_));
 sg13g2_a22oi_1 _16528_ (.Y(_02486_),
    .B1(net4021),
    .B2(_02485_),
    .A2(net4452),
    .A1(_09647_));
 sg13g2_o21ai_1 _16529_ (.B1(_02486_),
    .Y(_01168_),
    .A1(net4750),
    .A2(_05836_));
 sg13g2_nor2_2 _16530_ (.A(net4974),
    .B(_05521_),
    .Y(_02487_));
 sg13g2_a22oi_1 _16531_ (.Y(_02488_),
    .B1(net4020),
    .B2(_02487_),
    .A2(net4453),
    .A1(_09658_));
 sg13g2_o21ai_1 _16532_ (.B1(_02488_),
    .Y(_01169_),
    .A1(net4748),
    .A2(_05834_));
 sg13g2_nor2_2 _16533_ (.A(net4975),
    .B(_05523_),
    .Y(_02489_));
 sg13g2_a22oi_1 _16534_ (.Y(_02490_),
    .B1(net4021),
    .B2(_02489_),
    .A2(net4450),
    .A1(_09669_));
 sg13g2_o21ai_1 _16535_ (.B1(_02490_),
    .Y(_01170_),
    .A1(net4747),
    .A2(_05832_));
 sg13g2_nor2_2 _16536_ (.A(net4974),
    .B(_05524_),
    .Y(_02491_));
 sg13g2_a22oi_1 _16537_ (.Y(_02492_),
    .B1(net4020),
    .B2(_02491_),
    .A2(net4450),
    .A1(_09682_));
 sg13g2_o21ai_1 _16538_ (.B1(_02492_),
    .Y(_01171_),
    .A1(net4747),
    .A2(_05830_));
 sg13g2_nor2_2 _16539_ (.A(net4975),
    .B(_05525_),
    .Y(_02493_));
 sg13g2_a22oi_1 _16540_ (.Y(_02494_),
    .B1(net4020),
    .B2(_02493_),
    .A2(net4450),
    .A1(_09695_));
 sg13g2_o21ai_1 _16541_ (.B1(_02494_),
    .Y(_01172_),
    .A1(net4747),
    .A2(_05828_));
 sg13g2_nor2_2 _16542_ (.A(net4975),
    .B(_05526_),
    .Y(_02495_));
 sg13g2_a22oi_1 _16543_ (.Y(_02496_),
    .B1(net4020),
    .B2(_02495_),
    .A2(net4450),
    .A1(_09706_));
 sg13g2_o21ai_1 _16544_ (.B1(_02496_),
    .Y(_01173_),
    .A1(net4747),
    .A2(_05826_));
 sg13g2_nor2_2 _16545_ (.A(net4963),
    .B(_05527_),
    .Y(_02497_));
 sg13g2_a22oi_1 _16546_ (.Y(_02498_),
    .B1(net4020),
    .B2(_02497_),
    .A2(net4452),
    .A1(_09717_));
 sg13g2_o21ai_1 _16547_ (.B1(_02498_),
    .Y(_01174_),
    .A1(net4748),
    .A2(_05824_));
 sg13g2_nor2_2 _16548_ (.A(net4972),
    .B(_05528_),
    .Y(_02499_));
 sg13g2_a22oi_1 _16549_ (.Y(_02500_),
    .B1(net4020),
    .B2(_02499_),
    .A2(net4451),
    .A1(_09728_));
 sg13g2_o21ai_1 _16550_ (.B1(_02500_),
    .Y(_01175_),
    .A1(net4747),
    .A2(_05822_));
 sg13g2_nor2_2 _16551_ (.A(net4962),
    .B(_05529_),
    .Y(_02501_));
 sg13g2_a22oi_1 _16552_ (.Y(_02502_),
    .B1(net4021),
    .B2(_02501_),
    .A2(net4452),
    .A1(_09739_));
 sg13g2_o21ai_1 _16553_ (.B1(_02502_),
    .Y(_01176_),
    .A1(net4742),
    .A2(_05820_));
 sg13g2_nor2_2 _16554_ (.A(net4962),
    .B(_05530_),
    .Y(_02503_));
 sg13g2_a22oi_1 _16555_ (.Y(_02504_),
    .B1(net4021),
    .B2(_02503_),
    .A2(net4452),
    .A1(_09750_));
 sg13g2_o21ai_1 _16556_ (.B1(_02504_),
    .Y(_01177_),
    .A1(net4748),
    .A2(_05818_));
 sg13g2_nor2_2 _16557_ (.A(net4962),
    .B(_05531_),
    .Y(_02505_));
 sg13g2_a22oi_1 _16558_ (.Y(_02506_),
    .B1(net4021),
    .B2(_02505_),
    .A2(net4452),
    .A1(_09761_));
 sg13g2_o21ai_1 _16559_ (.B1(_02506_),
    .Y(_01178_),
    .A1(net4746),
    .A2(_05816_));
 sg13g2_nor2_2 _16560_ (.A(net4961),
    .B(_05532_),
    .Y(_02507_));
 sg13g2_a22oi_1 _16561_ (.Y(_02508_),
    .B1(net4019),
    .B2(_02507_),
    .A2(net4451),
    .A1(_09772_));
 sg13g2_o21ai_1 _16562_ (.B1(_02508_),
    .Y(_01179_),
    .A1(net4742),
    .A2(_05814_));
 sg13g2_nor2_2 _16563_ (.A(net4960),
    .B(_05533_),
    .Y(_02509_));
 sg13g2_a22oi_1 _16564_ (.Y(_02510_),
    .B1(net4022),
    .B2(_02509_),
    .A2(net4449),
    .A1(_09783_));
 sg13g2_o21ai_1 _16565_ (.B1(_02510_),
    .Y(_01180_),
    .A1(net4744),
    .A2(_05812_));
 sg13g2_nor2_2 _16566_ (.A(net4960),
    .B(_05534_),
    .Y(_02511_));
 sg13g2_a22oi_1 _16567_ (.Y(_02512_),
    .B1(net4022),
    .B2(_02511_),
    .A2(net4449),
    .A1(_09794_));
 sg13g2_o21ai_1 _16568_ (.B1(_02512_),
    .Y(_01181_),
    .A1(net4745),
    .A2(_05810_));
 sg13g2_nor2_2 _16569_ (.A(net4915),
    .B(_05535_),
    .Y(_02513_));
 sg13g2_a22oi_1 _16570_ (.Y(_02514_),
    .B1(net4019),
    .B2(_02513_),
    .A2(net4448),
    .A1(_09805_));
 sg13g2_o21ai_1 _16571_ (.B1(_02514_),
    .Y(_01182_),
    .A1(net4741),
    .A2(_05808_));
 sg13g2_nor2_2 _16572_ (.A(net4916),
    .B(_05536_),
    .Y(_02515_));
 sg13g2_a22oi_1 _16573_ (.Y(_02516_),
    .B1(net4022),
    .B2(_02515_),
    .A2(net4449),
    .A1(_09816_));
 sg13g2_o21ai_1 _16574_ (.B1(_02516_),
    .Y(_01183_),
    .A1(net4744),
    .A2(_05806_));
 sg13g2_nor2_2 _16575_ (.A(net4916),
    .B(_05537_),
    .Y(_02517_));
 sg13g2_a22oi_1 _16576_ (.Y(_02518_),
    .B1(net4019),
    .B2(_02517_),
    .A2(net4448),
    .A1(_09827_));
 sg13g2_o21ai_1 _16577_ (.B1(_02518_),
    .Y(_01184_),
    .A1(net4741),
    .A2(_05804_));
 sg13g2_nor2_2 _16578_ (.A(net4914),
    .B(_05538_),
    .Y(_02519_));
 sg13g2_a22oi_1 _16579_ (.Y(_02520_),
    .B1(net4019),
    .B2(_02519_),
    .A2(net4449),
    .A1(_09840_));
 sg13g2_o21ai_1 _16580_ (.B1(_02520_),
    .Y(_01185_),
    .A1(net4741),
    .A2(_05802_));
 sg13g2_nor2_2 _16581_ (.A(net4952),
    .B(_05539_),
    .Y(_02521_));
 sg13g2_a22oi_1 _16582_ (.Y(_02522_),
    .B1(net4019),
    .B2(_02521_),
    .A2(net4448),
    .A1(_09851_));
 sg13g2_o21ai_1 _16583_ (.B1(_02522_),
    .Y(_01186_),
    .A1(net4741),
    .A2(_05800_));
 sg13g2_nor2_2 _16584_ (.A(net4952),
    .B(_05540_),
    .Y(_02523_));
 sg13g2_a22oi_1 _16585_ (.Y(_02524_),
    .B1(net4019),
    .B2(_02523_),
    .A2(net4448),
    .A1(_09862_));
 sg13g2_o21ai_1 _16586_ (.B1(_02524_),
    .Y(_01187_),
    .A1(net4741),
    .A2(_05798_));
 sg13g2_nor2_2 _16587_ (.A(net4952),
    .B(_05541_),
    .Y(_02525_));
 sg13g2_a22oi_1 _16588_ (.Y(_02526_),
    .B1(net4019),
    .B2(_02525_),
    .A2(net4448),
    .A1(_09875_));
 sg13g2_o21ai_1 _16589_ (.B1(_02526_),
    .Y(_01188_),
    .A1(net4741),
    .A2(_05796_));
 sg13g2_nor2_2 _16590_ (.A(net4952),
    .B(_05542_),
    .Y(_02527_));
 sg13g2_a22oi_1 _16591_ (.Y(_02528_),
    .B1(net4019),
    .B2(_02527_),
    .A2(net4448),
    .A1(_09886_));
 sg13g2_o21ai_1 _16592_ (.B1(_02528_),
    .Y(_01189_),
    .A1(net4743),
    .A2(_05794_));
 sg13g2_a22oi_1 _16593_ (.Y(_02529_),
    .B1(_09897_),
    .B2(net4451),
    .A2(net2888),
    .A1(net4890));
 sg13g2_inv_1 _16594_ (.Y(_01190_),
    .A(_02529_));
 sg13g2_a22oi_1 _16595_ (.Y(_02530_),
    .B1(_09908_),
    .B2(net4450),
    .A2(net2244),
    .A1(net4890));
 sg13g2_inv_1 _16596_ (.Y(_01191_),
    .A(_02530_));
 sg13g2_a22oi_1 _16597_ (.Y(_02531_),
    .B1(_09919_),
    .B2(net4450),
    .A2(net2454),
    .A1(net4890));
 sg13g2_inv_1 _16598_ (.Y(_01192_),
    .A(_02531_));
 sg13g2_a22oi_1 _16599_ (.Y(_02532_),
    .B1(_09930_),
    .B2(net4451),
    .A2(net2837),
    .A1(net4880));
 sg13g2_inv_1 _16600_ (.Y(_01193_),
    .A(_02532_));
 sg13g2_a22oi_1 _16601_ (.Y(_02533_),
    .B1(_09941_),
    .B2(net4448),
    .A2(net4855),
    .A1(net4882));
 sg13g2_inv_1 _16602_ (.Y(_01194_),
    .A(_02533_));
 sg13g2_a22oi_1 _16603_ (.Y(_02534_),
    .B1(_09952_),
    .B2(net4448),
    .A2(net2893),
    .A1(net4880));
 sg13g2_inv_1 _16604_ (.Y(_01195_),
    .A(_02534_));
 sg13g2_a22oi_1 _16605_ (.Y(_02535_),
    .B1(_09963_),
    .B2(net4450),
    .A2(net2922),
    .A1(net4890));
 sg13g2_inv_1 _16606_ (.Y(_01196_),
    .A(_02535_));
 sg13g2_a22oi_1 _16607_ (.Y(_02536_),
    .B1(_09976_),
    .B2(net4452),
    .A2(net2453),
    .A1(net4891));
 sg13g2_inv_1 _16608_ (.Y(_01197_),
    .A(_02536_));
 sg13g2_nand2b_1 _16609_ (.Y(_02537_),
    .B(_02363_),
    .A_N(net2801));
 sg13g2_nand2_1 _16610_ (.Y(_02538_),
    .A(net4116),
    .B(_02537_));
 sg13g2_and2_1 _16611_ (.A(net4125),
    .B(net4115),
    .X(_02539_));
 sg13g2_o21ai_1 _16612_ (.B1(_02538_),
    .Y(_02540_),
    .A1(_10023_),
    .A2(net4070));
 sg13g2_o21ai_1 _16613_ (.B1(_02540_),
    .Y(_01198_),
    .A1(net4749),
    .A2(_05839_));
 sg13g2_nand2_1 _16614_ (.Y(_02541_),
    .A(net2029),
    .B(_02356_));
 sg13g2_a22oi_1 _16615_ (.Y(_02542_),
    .B1(_02541_),
    .B2(_02353_),
    .A2(_02391_),
    .A1(_02369_));
 sg13g2_o21ai_1 _16616_ (.B1(_02542_),
    .Y(_02543_),
    .A1(_10036_),
    .A2(net4070));
 sg13g2_o21ai_1 _16617_ (.B1(_02543_),
    .Y(_01199_),
    .A1(net4748),
    .A2(_05837_));
 sg13g2_nor2_1 _16618_ (.A(_10049_),
    .B(net4071),
    .Y(_02544_));
 sg13g2_o21ai_1 _16619_ (.B1(_02353_),
    .Y(_02545_),
    .A1(net2029),
    .A2(_02357_));
 sg13g2_a21oi_1 _16620_ (.A1(_02371_),
    .A2(_02391_),
    .Y(_02546_),
    .B1(_02544_));
 sg13g2_a22oi_1 _16621_ (.Y(_02547_),
    .B1(_02545_),
    .B2(_02546_),
    .A2(net4823),
    .A1(net4892));
 sg13g2_inv_1 _16622_ (.Y(_01200_),
    .A(_02547_));
 sg13g2_o21ai_1 _16623_ (.B1(net4117),
    .Y(_02548_),
    .A1(net5015),
    .A2(_02373_));
 sg13g2_o21ai_1 _16624_ (.B1(_02548_),
    .Y(_02549_),
    .A1(_10062_),
    .A2(net4071));
 sg13g2_o21ai_1 _16625_ (.B1(_02549_),
    .Y(_01201_),
    .A1(net4746),
    .A2(net4733));
 sg13g2_o21ai_1 _16626_ (.B1(net4116),
    .Y(_02550_),
    .A1(net5015),
    .A2(_02375_));
 sg13g2_o21ai_1 _16627_ (.B1(_02550_),
    .Y(_02551_),
    .A1(_10073_),
    .A2(net4070));
 sg13g2_o21ai_1 _16628_ (.B1(_02551_),
    .Y(_01202_),
    .A1(net4749),
    .A2(net4737));
 sg13g2_o21ai_1 _16629_ (.B1(net4116),
    .Y(_02552_),
    .A1(net5015),
    .A2(_02379_));
 sg13g2_o21ai_1 _16630_ (.B1(_02552_),
    .Y(_02553_),
    .A1(_10086_),
    .A2(net4070));
 sg13g2_o21ai_1 _16631_ (.B1(_02553_),
    .Y(_01203_),
    .A1(net4747),
    .A2(_05829_));
 sg13g2_o21ai_1 _16632_ (.B1(net4116),
    .Y(_02554_),
    .A1(net5016),
    .A2(_02381_));
 sg13g2_o21ai_1 _16633_ (.B1(_02554_),
    .Y(_02555_),
    .A1(_10099_),
    .A2(net4070));
 sg13g2_o21ai_1 _16634_ (.B1(_02555_),
    .Y(_01204_),
    .A1(net4748),
    .A2(_05827_));
 sg13g2_o21ai_1 _16635_ (.B1(net4117),
    .Y(_02556_),
    .A1(net5015),
    .A2(_02383_));
 sg13g2_o21ai_1 _16636_ (.B1(_02556_),
    .Y(_02557_),
    .A1(_10112_),
    .A2(net4071));
 sg13g2_o21ai_1 _16637_ (.B1(_02557_),
    .Y(_01205_),
    .A1(net4748),
    .A2(_05825_));
 sg13g2_o21ai_1 _16638_ (.B1(net4116),
    .Y(_02558_),
    .A1(net5013),
    .A2(_02385_));
 sg13g2_o21ai_1 _16639_ (.B1(_02558_),
    .Y(_02559_),
    .A1(_10125_),
    .A2(net4070));
 sg13g2_o21ai_1 _16640_ (.B1(_02559_),
    .Y(_01206_),
    .A1(net4743),
    .A2(_05823_));
 sg13g2_o21ai_1 _16641_ (.B1(net4117),
    .Y(_02560_),
    .A1(net5013),
    .A2(_02387_));
 sg13g2_o21ai_1 _16642_ (.B1(_02560_),
    .Y(_02561_),
    .A1(_10136_),
    .A2(net4070));
 sg13g2_o21ai_1 _16643_ (.B1(_02561_),
    .Y(_01207_),
    .A1(net4747),
    .A2(_05821_));
 sg13g2_o21ai_1 _16644_ (.B1(net4117),
    .Y(_02562_),
    .A1(net5013),
    .A2(_02389_));
 sg13g2_o21ai_1 _16645_ (.B1(_02562_),
    .Y(_02563_),
    .A1(_10149_),
    .A2(net4071));
 sg13g2_o21ai_1 _16646_ (.B1(_02563_),
    .Y(_01208_),
    .A1(net4743),
    .A2(_05819_));
 sg13g2_o21ai_1 _16647_ (.B1(net4118),
    .Y(_02564_),
    .A1(net5013),
    .A2(_02394_));
 sg13g2_o21ai_1 _16648_ (.B1(_02564_),
    .Y(_02565_),
    .A1(_10162_),
    .A2(net4072));
 sg13g2_o21ai_1 _16649_ (.B1(_02565_),
    .Y(_01209_),
    .A1(net4750),
    .A2(_05817_));
 sg13g2_o21ai_1 _16650_ (.B1(net4118),
    .Y(_02566_),
    .A1(net5014),
    .A2(_02403_));
 sg13g2_o21ai_1 _16651_ (.B1(_02566_),
    .Y(_02567_),
    .A1(_10175_),
    .A2(net4072));
 sg13g2_o21ai_1 _16652_ (.B1(_02567_),
    .Y(_01210_),
    .A1(net4746),
    .A2(_05815_));
 sg13g2_o21ai_1 _16653_ (.B1(net4114),
    .Y(_02568_),
    .A1(net5012),
    .A2(_02405_));
 sg13g2_o21ai_1 _16654_ (.B1(_02568_),
    .Y(_02569_),
    .A1(_10188_),
    .A2(net4069));
 sg13g2_o21ai_1 _16655_ (.B1(_02569_),
    .Y(_01211_),
    .A1(net4745),
    .A2(_05813_));
 sg13g2_o21ai_1 _16656_ (.B1(net4116),
    .Y(_02570_),
    .A1(net5013),
    .A2(_02407_));
 sg13g2_o21ai_1 _16657_ (.B1(_02570_),
    .Y(_02571_),
    .A1(_10199_),
    .A2(net4071));
 sg13g2_o21ai_1 _16658_ (.B1(_02571_),
    .Y(_01212_),
    .A1(net4746),
    .A2(_05811_));
 sg13g2_o21ai_1 _16659_ (.B1(net4114),
    .Y(_02572_),
    .A1(net5012),
    .A2(_02409_));
 sg13g2_o21ai_1 _16660_ (.B1(_02572_),
    .Y(_02573_),
    .A1(_10210_),
    .A2(net4069));
 sg13g2_o21ai_1 _16661_ (.B1(_02573_),
    .Y(_01213_),
    .A1(net4744),
    .A2(_05809_));
 sg13g2_o21ai_1 _16662_ (.B1(net4113),
    .Y(_02574_),
    .A1(net5011),
    .A2(_02411_));
 sg13g2_o21ai_1 _16663_ (.B1(_02574_),
    .Y(_02575_),
    .A1(_02164_),
    .A2(net4068));
 sg13g2_o21ai_1 _16664_ (.B1(_02575_),
    .Y(_01214_),
    .A1(net4743),
    .A2(_05807_));
 sg13g2_o21ai_1 _16665_ (.B1(net4113),
    .Y(_02576_),
    .A1(net5011),
    .A2(_02413_));
 sg13g2_o21ai_1 _16666_ (.B1(_02576_),
    .Y(_02577_),
    .A1(_02175_),
    .A2(net4068));
 sg13g2_o21ai_1 _16667_ (.B1(_02577_),
    .Y(_01215_),
    .A1(net4744),
    .A2(_05805_));
 sg13g2_o21ai_1 _16668_ (.B1(net4113),
    .Y(_02578_),
    .A1(net5011),
    .A2(_02415_));
 sg13g2_o21ai_1 _16669_ (.B1(_02578_),
    .Y(_02579_),
    .A1(_02188_),
    .A2(net4068));
 sg13g2_o21ai_1 _16670_ (.B1(_02579_),
    .Y(_01216_),
    .A1(net4745),
    .A2(_05803_));
 sg13g2_o21ai_1 _16671_ (.B1(net4113),
    .Y(_02580_),
    .A1(net5011),
    .A2(_02417_));
 sg13g2_o21ai_1 _16672_ (.B1(_02580_),
    .Y(_02581_),
    .A1(_02201_),
    .A2(net4068));
 sg13g2_o21ai_1 _16673_ (.B1(_02581_),
    .Y(_01217_),
    .A1(net4744),
    .A2(_05801_));
 sg13g2_o21ai_1 _16674_ (.B1(net4113),
    .Y(_02582_),
    .A1(net5012),
    .A2(_02422_));
 sg13g2_o21ai_1 _16675_ (.B1(_02582_),
    .Y(_02583_),
    .A1(_02214_),
    .A2(net4069));
 sg13g2_o21ai_1 _16676_ (.B1(_02583_),
    .Y(_01218_),
    .A1(net4744),
    .A2(_05799_));
 sg13g2_o21ai_1 _16677_ (.B1(net4113),
    .Y(_02584_),
    .A1(net5011),
    .A2(_02426_));
 sg13g2_o21ai_1 _16678_ (.B1(_02584_),
    .Y(_02585_),
    .A1(_02225_),
    .A2(net4068));
 sg13g2_o21ai_1 _16679_ (.B1(_02585_),
    .Y(_01219_),
    .A1(net4744),
    .A2(_05797_));
 sg13g2_o21ai_1 _16680_ (.B1(net4114),
    .Y(_02586_),
    .A1(net5011),
    .A2(_02430_));
 sg13g2_o21ai_1 _16681_ (.B1(_02586_),
    .Y(_02587_),
    .A1(_02238_),
    .A2(net4068));
 sg13g2_o21ai_1 _16682_ (.B1(_02587_),
    .Y(_01220_),
    .A1(net4745),
    .A2(_05795_));
 sg13g2_o21ai_1 _16683_ (.B1(net4113),
    .Y(_02588_),
    .A1(net5011),
    .A2(_02434_));
 sg13g2_o21ai_1 _16684_ (.B1(_02588_),
    .Y(_02589_),
    .A1(_02251_),
    .A2(net4068));
 sg13g2_o21ai_1 _16685_ (.B1(_02589_),
    .Y(_01221_),
    .A1(net4744),
    .A2(_05793_));
 sg13g2_o21ai_1 _16686_ (.B1(net4115),
    .Y(_02590_),
    .A1(net5012),
    .A2(_02438_));
 sg13g2_o21ai_1 _16687_ (.B1(_02590_),
    .Y(_02591_),
    .A1(_02262_),
    .A2(net4069));
 sg13g2_o21ai_1 _16688_ (.B1(_02591_),
    .Y(_01222_),
    .A1(net4742),
    .A2(_05792_));
 sg13g2_o21ai_1 _16689_ (.B1(net4116),
    .Y(_02592_),
    .A1(net5013),
    .A2(_02442_));
 sg13g2_o21ai_1 _16690_ (.B1(_02592_),
    .Y(_02593_),
    .A1(_02273_),
    .A2(net4070));
 sg13g2_o21ai_1 _16691_ (.B1(_02593_),
    .Y(_01223_),
    .A1(net4742),
    .A2(_05791_));
 sg13g2_o21ai_1 _16692_ (.B1(net4118),
    .Y(_02594_),
    .A1(net5012),
    .A2(_02446_));
 sg13g2_o21ai_1 _16693_ (.B1(_02594_),
    .Y(_02595_),
    .A1(_02286_),
    .A2(net4072));
 sg13g2_o21ai_1 _16694_ (.B1(_02595_),
    .Y(_01224_),
    .A1(net4746),
    .A2(_05790_));
 sg13g2_o21ai_1 _16695_ (.B1(net4115),
    .Y(_02596_),
    .A1(net5012),
    .A2(_02450_));
 sg13g2_o21ai_1 _16696_ (.B1(_02596_),
    .Y(_02597_),
    .A1(_02299_),
    .A2(net4072));
 sg13g2_o21ai_1 _16697_ (.B1(_02597_),
    .Y(_01225_),
    .A1(net4742),
    .A2(_05789_));
 sg13g2_o21ai_1 _16698_ (.B1(net4113),
    .Y(_02598_),
    .A1(net5011),
    .A2(_02454_));
 sg13g2_o21ai_1 _16699_ (.B1(_02598_),
    .Y(_02599_),
    .A1(_02312_),
    .A2(net4068));
 sg13g2_o21ai_1 _16700_ (.B1(_02599_),
    .Y(_01226_),
    .A1(net4743),
    .A2(_05788_));
 sg13g2_o21ai_1 _16701_ (.B1(net4115),
    .Y(_02600_),
    .A1(\soc_inst.cpu_core.if_instr[6] ),
    .A2(_02458_));
 sg13g2_o21ai_1 _16702_ (.B1(_02600_),
    .Y(_02601_),
    .A1(_02323_),
    .A2(net4069));
 sg13g2_o21ai_1 _16703_ (.B1(_02601_),
    .Y(_01227_),
    .A1(net4742),
    .A2(_05787_));
 sg13g2_o21ai_1 _16704_ (.B1(net4116),
    .Y(_02602_),
    .A1(net5013),
    .A2(_02462_));
 sg13g2_o21ai_1 _16705_ (.B1(_02602_),
    .Y(_02603_),
    .A1(_02336_),
    .A2(net4071));
 sg13g2_o21ai_1 _16706_ (.B1(_02603_),
    .Y(_01228_),
    .A1(net4746),
    .A2(_05786_));
 sg13g2_o21ai_1 _16707_ (.B1(net4118),
    .Y(_02604_),
    .A1(net5012),
    .A2(_02465_));
 sg13g2_o21ai_1 _16708_ (.B1(_02604_),
    .Y(_02605_),
    .A1(_02349_),
    .A2(net4071));
 sg13g2_o21ai_1 _16709_ (.B1(_02605_),
    .Y(_01229_),
    .A1(net4750),
    .A2(_05785_));
 sg13g2_nand2_1 _16710_ (.Y(_02606_),
    .A(net4889),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[0] ));
 sg13g2_o21ai_1 _16711_ (.B1(_02606_),
    .Y(_01230_),
    .A1(net4889),
    .A2(_05763_));
 sg13g2_mux2_1 _16712_ (.A0(net2680),
    .A1(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .S(net4927),
    .X(_01231_));
 sg13g2_mux2_1 _16713_ (.A0(net2557),
    .A1(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .S(net4930),
    .X(_01232_));
 sg13g2_a22oi_1 _16714_ (.Y(_02607_),
    .B1(net2029),
    .B2(net4130),
    .A2(net2158),
    .A1(net4930));
 sg13g2_inv_1 _16715_ (.Y(_01233_),
    .A(_02607_));
 sg13g2_mux2_1 _16716_ (.A0(net2289),
    .A1(_00273_),
    .S(net4980),
    .X(_01234_));
 sg13g2_mux2_1 _16717_ (.A0(net2281),
    .A1(_00274_),
    .S(net4980),
    .X(_01235_));
 sg13g2_nor2_1 _16718_ (.A(net4970),
    .B(\soc_inst.cpu_core.id_instr[2] ),
    .Y(_02608_));
 sg13g2_a21oi_1 _16719_ (.A1(_05475_),
    .A2(net4970),
    .Y(_01236_),
    .B1(_02608_));
 sg13g2_mux2_1 _16720_ (.A0(\soc_inst.cpu_core.id_instr[3] ),
    .A1(net2442),
    .S(net4941),
    .X(_01237_));
 sg13g2_mux2_1 _16721_ (.A0(net2341),
    .A1(_00275_),
    .S(net4980),
    .X(_01238_));
 sg13g2_o21ai_1 _16722_ (.B1(_09212_),
    .Y(_01239_),
    .A1(_05476_),
    .A2(net4752));
 sg13g2_mux2_1 _16723_ (.A0(net4878),
    .A1(net2709),
    .S(net4940),
    .X(_01240_));
 sg13g2_nor2_1 _16724_ (.A(net4927),
    .B(net960),
    .Y(_02609_));
 sg13g2_a21oi_1 _16725_ (.A1(net4892),
    .A2(_05763_),
    .Y(_01241_),
    .B1(_02609_));
 sg13g2_mux2_1 _16726_ (.A0(net2183),
    .A1(\soc_inst.cpu_core.ex_instr[8] ),
    .S(net4928),
    .X(_01242_));
 sg13g2_mux2_1 _16727_ (.A0(net1981),
    .A1(\soc_inst.cpu_core.ex_instr[9] ),
    .S(net4930),
    .X(_01243_));
 sg13g2_mux2_1 _16728_ (.A0(net841),
    .A1(net2086),
    .S(net4928),
    .X(_01244_));
 sg13g2_mux2_1 _16729_ (.A0(net1253),
    .A1(net2066),
    .S(net4939),
    .X(_01245_));
 sg13g2_mux2_1 _16730_ (.A0(\soc_inst.cpu_core.id_funct3[0] ),
    .A1(net2609),
    .S(net4962),
    .X(_01246_));
 sg13g2_mux2_1 _16731_ (.A0(net2498),
    .A1(net2252),
    .S(net4962),
    .X(_01247_));
 sg13g2_mux2_1 _16732_ (.A0(net2386),
    .A1(net1870),
    .S(net4924),
    .X(_01248_));
 sg13g2_mux2_1 _16733_ (.A0(net1048),
    .A1(\soc_inst.cpu_core.ex_instr[15] ),
    .S(net4940),
    .X(_01249_));
 sg13g2_mux2_1 _16734_ (.A0(net2151),
    .A1(\soc_inst.cpu_core.ex_instr[16] ),
    .S(net4926),
    .X(_01250_));
 sg13g2_mux2_1 _16735_ (.A0(net1003),
    .A1(\soc_inst.cpu_core.ex_instr[17] ),
    .S(net4898),
    .X(_01251_));
 sg13g2_mux2_1 _16736_ (.A0(net1064),
    .A1(net1529),
    .S(net4901),
    .X(_01252_));
 sg13g2_mux2_1 _16737_ (.A0(net1242),
    .A1(\soc_inst.cpu_core.ex_instr[19] ),
    .S(net4900),
    .X(_01253_));
 sg13g2_mux2_1 _16738_ (.A0(\soc_inst.cpu_core.id_imm12[0] ),
    .A1(net2041),
    .S(net4958),
    .X(_01254_));
 sg13g2_mux2_1 _16739_ (.A0(\soc_inst.cpu_core.id_imm12[1] ),
    .A1(net2535),
    .S(net4917),
    .X(_01255_));
 sg13g2_mux2_1 _16740_ (.A0(net2330),
    .A1(\soc_inst.cpu_core.ex_instr[22] ),
    .S(net4955),
    .X(_01256_));
 sg13g2_a21oi_1 _16741_ (.A1(net4958),
    .A2(_05773_),
    .Y(_01257_),
    .B1(_09239_));
 sg13g2_mux2_1 _16742_ (.A0(net2354),
    .A1(net2362),
    .S(net4923),
    .X(_01258_));
 sg13g2_nor2_1 _16743_ (.A(net4919),
    .B(net720),
    .Y(_02610_));
 sg13g2_a21oi_1 _16744_ (.A1(net4919),
    .A2(_05775_),
    .Y(_01259_),
    .B1(_02610_));
 sg13g2_mux2_1 _16745_ (.A0(net2139),
    .A1(net2067),
    .S(net4923),
    .X(_01260_));
 sg13g2_mux2_1 _16746_ (.A0(\soc_inst.cpu_core.id_imm12[7] ),
    .A1(net2078),
    .S(net4922),
    .X(_01261_));
 sg13g2_mux2_1 _16747_ (.A0(\soc_inst.cpu_core.id_imm12[8] ),
    .A1(net2082),
    .S(net4917),
    .X(_01262_));
 sg13g2_nor2_1 _16748_ (.A(net4917),
    .B(net567),
    .Y(_02611_));
 sg13g2_a21oi_1 _16749_ (.A1(net4955),
    .A2(_05778_),
    .Y(_01263_),
    .B1(_02611_));
 sg13g2_nor2_1 _16750_ (.A(net4922),
    .B(net583),
    .Y(_02612_));
 sg13g2_a21oi_1 _16751_ (.A1(net4922),
    .A2(_05781_),
    .Y(_01264_),
    .B1(_02612_));
 sg13g2_mux2_1 _16752_ (.A0(\soc_inst.cpu_core.id_imm12[11] ),
    .A1(net2269),
    .S(net4960),
    .X(_01265_));
 sg13g2_nor2_1 _16753_ (.A(\soc_inst.cpu_core.id_int_is_interrupt ),
    .B(net4964),
    .Y(_02613_));
 sg13g2_a22oi_1 _16754_ (.Y(_01266_),
    .B1(net4661),
    .B2(_05677_),
    .A2(_05734_),
    .A1(net4938));
 sg13g2_a22oi_1 _16755_ (.Y(_01267_),
    .B1(net4661),
    .B2(_05678_),
    .A2(_05735_),
    .A1(net4972));
 sg13g2_a22oi_1 _16756_ (.Y(_01268_),
    .B1(net4661),
    .B2(_05679_),
    .A2(_05736_),
    .A1(net4972));
 sg13g2_a22oi_1 _16757_ (.Y(_01269_),
    .B1(net4661),
    .B2(_05680_),
    .A2(_05737_),
    .A1(net4972));
 sg13g2_a22oi_1 _16758_ (.Y(_01270_),
    .B1(net4661),
    .B2(_05681_),
    .A2(_05738_),
    .A1(net4972));
 sg13g2_a22oi_1 _16759_ (.Y(_01271_),
    .B1(net4661),
    .B2(_05682_),
    .A2(_05739_),
    .A1(net4938));
 sg13g2_a22oi_1 _16760_ (.Y(_01272_),
    .B1(net4661),
    .B2(_05683_),
    .A2(_05740_),
    .A1(net4938));
 sg13g2_a22oi_1 _16761_ (.Y(_01273_),
    .B1(net4662),
    .B2(_05684_),
    .A2(_05741_),
    .A1(net4966));
 sg13g2_a22oi_1 _16762_ (.Y(_01274_),
    .B1(net4662),
    .B2(_05685_),
    .A2(_05742_),
    .A1(net4961));
 sg13g2_a22oi_1 _16763_ (.Y(_01275_),
    .B1(net4662),
    .B2(_05686_),
    .A2(_05743_),
    .A1(net4963));
 sg13g2_a22oi_1 _16764_ (.Y(_01276_),
    .B1(net4661),
    .B2(_05687_),
    .A2(_05744_),
    .A1(net4938));
 sg13g2_a22oi_1 _16765_ (.Y(_01277_),
    .B1(net4662),
    .B2(_05689_),
    .A2(_05745_),
    .A1(net4962));
 sg13g2_a22oi_1 _16766_ (.Y(_01278_),
    .B1(net4662),
    .B2(_05691_),
    .A2(_05746_),
    .A1(net4960));
 sg13g2_a22oi_1 _16767_ (.Y(_01279_),
    .B1(net4663),
    .B2(_05692_),
    .A2(_05747_),
    .A1(net4964));
 sg13g2_a22oi_1 _16768_ (.Y(_01280_),
    .B1(net4662),
    .B2(_05693_),
    .A2(_05748_),
    .A1(net4960));
 sg13g2_a22oi_1 _16769_ (.Y(_01281_),
    .B1(net4663),
    .B2(_05694_),
    .A2(_05749_),
    .A1(net4955));
 sg13g2_a22oi_1 _16770_ (.Y(_01282_),
    .B1(net4660),
    .B2(_05696_),
    .A2(_05750_),
    .A1(net4954));
 sg13g2_a22oi_1 _16771_ (.Y(_01283_),
    .B1(net4660),
    .B2(_05697_),
    .A2(_05751_),
    .A1(net4954));
 sg13g2_a22oi_1 _16772_ (.Y(_01284_),
    .B1(net4660),
    .B2(_05698_),
    .A2(_05752_),
    .A1(net4954));
 sg13g2_a22oi_1 _16773_ (.Y(_01285_),
    .B1(net4660),
    .B2(_05699_),
    .A2(_05753_),
    .A1(net4952));
 sg13g2_a22oi_1 _16774_ (.Y(_01286_),
    .B1(net4660),
    .B2(_05700_),
    .A2(_05754_),
    .A1(net4954));
 sg13g2_a22oi_1 _16775_ (.Y(_01287_),
    .B1(net4660),
    .B2(_05702_),
    .A2(_05755_),
    .A1(net4952));
 sg13g2_a22oi_1 _16776_ (.Y(_01288_),
    .B1(net4660),
    .B2(_05703_),
    .A2(_05756_),
    .A1(net4957));
 sg13g2_a22oi_1 _16777_ (.Y(_01289_),
    .B1(net4660),
    .B2(_05704_),
    .A2(_05757_),
    .A1(net4954));
 sg13g2_mux2_1 _16778_ (.A0(\soc_inst.cpu_core.id_rs1_data[0] ),
    .A1(net1213),
    .S(net4978),
    .X(_01290_));
 sg13g2_mux2_1 _16779_ (.A0(net1250),
    .A1(net808),
    .S(net4907),
    .X(_01291_));
 sg13g2_mux2_1 _16780_ (.A0(\soc_inst.cpu_core.id_rs1_data[2] ),
    .A1(net801),
    .S(net4971),
    .X(_01292_));
 sg13g2_mux2_1 _16781_ (.A0(\soc_inst.cpu_core.id_rs1_data[3] ),
    .A1(net857),
    .S(net4986),
    .X(_01293_));
 sg13g2_nand2_1 _16782_ (.Y(_02614_),
    .A(net4941),
    .B(net257));
 sg13g2_o21ai_1 _16783_ (.B1(_02614_),
    .Y(_01294_),
    .A1(net4940),
    .A2(_05656_));
 sg13g2_nand2_1 _16784_ (.Y(_02615_),
    .A(net4945),
    .B(net305));
 sg13g2_o21ai_1 _16785_ (.B1(_02615_),
    .Y(_01295_),
    .A1(net4945),
    .A2(_05654_));
 sg13g2_nand2_1 _16786_ (.Y(_02616_),
    .A(net4944),
    .B(net352));
 sg13g2_o21ai_1 _16787_ (.B1(_02616_),
    .Y(_01296_),
    .A1(net4943),
    .A2(_05653_));
 sg13g2_nand2_1 _16788_ (.Y(_02617_),
    .A(net4943),
    .B(net271));
 sg13g2_o21ai_1 _16789_ (.B1(_02617_),
    .Y(_01297_),
    .A1(net4944),
    .A2(_05652_));
 sg13g2_mux2_1 _16790_ (.A0(\soc_inst.cpu_core.id_rs1_data[8] ),
    .A1(net1144),
    .S(net4935),
    .X(_01298_));
 sg13g2_mux2_1 _16791_ (.A0(\soc_inst.cpu_core.id_rs1_data[9] ),
    .A1(net2589),
    .S(net4935),
    .X(_01299_));
 sg13g2_mux2_1 _16792_ (.A0(net2550),
    .A1(net2456),
    .S(net4972),
    .X(_01300_));
 sg13g2_mux2_1 _16793_ (.A0(net764),
    .A1(net637),
    .S(net4920),
    .X(_01301_));
 sg13g2_mux2_1 _16794_ (.A0(\soc_inst.cpu_core.id_rs1_data[12] ),
    .A1(net2107),
    .S(net4920),
    .X(_01302_));
 sg13g2_mux2_1 _16795_ (.A0(\soc_inst.cpu_core.id_rs1_data[13] ),
    .A1(net780),
    .S(net4918),
    .X(_01303_));
 sg13g2_nand2_1 _16796_ (.Y(_02618_),
    .A(net4907),
    .B(net835));
 sg13g2_o21ai_1 _16797_ (.B1(_02618_),
    .Y(_01304_),
    .A1(net4907),
    .A2(_05660_));
 sg13g2_nand2_1 _16798_ (.Y(_02619_),
    .A(net4923),
    .B(net444));
 sg13g2_o21ai_1 _16799_ (.B1(_02619_),
    .Y(_01305_),
    .A1(net4919),
    .A2(_05658_));
 sg13g2_mux2_1 _16800_ (.A0(net1516),
    .A1(net1137),
    .S(net4956),
    .X(_01306_));
 sg13g2_mux2_1 _16801_ (.A0(net2339),
    .A1(net2223),
    .S(net4911),
    .X(_01307_));
 sg13g2_nand2_1 _16802_ (.Y(_02620_),
    .A(net4913),
    .B(net873));
 sg13g2_o21ai_1 _16803_ (.B1(_02620_),
    .Y(_01308_),
    .A1(net4910),
    .A2(_05676_));
 sg13g2_nand2_1 _16804_ (.Y(_02621_),
    .A(net4913),
    .B(net737));
 sg13g2_o21ai_1 _16805_ (.B1(_02621_),
    .Y(_01309_),
    .A1(net4910),
    .A2(_05674_));
 sg13g2_mux2_1 _16806_ (.A0(\soc_inst.cpu_core.id_rs1_data[20] ),
    .A1(net1314),
    .S(net4915),
    .X(_01310_));
 sg13g2_nand2_1 _16807_ (.Y(_02622_),
    .A(net4913),
    .B(net730));
 sg13g2_o21ai_1 _16808_ (.B1(_02622_),
    .Y(_01311_),
    .A1(net4910),
    .A2(_05672_));
 sg13g2_nand2_1 _16809_ (.Y(_02623_),
    .A(net4913),
    .B(net647));
 sg13g2_o21ai_1 _16810_ (.B1(_02623_),
    .Y(_01312_),
    .A1(net4910),
    .A2(_05670_));
 sg13g2_nand2_1 _16811_ (.Y(_02624_),
    .A(net4915),
    .B(net755));
 sg13g2_o21ai_1 _16812_ (.B1(_02624_),
    .Y(_01313_),
    .A1(net4915),
    .A2(_05668_));
 sg13g2_mux2_1 _16813_ (.A0(net1393),
    .A1(net1256),
    .S(net4992),
    .X(_01314_));
 sg13g2_mux2_1 _16814_ (.A0(\soc_inst.cpu_core.id_rs1_data[25] ),
    .A1(net877),
    .S(net4991),
    .X(_01315_));
 sg13g2_nand2_1 _16815_ (.Y(_02625_),
    .A(net4923),
    .B(net2264));
 sg13g2_o21ai_1 _16816_ (.B1(_02625_),
    .Y(_01316_),
    .A1(net4923),
    .A2(_05666_));
 sg13g2_mux2_1 _16817_ (.A0(net942),
    .A1(net934),
    .S(net4988),
    .X(_01317_));
 sg13g2_mux2_1 _16818_ (.A0(net1030),
    .A1(net916),
    .S(net4989),
    .X(_01318_));
 sg13g2_mux2_1 _16819_ (.A0(\soc_inst.cpu_core.id_rs1_data[29] ),
    .A1(net847),
    .S(net4990),
    .X(_01319_));
 sg13g2_nand2_1 _16820_ (.Y(_02626_),
    .A(net4912),
    .B(net2092));
 sg13g2_o21ai_1 _16821_ (.B1(_02626_),
    .Y(_01320_),
    .A1(net4912),
    .A2(_05663_));
 sg13g2_mux2_1 _16822_ (.A0(\soc_inst.cpu_core.id_rs1_data[31] ),
    .A1(net2633),
    .S(net4923),
    .X(_01321_));
 sg13g2_nor2_1 _16823_ (.A(\soc_inst.cpu_core.ex_alu_result[0] ),
    .B(net4976),
    .Y(_02627_));
 sg13g2_a21oi_1 _16824_ (.A1(net4984),
    .A2(_05483_),
    .Y(_01322_),
    .B1(_02627_));
 sg13g2_nor2_1 _16825_ (.A(net2804),
    .B(net4976),
    .Y(_02628_));
 sg13g2_a21oi_1 _16826_ (.A1(net4984),
    .A2(_05482_),
    .Y(_01323_),
    .B1(_02628_));
 sg13g2_nor2_1 _16827_ (.A(net4993),
    .B(net2751),
    .Y(_02629_));
 sg13g2_a21oi_1 _16828_ (.A1(net4993),
    .A2(_05484_),
    .Y(_01324_),
    .B1(_02629_));
 sg13g2_nor2_1 _16829_ (.A(net4993),
    .B(net2777),
    .Y(_02630_));
 sg13g2_a21oi_1 _16830_ (.A1(net4993),
    .A2(_05485_),
    .Y(_01325_),
    .B1(_02630_));
 sg13g2_nor2_1 _16831_ (.A(net4993),
    .B(net2743),
    .Y(_02631_));
 sg13g2_a21oi_1 _16832_ (.A1(net4993),
    .A2(_05487_),
    .Y(_01326_),
    .B1(_02631_));
 sg13g2_nor2_1 _16833_ (.A(net4994),
    .B(\soc_inst.cpu_core.ex_alu_result[5] ),
    .Y(_02632_));
 sg13g2_a21oi_1 _16834_ (.A1(net4994),
    .A2(_05486_),
    .Y(_01327_),
    .B1(_02632_));
 sg13g2_nor2_1 _16835_ (.A(net4994),
    .B(\soc_inst.cpu_core.ex_alu_result[6] ),
    .Y(_02633_));
 sg13g2_a21oi_1 _16836_ (.A1(net4993),
    .A2(_05488_),
    .Y(_01328_),
    .B1(_02633_));
 sg13g2_nor2_1 _16837_ (.A(net4994),
    .B(\soc_inst.cpu_core.ex_alu_result[7] ),
    .Y(_02634_));
 sg13g2_a21oi_1 _16838_ (.A1(net4994),
    .A2(_05489_),
    .Y(_01329_),
    .B1(_02634_));
 sg13g2_nor2_1 _16839_ (.A(net4984),
    .B(\soc_inst.cpu_core.ex_alu_result[8] ),
    .Y(_02635_));
 sg13g2_a21oi_1 _16840_ (.A1(_05418_),
    .A2(net4984),
    .Y(_01330_),
    .B1(_02635_));
 sg13g2_nor2_1 _16841_ (.A(net4983),
    .B(\soc_inst.cpu_core.ex_alu_result[9] ),
    .Y(_02636_));
 sg13g2_a21oi_1 _16842_ (.A1(_05419_),
    .A2(net4983),
    .Y(_01331_),
    .B1(_02636_));
 sg13g2_nor2_1 _16843_ (.A(net4975),
    .B(\soc_inst.cpu_core.ex_alu_result[10] ),
    .Y(_02637_));
 sg13g2_a21oi_1 _16844_ (.A1(_05421_),
    .A2(net4973),
    .Y(_01332_),
    .B1(_02637_));
 sg13g2_nor2_1 _16845_ (.A(net4973),
    .B(\soc_inst.cpu_core.ex_alu_result[11] ),
    .Y(_02638_));
 sg13g2_a21oi_1 _16846_ (.A1(_05420_),
    .A2(net4986),
    .Y(_01333_),
    .B1(_02638_));
 sg13g2_nor2_1 _16847_ (.A(net4988),
    .B(net2833),
    .Y(_02639_));
 sg13g2_a21oi_1 _16848_ (.A1(_05423_),
    .A2(net4993),
    .Y(_01334_),
    .B1(_02639_));
 sg13g2_nor2_1 _16849_ (.A(net4969),
    .B(net2649),
    .Y(_02640_));
 sg13g2_a21oi_1 _16850_ (.A1(_05422_),
    .A2(net4988),
    .Y(_01335_),
    .B1(_02640_));
 sg13g2_nor2_2 _16851_ (.A(net4988),
    .B(\soc_inst.cpu_core.ex_alu_result[14] ),
    .Y(_02641_));
 sg13g2_a21oi_1 _16852_ (.A1(_05425_),
    .A2(net4997),
    .Y(_01336_),
    .B1(_02641_));
 sg13g2_nor2_2 _16853_ (.A(net4967),
    .B(net2673),
    .Y(_02642_));
 sg13g2_a21oi_1 _16854_ (.A1(_05424_),
    .A2(net4983),
    .Y(_01337_),
    .B1(_02642_));
 sg13g2_nor2_1 _16855_ (.A(net4968),
    .B(net1109),
    .Y(_02643_));
 sg13g2_a21oi_1 _16856_ (.A1(_05426_),
    .A2(net4987),
    .Y(_01338_),
    .B1(_02643_));
 sg13g2_mux2_1 _16857_ (.A0(net1996),
    .A1(net2813),
    .S(net4987),
    .X(_01339_));
 sg13g2_nor2_1 _16858_ (.A(net4957),
    .B(net1128),
    .Y(_02644_));
 sg13g2_a21oi_1 _16859_ (.A1(_05428_),
    .A2(net4987),
    .Y(_01340_),
    .B1(_02644_));
 sg13g2_nor2_1 _16860_ (.A(net4957),
    .B(net898),
    .Y(_02645_));
 sg13g2_a21oi_1 _16861_ (.A1(_05427_),
    .A2(net4987),
    .Y(_01341_),
    .B1(_02645_));
 sg13g2_nor2_1 _16862_ (.A(net4959),
    .B(net736),
    .Y(_02646_));
 sg13g2_a21oi_1 _16863_ (.A1(_05430_),
    .A2(net4968),
    .Y(_01342_),
    .B1(_02646_));
 sg13g2_nor2_1 _16864_ (.A(net4959),
    .B(net2643),
    .Y(_02647_));
 sg13g2_a21oi_1 _16865_ (.A1(_05429_),
    .A2(net4967),
    .Y(_01343_),
    .B1(_02647_));
 sg13g2_nor2_1 _16866_ (.A(net4968),
    .B(net2213),
    .Y(_02648_));
 sg13g2_a21oi_1 _16867_ (.A1(_05432_),
    .A2(net4968),
    .Y(_01344_),
    .B1(_02648_));
 sg13g2_nor2_1 _16868_ (.A(net4959),
    .B(net1974),
    .Y(_02649_));
 sg13g2_a21oi_1 _16869_ (.A1(_05431_),
    .A2(net4967),
    .Y(_01345_),
    .B1(_02649_));
 sg13g2_mux2_1 _16870_ (.A0(\soc_inst.cpu_core.ex_alu_result[24] ),
    .A1(net2267),
    .S(net4980),
    .X(_01346_));
 sg13g2_mux2_1 _16871_ (.A0(\soc_inst.cpu_core.ex_alu_result[25] ),
    .A1(net2346),
    .S(net4941),
    .X(_01347_));
 sg13g2_mux2_1 _16872_ (.A0(\soc_inst.cpu_core.ex_alu_result[26] ),
    .A1(net2153),
    .S(net4980),
    .X(_01348_));
 sg13g2_mux2_1 _16873_ (.A0(\soc_inst.cpu_core.ex_alu_result[27] ),
    .A1(net2412),
    .S(net4948),
    .X(_01349_));
 sg13g2_mux2_1 _16874_ (.A0(\soc_inst.cpu_core.ex_alu_result[28] ),
    .A1(net2259),
    .S(net4958),
    .X(_01350_));
 sg13g2_nand2_1 _16875_ (.Y(_02650_),
    .A(net633),
    .B(net4955));
 sg13g2_o21ai_1 _16876_ (.B1(_02650_),
    .Y(_01351_),
    .A1(net4955),
    .A2(_05779_));
 sg13g2_nor2_1 _16877_ (.A(net4971),
    .B(\soc_inst.cpu_core.ex_alu_result[30] ),
    .Y(_02651_));
 sg13g2_a21oi_1 _16878_ (.A1(_05434_),
    .A2(net4973),
    .Y(_01352_),
    .B1(_02651_));
 sg13g2_mux2_1 _16879_ (.A0(\soc_inst.cpu_core.ex_alu_result[31] ),
    .A1(net2254),
    .S(net4963),
    .X(_01353_));
 sg13g2_nand2_1 _16880_ (.Y(_02652_),
    .A(net4978),
    .B(net336));
 sg13g2_o21ai_1 _16881_ (.B1(_02652_),
    .Y(_01354_),
    .A1(net4948),
    .A2(_05651_));
 sg13g2_mux2_1 _16882_ (.A0(net1057),
    .A1(net896),
    .S(net4950),
    .X(_01355_));
 sg13g2_mux2_1 _16883_ (.A0(net1404),
    .A1(net1265),
    .S(net4947),
    .X(_01356_));
 sg13g2_mux2_1 _16884_ (.A0(net875),
    .A1(net783),
    .S(net4946),
    .X(_01357_));
 sg13g2_nand2_1 _16885_ (.Y(_02653_),
    .A(net4946),
    .B(net399));
 sg13g2_o21ai_1 _16886_ (.B1(_02653_),
    .Y(_01358_),
    .A1(net4946),
    .A2(_05657_));
 sg13g2_nand2_1 _16887_ (.Y(_02654_),
    .A(net4946),
    .B(net364));
 sg13g2_o21ai_1 _16888_ (.B1(_02654_),
    .Y(_01359_),
    .A1(net4946),
    .A2(_05655_));
 sg13g2_mux2_1 _16889_ (.A0(net1261),
    .A1(net1147),
    .S(net4947),
    .X(_01360_));
 sg13g2_mux2_1 _16890_ (.A0(net1606),
    .A1(net1201),
    .S(net4944),
    .X(_01361_));
 sg13g2_nand2_1 _16891_ (.Y(_02655_),
    .A(net4945),
    .B(net707));
 sg13g2_o21ai_1 _16892_ (.B1(_02655_),
    .Y(_01362_),
    .A1(net4945),
    .A2(_05662_));
 sg13g2_mux2_1 _16893_ (.A0(\soc_inst.cpu_core.id_rs2_data[9] ),
    .A1(net940),
    .S(net4978),
    .X(_01363_));
 sg13g2_nand2_1 _16894_ (.Y(_02656_),
    .A(net4979),
    .B(net717));
 sg13g2_o21ai_1 _16895_ (.B1(_02656_),
    .Y(_01364_),
    .A1(net4978),
    .A2(_05661_));
 sg13g2_mux2_1 _16896_ (.A0(\soc_inst.cpu_core.id_rs2_data[11] ),
    .A1(net1476),
    .S(net4978),
    .X(_01365_));
 sg13g2_mux2_1 _16897_ (.A0(net1373),
    .A1(net1102),
    .S(net4978),
    .X(_01366_));
 sg13g2_mux2_1 _16898_ (.A0(net2257),
    .A1(net2162),
    .S(net4918),
    .X(_01367_));
 sg13g2_mux2_1 _16899_ (.A0(net1334),
    .A1(net1293),
    .S(net4924),
    .X(_01368_));
 sg13g2_nand2_1 _16900_ (.Y(_02657_),
    .A(net4947),
    .B(net372));
 sg13g2_o21ai_1 _16901_ (.B1(_02657_),
    .Y(_01369_),
    .A1(net4946),
    .A2(_05659_));
 sg13g2_mux2_1 _16902_ (.A0(net1283),
    .A1(net1066),
    .S(net4990),
    .X(_01370_));
 sg13g2_mux2_1 _16903_ (.A0(net2444),
    .A1(\soc_inst.cpu_core.ex_rs2_data[17] ),
    .S(net4913),
    .X(_01371_));
 sg13g2_mux2_1 _16904_ (.A0(\soc_inst.cpu_core.id_rs2_data[18] ),
    .A1(net1085),
    .S(net4989),
    .X(_01372_));
 sg13g2_nand2_1 _16905_ (.Y(_02658_),
    .A(net4995),
    .B(net311));
 sg13g2_o21ai_1 _16906_ (.B1(_02658_),
    .Y(_01373_),
    .A1(net4996),
    .A2(_05675_));
 sg13g2_nand2_1 _16907_ (.Y(_02659_),
    .A(net4915),
    .B(\soc_inst.cpu_core.ex_rs2_data[20] ));
 sg13g2_o21ai_1 _16908_ (.B1(_02659_),
    .Y(_01374_),
    .A1(net4915),
    .A2(_05673_));
 sg13g2_mux2_1 _16909_ (.A0(net1282),
    .A1(net1174),
    .S(net4989),
    .X(_01375_));
 sg13g2_nand2_1 _16910_ (.Y(_02660_),
    .A(net4932),
    .B(\soc_inst.cpu_core.ex_rs2_data[22] ));
 sg13g2_o21ai_1 _16911_ (.B1(_02660_),
    .Y(_01376_),
    .A1(net4932),
    .A2(_05671_));
 sg13g2_nand2_1 _16912_ (.Y(_02661_),
    .A(net4957),
    .B(net1972));
 sg13g2_o21ai_1 _16913_ (.B1(_02661_),
    .Y(_01377_),
    .A1(net4957),
    .A2(_05669_));
 sg13g2_nand2_1 _16914_ (.Y(_02662_),
    .A(net4946),
    .B(net497));
 sg13g2_o21ai_1 _16915_ (.B1(_02662_),
    .Y(_01378_),
    .A1(net4944),
    .A2(_05667_));
 sg13g2_mux2_1 _16916_ (.A0(net1248),
    .A1(net1172),
    .S(net4980),
    .X(_01379_));
 sg13g2_mux2_1 _16917_ (.A0(net2787),
    .A1(net2397),
    .S(net4936),
    .X(_01380_));
 sg13g2_nand2_1 _16918_ (.Y(_02663_),
    .A(net4995),
    .B(net316));
 sg13g2_o21ai_1 _16919_ (.B1(_02663_),
    .Y(_01381_),
    .A1(net4994),
    .A2(_05665_));
 sg13g2_nand2_1 _16920_ (.Y(_02664_),
    .A(net4981),
    .B(net1874));
 sg13g2_o21ai_1 _16921_ (.B1(_02664_),
    .Y(_01382_),
    .A1(net4980),
    .A2(_05664_));
 sg13g2_mux2_1 _16922_ (.A0(net1607),
    .A1(net713),
    .S(net4936),
    .X(_01383_));
 sg13g2_mux2_1 _16923_ (.A0(net2756),
    .A1(net2466),
    .S(net4940),
    .X(_01384_));
 sg13g2_mux2_1 _16924_ (.A0(\soc_inst.cpu_core.id_rs2_data[31] ),
    .A1(net863),
    .S(net4996),
    .X(_01385_));
 sg13g2_nor2_2 _16925_ (.A(net2745),
    .B(net2349),
    .Y(_02665_));
 sg13g2_nor3_1 _16926_ (.A(\soc_inst.cpu_core.alu.op[0] ),
    .B(\soc_inst.cpu_core.alu.op[1] ),
    .C(\soc_inst.cpu_core.alu.op[2] ),
    .Y(_02666_));
 sg13g2_nor2b_2 _16927_ (.A(\soc_inst.cpu_core.alu.op[1] ),
    .B_N(\soc_inst.cpu_core.alu.op[0] ),
    .Y(_02667_));
 sg13g2_and2_1 _16928_ (.A(\soc_inst.cpu_core.alu.op[2] ),
    .B(_02667_),
    .X(_02668_));
 sg13g2_nand2_2 _16929_ (.Y(_02669_),
    .A(\soc_inst.cpu_core.alu.op[2] ),
    .B(_02667_));
 sg13g2_and2_1 _16930_ (.A(net4865),
    .B(_02666_),
    .X(_02670_));
 sg13g2_nand2_2 _16931_ (.Y(_02671_),
    .A(net2747),
    .B(_02666_));
 sg13g2_nand3_1 _16932_ (.B(_02669_),
    .C(net4444),
    .A(net4865),
    .Y(_02672_));
 sg13g2_and2_1 _16933_ (.A(net4741),
    .B(_02672_),
    .X(_02673_));
 sg13g2_nand2_1 _16934_ (.Y(_02674_),
    .A(net4741),
    .B(_02672_));
 sg13g2_nand2b_1 _16935_ (.Y(_02675_),
    .B(net4854),
    .A_N(\soc_inst.cpu_core.alu.b[31] ));
 sg13g2_xor2_1 _16936_ (.B(net4854),
    .A(\soc_inst.cpu_core.alu.b[31] ),
    .X(_02676_));
 sg13g2_nand2_1 _16937_ (.Y(_02677_),
    .A(_05809_),
    .B(_05810_));
 sg13g2_nor2_1 _16938_ (.A(_05809_),
    .B(_05810_),
    .Y(_02678_));
 sg13g2_xor2_1 _16939_ (.B(\soc_inst.cpu_core.alu.a[15] ),
    .A(\soc_inst.cpu_core.alu.b[15] ),
    .X(_02679_));
 sg13g2_xnor2_1 _16940_ (.Y(_02680_),
    .A(\soc_inst.cpu_core.alu.b[15] ),
    .B(\soc_inst.cpu_core.alu.a[15] ));
 sg13g2_nor2_2 _16941_ (.A(_05811_),
    .B(_05812_),
    .Y(_02681_));
 sg13g2_nand2_1 _16942_ (.Y(_02682_),
    .A(_05811_),
    .B(_05812_));
 sg13g2_nor2b_2 _16943_ (.A(_02681_),
    .B_N(_02682_),
    .Y(_02683_));
 sg13g2_nand2b_2 _16944_ (.Y(_02684_),
    .B(_02682_),
    .A_N(_02681_));
 sg13g2_nand2_1 _16945_ (.Y(_02685_),
    .A(_05811_),
    .B(\soc_inst.cpu_core.alu.a[14] ));
 sg13g2_xor2_1 _16946_ (.B(net4863),
    .A(\soc_inst.cpu_core.alu.b[13] ),
    .X(_02686_));
 sg13g2_xnor2_1 _16947_ (.Y(_02687_),
    .A(\soc_inst.cpu_core.alu.b[13] ),
    .B(net4863));
 sg13g2_nor2_1 _16948_ (.A(\soc_inst.cpu_core.alu.b[11] ),
    .B(\soc_inst.cpu_core.alu.a[11] ),
    .Y(_02688_));
 sg13g2_inv_1 _16949_ (.Y(_02689_),
    .A(_02688_));
 sg13g2_nand2_2 _16950_ (.Y(_02690_),
    .A(\soc_inst.cpu_core.alu.b[11] ),
    .B(\soc_inst.cpu_core.alu.a[11] ));
 sg13g2_nor2b_2 _16951_ (.A(_02688_),
    .B_N(_02690_),
    .Y(_02691_));
 sg13g2_nor2_1 _16952_ (.A(\soc_inst.cpu_core.alu.b[10] ),
    .B(\soc_inst.cpu_core.alu.a[10] ),
    .Y(_02692_));
 sg13g2_nand2_1 _16953_ (.Y(_02693_),
    .A(_05819_),
    .B(_05820_));
 sg13g2_nand2_2 _16954_ (.Y(_02694_),
    .A(net1960),
    .B(net2719));
 sg13g2_and2_1 _16955_ (.A(_02693_),
    .B(_02694_),
    .X(_02695_));
 sg13g2_nand2_1 _16956_ (.Y(_02696_),
    .A(_02693_),
    .B(_02694_));
 sg13g2_nor2_1 _16957_ (.A(_02691_),
    .B(_02695_),
    .Y(_02697_));
 sg13g2_nand2_1 _16958_ (.Y(_02698_),
    .A(_05821_),
    .B(_05822_));
 sg13g2_nand2_2 _16959_ (.Y(_02699_),
    .A(\soc_inst.cpu_core.alu.b[9] ),
    .B(\soc_inst.cpu_core.alu.a[9] ));
 sg13g2_and2_1 _16960_ (.A(_02698_),
    .B(_02699_),
    .X(_02700_));
 sg13g2_nand2_2 _16961_ (.Y(_02701_),
    .A(_02698_),
    .B(_02699_));
 sg13g2_nand2_1 _16962_ (.Y(_02702_),
    .A(_05823_),
    .B(\soc_inst.cpu_core.alu.a[8] ));
 sg13g2_nand2b_1 _16963_ (.Y(_02703_),
    .B(_02701_),
    .A_N(_02702_));
 sg13g2_o21ai_1 _16964_ (.B1(_02703_),
    .Y(_02704_),
    .A1(\soc_inst.cpu_core.alu.b[9] ),
    .A2(_05822_));
 sg13g2_nand2_1 _16965_ (.Y(_02705_),
    .A(_05825_),
    .B(\soc_inst.cpu_core.alu.a[7] ));
 sg13g2_or2_1 _16966_ (.X(_02706_),
    .B(\soc_inst.cpu_core.alu.a[7] ),
    .A(\soc_inst.cpu_core.alu.b[7] ));
 sg13g2_nand2_1 _16967_ (.Y(_02707_),
    .A(\soc_inst.cpu_core.alu.b[7] ),
    .B(\soc_inst.cpu_core.alu.a[7] ));
 sg13g2_inv_1 _16968_ (.Y(_02708_),
    .A(_02707_));
 sg13g2_and2_1 _16969_ (.A(_02706_),
    .B(_02707_),
    .X(_02709_));
 sg13g2_nor2_1 _16970_ (.A(\soc_inst.cpu_core.alu.b[6] ),
    .B(_05828_),
    .Y(_02710_));
 sg13g2_nand2_1 _16971_ (.Y(_02711_),
    .A(_05827_),
    .B(_05828_));
 sg13g2_nand2_1 _16972_ (.Y(_02712_),
    .A(\soc_inst.cpu_core.alu.b[6] ),
    .B(\soc_inst.cpu_core.alu.a[6] ));
 sg13g2_inv_1 _16973_ (.Y(_02713_),
    .A(_02712_));
 sg13g2_and2_1 _16974_ (.A(_02711_),
    .B(_02712_),
    .X(_02714_));
 sg13g2_nand2_1 _16975_ (.Y(_02715_),
    .A(_02711_),
    .B(_02712_));
 sg13g2_nand2_1 _16976_ (.Y(_02716_),
    .A(_05829_),
    .B(\soc_inst.cpu_core.alu.a[5] ));
 sg13g2_nand2_1 _16977_ (.Y(_02717_),
    .A(_05829_),
    .B(_05830_));
 sg13g2_nand2_1 _16978_ (.Y(_02718_),
    .A(\soc_inst.cpu_core.alu.b[5] ),
    .B(\soc_inst.cpu_core.alu.a[5] ));
 sg13g2_and2_1 _16979_ (.A(_02717_),
    .B(_02718_),
    .X(_02719_));
 sg13g2_nand2_1 _16980_ (.Y(_02720_),
    .A(_02717_),
    .B(_02718_));
 sg13g2_nand2_1 _16981_ (.Y(_02721_),
    .A(net4737),
    .B(\soc_inst.cpu_core.alu.a[4] ));
 sg13g2_inv_1 _16982_ (.Y(_02722_),
    .A(_02721_));
 sg13g2_nand2_1 _16983_ (.Y(_02723_),
    .A(net4737),
    .B(_05832_));
 sg13g2_nor2_2 _16984_ (.A(net4737),
    .B(_05832_),
    .Y(_02724_));
 sg13g2_xnor2_1 _16985_ (.Y(_02725_),
    .A(net4806),
    .B(\soc_inst.cpu_core.alu.a[4] ));
 sg13g2_nand2_1 _16986_ (.Y(_02726_),
    .A(net4733),
    .B(\soc_inst.cpu_core.alu.a[3] ));
 sg13g2_and2_1 _16987_ (.A(net4814),
    .B(\soc_inst.cpu_core.alu.a[3] ),
    .X(_02727_));
 sg13g2_nand2_1 _16988_ (.Y(_02728_),
    .A(net4816),
    .B(\soc_inst.cpu_core.alu.a[3] ));
 sg13g2_nor2_1 _16989_ (.A(net4816),
    .B(\soc_inst.cpu_core.alu.a[3] ),
    .Y(_02729_));
 sg13g2_nor2_2 _16990_ (.A(_02727_),
    .B(_02729_),
    .Y(_02730_));
 sg13g2_nor2b_1 _16991_ (.A(net4823),
    .B_N(net4864),
    .Y(_02731_));
 sg13g2_and2_1 _16992_ (.A(net4823),
    .B(net4864),
    .X(_02732_));
 sg13g2_xor2_1 _16993_ (.B(net4864),
    .A(net4822),
    .X(_02733_));
 sg13g2_xnor2_1 _16994_ (.Y(_02734_),
    .A(net4823),
    .B(net4864));
 sg13g2_nor2b_1 _16995_ (.A(net4837),
    .B_N(\soc_inst.cpu_core.alu.a[1] ),
    .Y(_02735_));
 sg13g2_nand2_1 _16996_ (.Y(_02736_),
    .A(net4837),
    .B(\soc_inst.cpu_core.alu.a[1] ));
 sg13g2_xnor2_1 _16997_ (.Y(_02737_),
    .A(net4837),
    .B(\soc_inst.cpu_core.alu.a[1] ));
 sg13g2_nand2b_1 _16998_ (.Y(_02738_),
    .B(net4848),
    .A_N(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_a21o_1 _16999_ (.A2(_02738_),
    .A1(_02737_),
    .B1(_02735_),
    .X(_02739_));
 sg13g2_a21oi_1 _17000_ (.A1(_02734_),
    .A2(_02739_),
    .Y(_02740_),
    .B1(_02731_));
 sg13g2_o21ai_1 _17001_ (.B1(_02726_),
    .Y(_02741_),
    .A1(_02730_),
    .A2(_02740_));
 sg13g2_a21oi_2 _17002_ (.B1(_02722_),
    .Y(_02742_),
    .A2(_02741_),
    .A1(_02725_));
 sg13g2_o21ai_1 _17003_ (.B1(_02716_),
    .Y(_02743_),
    .A1(_02719_),
    .A2(_02742_));
 sg13g2_a21oi_1 _17004_ (.A1(_02715_),
    .A2(_02743_),
    .Y(_02744_),
    .B1(_02710_));
 sg13g2_o21ai_1 _17005_ (.B1(_02705_),
    .Y(_02745_),
    .A1(_02709_),
    .A2(_02744_));
 sg13g2_nand2_1 _17006_ (.Y(_02746_),
    .A(_05823_),
    .B(_05824_));
 sg13g2_nand2_2 _17007_ (.Y(_02747_),
    .A(net2474),
    .B(net2380));
 sg13g2_and2_1 _17008_ (.A(_02746_),
    .B(_02747_),
    .X(_02748_));
 sg13g2_nand2_2 _17009_ (.Y(_02749_),
    .A(_02746_),
    .B(_02747_));
 sg13g2_nand2_1 _17010_ (.Y(_02750_),
    .A(_02745_),
    .B(_02749_));
 sg13g2_inv_1 _17011_ (.Y(_02751_),
    .A(_02750_));
 sg13g2_nand2_1 _17012_ (.Y(_02752_),
    .A(_02701_),
    .B(_02751_));
 sg13g2_a21oi_1 _17013_ (.A1(_02701_),
    .A2(_02751_),
    .Y(_02753_),
    .B1(_02704_));
 sg13g2_nand2_1 _17014_ (.Y(_02754_),
    .A(_05817_),
    .B(\soc_inst.cpu_core.alu.a[11] ));
 sg13g2_nor2_1 _17015_ (.A(\soc_inst.cpu_core.alu.b[10] ),
    .B(_05820_),
    .Y(_02755_));
 sg13g2_a21oi_1 _17016_ (.A1(_02696_),
    .A2(_02704_),
    .Y(_02756_),
    .B1(_02755_));
 sg13g2_or2_1 _17017_ (.X(_02757_),
    .B(_02756_),
    .A(_02691_));
 sg13g2_nand4_1 _17018_ (.B(_02701_),
    .C(_02745_),
    .A(_02697_),
    .Y(_02758_),
    .D(_02749_));
 sg13g2_nand3_1 _17019_ (.B(_02757_),
    .C(_02758_),
    .A(_02754_),
    .Y(_02759_));
 sg13g2_nand2_1 _17020_ (.Y(_02760_),
    .A(net1895),
    .B(\soc_inst.cpu_core.alu.a[12] ));
 sg13g2_xnor2_1 _17021_ (.Y(_02761_),
    .A(\soc_inst.cpu_core.alu.b[12] ),
    .B(\soc_inst.cpu_core.alu.a[12] ));
 sg13g2_nand2_1 _17022_ (.Y(_02762_),
    .A(_02759_),
    .B(_02761_));
 sg13g2_nand3_1 _17023_ (.B(_02759_),
    .C(_02761_),
    .A(_02687_),
    .Y(_02763_));
 sg13g2_nand2_1 _17024_ (.Y(_02764_),
    .A(_05815_),
    .B(\soc_inst.cpu_core.alu.a[12] ));
 sg13g2_nor2_1 _17025_ (.A(_02686_),
    .B(_02764_),
    .Y(_02765_));
 sg13g2_nand2b_1 _17026_ (.Y(_02766_),
    .B(_02687_),
    .A_N(_02764_));
 sg13g2_a21oi_1 _17027_ (.A1(_05813_),
    .A2(net4863),
    .Y(_02767_),
    .B1(_02765_));
 sg13g2_o21ai_1 _17028_ (.B1(_02685_),
    .Y(_02768_),
    .A1(_02683_),
    .A2(_02767_));
 sg13g2_and2_1 _17029_ (.A(_02680_),
    .B(_02768_),
    .X(_02769_));
 sg13g2_and4_1 _17030_ (.A(_02680_),
    .B(_02684_),
    .C(_02687_),
    .D(_02761_),
    .X(_02770_));
 sg13g2_a221oi_1 _17031_ (.B2(_02770_),
    .C1(_02769_),
    .B1(_02759_),
    .A1(_05809_),
    .Y(_02771_),
    .A2(\soc_inst.cpu_core.alu.a[15] ));
 sg13g2_nand2_2 _17032_ (.Y(_02772_),
    .A(_05805_),
    .B(_05806_));
 sg13g2_nand2_1 _17033_ (.Y(_02773_),
    .A(\soc_inst.cpu_core.alu.b[17] ),
    .B(\soc_inst.cpu_core.alu.a[17] ));
 sg13g2_and2_1 _17034_ (.A(_02772_),
    .B(_02773_),
    .X(_02774_));
 sg13g2_nor2_2 _17035_ (.A(\soc_inst.cpu_core.alu.b[16] ),
    .B(\soc_inst.cpu_core.alu.a[16] ),
    .Y(_02775_));
 sg13g2_nand2_2 _17036_ (.Y(_02776_),
    .A(\soc_inst.cpu_core.alu.b[16] ),
    .B(\soc_inst.cpu_core.alu.a[16] ));
 sg13g2_nor2b_2 _17037_ (.A(_02775_),
    .B_N(_02776_),
    .Y(_02777_));
 sg13g2_nor3_1 _17038_ (.A(_02771_),
    .B(net4215),
    .C(net4443),
    .Y(_02778_));
 sg13g2_nor2_1 _17039_ (.A(\soc_inst.cpu_core.alu.b[23] ),
    .B(net4859),
    .Y(_02779_));
 sg13g2_nand2_2 _17040_ (.Y(_02780_),
    .A(\soc_inst.cpu_core.alu.b[23] ),
    .B(net4859));
 sg13g2_nor2b_1 _17041_ (.A(_02779_),
    .B_N(_02780_),
    .Y(_02781_));
 sg13g2_nand2b_1 _17042_ (.Y(_02782_),
    .B(_02780_),
    .A_N(_02779_));
 sg13g2_nand2_1 _17043_ (.Y(_02783_),
    .A(\soc_inst.cpu_core.alu.b[22] ),
    .B(\soc_inst.cpu_core.alu.a[22] ));
 sg13g2_xnor2_1 _17044_ (.Y(_02784_),
    .A(\soc_inst.cpu_core.alu.b[22] ),
    .B(\soc_inst.cpu_core.alu.a[22] ));
 sg13g2_inv_2 _17045_ (.Y(_02785_),
    .A(_02784_));
 sg13g2_nor2_1 _17046_ (.A(_02781_),
    .B(_02785_),
    .Y(_02786_));
 sg13g2_nor2_2 _17047_ (.A(\soc_inst.cpu_core.alu.b[21] ),
    .B(\soc_inst.cpu_core.alu.a[21] ),
    .Y(_02787_));
 sg13g2_nand2_2 _17048_ (.Y(_02788_),
    .A(\soc_inst.cpu_core.alu.b[21] ),
    .B(\soc_inst.cpu_core.alu.a[21] ));
 sg13g2_nor2b_2 _17049_ (.A(_02787_),
    .B_N(_02788_),
    .Y(_02789_));
 sg13g2_nand2b_2 _17050_ (.Y(_02790_),
    .B(_02788_),
    .A_N(_02787_));
 sg13g2_nand2_2 _17051_ (.Y(_02791_),
    .A(\soc_inst.cpu_core.alu.b[20] ),
    .B(net4860));
 sg13g2_xor2_1 _17052_ (.B(net4860),
    .A(\soc_inst.cpu_core.alu.b[20] ),
    .X(_02792_));
 sg13g2_xnor2_1 _17053_ (.Y(_02793_),
    .A(\soc_inst.cpu_core.alu.b[20] ),
    .B(net4860));
 sg13g2_nor2_1 _17054_ (.A(\soc_inst.cpu_core.alu.b[19] ),
    .B(net4861),
    .Y(_02794_));
 sg13g2_xor2_1 _17055_ (.B(net4861),
    .A(\soc_inst.cpu_core.alu.b[19] ),
    .X(_02795_));
 sg13g2_xnor2_1 _17056_ (.Y(_02796_),
    .A(\soc_inst.cpu_core.alu.b[19] ),
    .B(net4861));
 sg13g2_nand2_2 _17057_ (.Y(_02797_),
    .A(\soc_inst.cpu_core.alu.b[18] ),
    .B(net4862));
 sg13g2_xor2_1 _17058_ (.B(net4862),
    .A(\soc_inst.cpu_core.alu.b[18] ),
    .X(_02798_));
 sg13g2_xnor2_1 _17059_ (.Y(_02799_),
    .A(\soc_inst.cpu_core.alu.b[18] ),
    .B(net4862));
 sg13g2_nand2_1 _17060_ (.Y(_02800_),
    .A(_02796_),
    .B(_02799_));
 sg13g2_nor3_1 _17061_ (.A(net4215),
    .B(net4443),
    .C(_02800_),
    .Y(_02801_));
 sg13g2_nand4_1 _17062_ (.B(_02790_),
    .C(_02793_),
    .A(_02786_),
    .Y(_02802_),
    .D(_02801_));
 sg13g2_nor2_1 _17063_ (.A(\soc_inst.cpu_core.alu.b[22] ),
    .B(_05796_),
    .Y(_02803_));
 sg13g2_and2_1 _17064_ (.A(_02782_),
    .B(_02803_),
    .X(_02804_));
 sg13g2_nand2_1 _17065_ (.Y(_02805_),
    .A(_05797_),
    .B(\soc_inst.cpu_core.alu.a[21] ));
 sg13g2_nand2_1 _17066_ (.Y(_02806_),
    .A(_05799_),
    .B(\soc_inst.cpu_core.alu.a[20] ));
 sg13g2_nor2b_1 _17067_ (.A(\soc_inst.cpu_core.alu.b[18] ),
    .B_N(\soc_inst.cpu_core.alu.a[18] ),
    .Y(_02807_));
 sg13g2_nand2_1 _17068_ (.Y(_02808_),
    .A(_05807_),
    .B(\soc_inst.cpu_core.alu.a[16] ));
 sg13g2_nand2_1 _17069_ (.Y(_02809_),
    .A(_05805_),
    .B(\soc_inst.cpu_core.alu.a[17] ));
 sg13g2_o21ai_1 _17070_ (.B1(_02809_),
    .Y(_02810_),
    .A1(net4215),
    .A2(_02808_));
 sg13g2_a21oi_1 _17071_ (.A1(_02799_),
    .A2(_02810_),
    .Y(_02811_),
    .B1(_02807_));
 sg13g2_nor2_1 _17072_ (.A(_02795_),
    .B(_02811_),
    .Y(_02812_));
 sg13g2_a21oi_1 _17073_ (.A1(_05801_),
    .A2(net4861),
    .Y(_02813_),
    .B1(_02812_));
 sg13g2_inv_1 _17074_ (.Y(_02814_),
    .A(_02813_));
 sg13g2_o21ai_1 _17075_ (.B1(_02806_),
    .Y(_02815_),
    .A1(_02792_),
    .A2(_02813_));
 sg13g2_nand2_1 _17076_ (.Y(_02816_),
    .A(_02790_),
    .B(_02815_));
 sg13g2_nand2_1 _17077_ (.Y(_02817_),
    .A(_02805_),
    .B(_02816_));
 sg13g2_a221oi_1 _17078_ (.B2(_02817_),
    .C1(_02804_),
    .B1(_02786_),
    .A1(_05793_),
    .Y(_02818_),
    .A2(net4859));
 sg13g2_o21ai_1 _17079_ (.B1(_02818_),
    .Y(_02819_),
    .A1(_02771_),
    .A2(_02802_));
 sg13g2_xor2_1 _17080_ (.B(net4856),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .X(_02820_));
 sg13g2_xnor2_1 _17081_ (.Y(_02821_),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .B(net4857));
 sg13g2_nor2_1 _17082_ (.A(\soc_inst.cpu_core.alu.b[27] ),
    .B(\soc_inst.cpu_core.alu.a[27] ),
    .Y(_02822_));
 sg13g2_inv_1 _17083_ (.Y(_02823_),
    .A(_02822_));
 sg13g2_nand2_1 _17084_ (.Y(_02824_),
    .A(\soc_inst.cpu_core.alu.b[27] ),
    .B(\soc_inst.cpu_core.alu.a[27] ));
 sg13g2_nor2b_2 _17085_ (.A(_02822_),
    .B_N(_02824_),
    .Y(_02825_));
 sg13g2_inv_1 _17086_ (.Y(_02826_),
    .A(_02825_));
 sg13g2_nor2_2 _17087_ (.A(\soc_inst.cpu_core.alu.b[25] ),
    .B(net4858),
    .Y(_02827_));
 sg13g2_inv_1 _17088_ (.Y(_02828_),
    .A(_02827_));
 sg13g2_nand2_2 _17089_ (.Y(_02829_),
    .A(\soc_inst.cpu_core.alu.b[25] ),
    .B(net4858));
 sg13g2_nor2b_2 _17090_ (.A(_02827_),
    .B_N(_02829_),
    .Y(_02830_));
 sg13g2_nand2_2 _17091_ (.Y(_02831_),
    .A(\soc_inst.cpu_core.alu.b[24] ),
    .B(\soc_inst.cpu_core.alu.a[24] ));
 sg13g2_inv_2 _17092_ (.Y(_02832_),
    .A(_02831_));
 sg13g2_or2_1 _17093_ (.X(_02833_),
    .B(\soc_inst.cpu_core.alu.a[24] ),
    .A(\soc_inst.cpu_core.alu.b[24] ));
 sg13g2_and2_1 _17094_ (.A(_02831_),
    .B(_02833_),
    .X(_02834_));
 sg13g2_nand2_2 _17095_ (.Y(_02835_),
    .A(_02831_),
    .B(_02833_));
 sg13g2_nor4_1 _17096_ (.A(_02820_),
    .B(_02825_),
    .C(net4442),
    .D(_02834_),
    .Y(_02836_));
 sg13g2_nand2_1 _17097_ (.Y(_02837_),
    .A(_05792_),
    .B(\soc_inst.cpu_core.alu.a[24] ));
 sg13g2_nor2_1 _17098_ (.A(net4442),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_a21oi_1 _17099_ (.A1(_05791_),
    .A2(net4858),
    .Y(_02839_),
    .B1(_02838_));
 sg13g2_nor2b_1 _17100_ (.A(\soc_inst.cpu_core.alu.b[26] ),
    .B_N(net4857),
    .Y(_02840_));
 sg13g2_nor2_1 _17101_ (.A(_02820_),
    .B(_02839_),
    .Y(_02841_));
 sg13g2_nor2_1 _17102_ (.A(_02840_),
    .B(_02841_),
    .Y(_02842_));
 sg13g2_nor2_1 _17103_ (.A(_02825_),
    .B(_02842_),
    .Y(_02843_));
 sg13g2_a221oi_1 _17104_ (.B2(_02836_),
    .C1(_02843_),
    .B1(_02819_),
    .A1(_05789_),
    .Y(_02844_),
    .A2(\soc_inst.cpu_core.alu.a[27] ));
 sg13g2_nand2_1 _17105_ (.Y(_02845_),
    .A(\soc_inst.cpu_core.alu.b[29] ),
    .B(\soc_inst.cpu_core.alu.a[29] ));
 sg13g2_xnor2_1 _17106_ (.Y(_02846_),
    .A(\soc_inst.cpu_core.alu.b[29] ),
    .B(\soc_inst.cpu_core.alu.a[29] ));
 sg13g2_nand2_1 _17107_ (.Y(_02847_),
    .A(\soc_inst.cpu_core.alu.b[28] ),
    .B(net4855));
 sg13g2_xor2_1 _17108_ (.B(net4855),
    .A(\soc_inst.cpu_core.alu.b[28] ),
    .X(_02848_));
 sg13g2_xnor2_1 _17109_ (.Y(_02849_),
    .A(\soc_inst.cpu_core.alu.b[28] ),
    .B(net4855));
 sg13g2_nand2_1 _17110_ (.Y(_02850_),
    .A(_02846_),
    .B(_02849_));
 sg13g2_nor2_1 _17111_ (.A(_02844_),
    .B(_02850_),
    .Y(_02851_));
 sg13g2_nor2b_1 _17112_ (.A(\soc_inst.cpu_core.alu.b[28] ),
    .B_N(net4855),
    .Y(_02852_));
 sg13g2_and2_1 _17113_ (.A(_02846_),
    .B(_02852_),
    .X(_02853_));
 sg13g2_a21oi_1 _17114_ (.A1(_05787_),
    .A2(\soc_inst.cpu_core.alu.a[29] ),
    .Y(_02854_),
    .B1(_02853_));
 sg13g2_o21ai_1 _17115_ (.B1(_02854_),
    .Y(_02855_),
    .A1(_02844_),
    .A2(_02850_));
 sg13g2_and2_1 _17116_ (.A(\soc_inst.cpu_core.alu.b[30] ),
    .B(\soc_inst.cpu_core.alu.a[30] ),
    .X(_02856_));
 sg13g2_xnor2_1 _17117_ (.Y(_02857_),
    .A(\soc_inst.cpu_core.alu.b[30] ),
    .B(\soc_inst.cpu_core.alu.a[30] ));
 sg13g2_and2_1 _17118_ (.A(_02855_),
    .B(_02857_),
    .X(_02858_));
 sg13g2_nor2b_1 _17119_ (.A(\soc_inst.cpu_core.alu.b[30] ),
    .B_N(\soc_inst.cpu_core.alu.a[30] ),
    .Y(_02859_));
 sg13g2_a21oi_2 _17120_ (.B1(_02859_),
    .Y(_02860_),
    .A2(_02857_),
    .A1(_02855_));
 sg13g2_nand2b_1 _17121_ (.Y(_02861_),
    .B(_02860_),
    .A_N(_02676_));
 sg13g2_nor2_2 _17122_ (.A(\soc_inst.cpu_core.alu.op[2] ),
    .B(net4865),
    .Y(_02862_));
 sg13g2_nor2b_2 _17123_ (.A(net2745),
    .B_N(\soc_inst.cpu_core.alu.op[1] ),
    .Y(_02863_));
 sg13g2_nand2_1 _17124_ (.Y(_02864_),
    .A(_02862_),
    .B(_02863_));
 sg13g2_a21oi_1 _17125_ (.A1(_02675_),
    .A2(_02861_),
    .Y(_02865_),
    .B1(_02864_));
 sg13g2_nand2_1 _17126_ (.Y(_02866_),
    .A(\soc_inst.cpu_core.alu.op[0] ),
    .B(\soc_inst.cpu_core.alu.op[1] ));
 sg13g2_and4_1 _17127_ (.A(\soc_inst.cpu_core.alu.op[0] ),
    .B(\soc_inst.cpu_core.alu.op[1] ),
    .C(_02675_),
    .D(_02862_),
    .X(_02867_));
 sg13g2_o21ai_1 _17128_ (.B1(_02867_),
    .Y(_02868_),
    .A1(_02676_),
    .A2(_02860_));
 sg13g2_nand2_1 _17129_ (.Y(_02869_),
    .A(\soc_inst.cpu_core.alu.a[21] ),
    .B(net4839));
 sg13g2_o21ai_1 _17130_ (.B1(_02869_),
    .Y(_02870_),
    .A1(_05800_),
    .A2(net4839));
 sg13g2_nand2_1 _17131_ (.Y(_02871_),
    .A(net4859),
    .B(net4840));
 sg13g2_o21ai_1 _17132_ (.B1(_02871_),
    .Y(_02872_),
    .A1(_05796_),
    .A2(net4840));
 sg13g2_mux2_1 _17133_ (.A0(_02870_),
    .A1(_02872_),
    .S(net4827),
    .X(_02873_));
 sg13g2_nor2b_1 _17134_ (.A(net4845),
    .B_N(\soc_inst.cpu_core.alu.a[16] ),
    .Y(_02874_));
 sg13g2_a21oi_1 _17135_ (.A1(\soc_inst.cpu_core.alu.a[17] ),
    .A2(net4846),
    .Y(_02875_),
    .B1(_02874_));
 sg13g2_nor2b_1 _17136_ (.A(net4839),
    .B_N(net4862),
    .Y(_02876_));
 sg13g2_a21oi_1 _17137_ (.A1(net4861),
    .A2(net4839),
    .Y(_02877_),
    .B1(_02876_));
 sg13g2_mux4_1 _17138_ (.S0(net4845),
    .A0(\soc_inst.cpu_core.alu.a[16] ),
    .A1(\soc_inst.cpu_core.alu.a[17] ),
    .A2(net4862),
    .A3(\soc_inst.cpu_core.alu.a[19] ),
    .S1(net4831),
    .X(_02878_));
 sg13g2_and2_1 _17139_ (.A(net4721),
    .B(_02878_),
    .X(_02879_));
 sg13g2_a21oi_1 _17140_ (.A1(net4820),
    .A2(_02873_),
    .Y(_02880_),
    .B1(_02879_));
 sg13g2_nor2b_1 _17141_ (.A(net4842),
    .B_N(net4855),
    .Y(_02881_));
 sg13g2_a21oi_1 _17142_ (.A1(\soc_inst.cpu_core.alu.a[29] ),
    .A2(net4842),
    .Y(_02882_),
    .B1(_02881_));
 sg13g2_nor2b_1 _17143_ (.A(net4843),
    .B_N(\soc_inst.cpu_core.alu.a[30] ),
    .Y(_02883_));
 sg13g2_a21o_1 _17144_ (.A2(net4842),
    .A1(net4853),
    .B1(_02883_),
    .X(_02884_));
 sg13g2_nand2_1 _17145_ (.Y(_02885_),
    .A(net4824),
    .B(_02884_));
 sg13g2_o21ai_1 _17146_ (.B1(_02885_),
    .Y(_02886_),
    .A1(net4824),
    .A2(_02882_));
 sg13g2_nor2b_1 _17147_ (.A(net4841),
    .B_N(\soc_inst.cpu_core.alu.a[24] ),
    .Y(_02887_));
 sg13g2_a21oi_1 _17148_ (.A1(net4858),
    .A2(net4841),
    .Y(_02888_),
    .B1(_02887_));
 sg13g2_mux2_1 _17149_ (.A0(net4856),
    .A1(\soc_inst.cpu_core.alu.a[27] ),
    .S(net4842),
    .X(_02889_));
 sg13g2_nand2_1 _17150_ (.Y(_02890_),
    .A(net4824),
    .B(_02889_));
 sg13g2_o21ai_1 _17151_ (.B1(_02890_),
    .Y(_02891_),
    .A1(net4825),
    .A2(_02888_));
 sg13g2_mux2_1 _17152_ (.A0(_02886_),
    .A1(_02891_),
    .S(net4718),
    .X(_02892_));
 sg13g2_nor2_1 _17153_ (.A(net4730),
    .B(_02892_),
    .Y(_02893_));
 sg13g2_a21oi_1 _17154_ (.A1(net4730),
    .A2(_02880_),
    .Y(_02894_),
    .B1(_02893_));
 sg13g2_nand3_1 _17155_ (.B(_02668_),
    .C(_02894_),
    .A(net4803),
    .Y(_02895_));
 sg13g2_nand2_1 _17156_ (.Y(_02896_),
    .A(net4863),
    .B(net4846));
 sg13g2_o21ai_1 _17157_ (.B1(_02896_),
    .Y(_02897_),
    .A1(_05816_),
    .A2(net4846));
 sg13g2_nand2_1 _17158_ (.Y(_02898_),
    .A(\soc_inst.cpu_core.alu.a[15] ),
    .B(net4847));
 sg13g2_o21ai_1 _17159_ (.B1(_02898_),
    .Y(_02899_),
    .A1(_05812_),
    .A2(net4846));
 sg13g2_mux2_1 _17160_ (.A0(_02897_),
    .A1(_02899_),
    .S(net4831),
    .X(_02900_));
 sg13g2_nand2_1 _17161_ (.Y(_02901_),
    .A(net4820),
    .B(_02900_));
 sg13g2_nand2_1 _17162_ (.Y(_02902_),
    .A(\soc_inst.cpu_core.alu.a[8] ),
    .B(_05839_));
 sg13g2_o21ai_1 _17163_ (.B1(_02902_),
    .Y(_02903_),
    .A1(_05822_),
    .A2(_05839_));
 sg13g2_nor2_1 _17164_ (.A(net4836),
    .B(_02903_),
    .Y(_02904_));
 sg13g2_nor2_1 _17165_ (.A(_05820_),
    .B(net4849),
    .Y(_02905_));
 sg13g2_a21oi_2 _17166_ (.B1(_02905_),
    .Y(_02906_),
    .A2(net4849),
    .A1(\soc_inst.cpu_core.alu.a[11] ));
 sg13g2_a21oi_1 _17167_ (.A1(net4837),
    .A2(_02906_),
    .Y(_02907_),
    .B1(_02904_));
 sg13g2_inv_1 _17168_ (.Y(_02908_),
    .A(_02907_));
 sg13g2_o21ai_1 _17169_ (.B1(_02901_),
    .Y(_02909_),
    .A1(net4820),
    .A2(_02908_));
 sg13g2_nor2_1 _17170_ (.A(net4803),
    .B(_02669_),
    .Y(_02910_));
 sg13g2_nand2_2 _17171_ (.Y(_02911_),
    .A(net4735),
    .B(_02668_));
 sg13g2_nand2_1 _17172_ (.Y(_02912_),
    .A(\soc_inst.cpu_core.alu.a[5] ),
    .B(net4852));
 sg13g2_o21ai_1 _17173_ (.B1(_02912_),
    .Y(_02913_),
    .A1(_05832_),
    .A2(net4852));
 sg13g2_inv_1 _17174_ (.Y(_02914_),
    .A(_02913_));
 sg13g2_nor2_1 _17175_ (.A(net4833),
    .B(_02913_),
    .Y(_02915_));
 sg13g2_nor2_1 _17176_ (.A(_05828_),
    .B(net4852),
    .Y(_02916_));
 sg13g2_nand2_1 _17177_ (.Y(_02917_),
    .A(\soc_inst.cpu_core.alu.a[7] ),
    .B(net4852));
 sg13g2_nor2b_1 _17178_ (.A(_02916_),
    .B_N(_02917_),
    .Y(_02918_));
 sg13g2_a21oi_1 _17179_ (.A1(net4836),
    .A2(_02918_),
    .Y(_02919_),
    .B1(_02915_));
 sg13g2_nand2_1 _17180_ (.Y(_02920_),
    .A(net4864),
    .B(_05839_));
 sg13g2_nand2_1 _17181_ (.Y(_02921_),
    .A(\soc_inst.cpu_core.alu.a[3] ),
    .B(net4849));
 sg13g2_nand2_1 _17182_ (.Y(_02922_),
    .A(_02920_),
    .B(_02921_));
 sg13g2_nor2b_2 _17183_ (.A(net4821),
    .B_N(net4834),
    .Y(_02923_));
 sg13g2_nor2_2 _17184_ (.A(net4821),
    .B(net4829),
    .Y(_02924_));
 sg13g2_or2_1 _17185_ (.X(_02925_),
    .B(net4834),
    .A(net4821));
 sg13g2_nor2b_1 _17186_ (.A(net4848),
    .B_N(\soc_inst.cpu_core.alu.a[0] ),
    .Y(_02926_));
 sg13g2_nand2_2 _17187_ (.Y(_02927_),
    .A(_05839_),
    .B(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_nor2_1 _17188_ (.A(net4659),
    .B(_02927_),
    .Y(_02928_));
 sg13g2_nand2_1 _17189_ (.Y(_02929_),
    .A(\soc_inst.cpu_core.alu.a[1] ),
    .B(net4848));
 sg13g2_a21oi_1 _17190_ (.A1(_02927_),
    .A2(_02929_),
    .Y(_02930_),
    .B1(net4659));
 sg13g2_a221oi_1 _17191_ (.B2(_02923_),
    .C1(_02930_),
    .B1(_02922_),
    .A1(net4822),
    .Y(_02931_),
    .A2(_02919_));
 sg13g2_o21ai_1 _17192_ (.B1(net4213),
    .Y(_02932_),
    .A1(net4733),
    .A2(_02909_));
 sg13g2_a21oi_1 _17193_ (.A1(net4733),
    .A2(_02931_),
    .Y(_02933_),
    .B1(_02932_));
 sg13g2_nor2b_2 _17194_ (.A(net4865),
    .B_N(\soc_inst.cpu_core.alu.op[2] ),
    .Y(_02934_));
 sg13g2_and2_1 _17195_ (.A(_02863_),
    .B(_02934_),
    .X(_02935_));
 sg13g2_nand2_2 _17196_ (.Y(_02936_),
    .A(_02863_),
    .B(_02934_));
 sg13g2_and2_1 _17197_ (.A(net4848),
    .B(\soc_inst.cpu_core.alu.a[0] ),
    .X(_02937_));
 sg13g2_nand2_1 _17198_ (.Y(_02938_),
    .A(net4848),
    .B(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_nand2_1 _17199_ (.Y(_02939_),
    .A(\soc_inst.cpu_core.alu.op[2] ),
    .B(net4865));
 sg13g2_nand3_1 _17200_ (.B(_02938_),
    .C(_02939_),
    .A(_02665_),
    .Y(_02940_));
 sg13g2_nand2_1 _17201_ (.Y(_02941_),
    .A(_02936_),
    .B(_02940_));
 sg13g2_o21ai_1 _17202_ (.B1(_02941_),
    .Y(_02942_),
    .A1(net4848),
    .A2(net2345));
 sg13g2_nor3_1 _17203_ (.A(net4814),
    .B(net4659),
    .C(_02927_),
    .Y(_02943_));
 sg13g2_and2_1 _17204_ (.A(_02667_),
    .B(_02862_),
    .X(_02944_));
 sg13g2_nand2_2 _17205_ (.Y(_02945_),
    .A(_02667_),
    .B(_02862_));
 sg13g2_nor2_1 _17206_ (.A(net4805),
    .B(_02945_),
    .Y(_02946_));
 sg13g2_nand2_2 _17207_ (.Y(_02947_),
    .A(net4736),
    .B(_02944_));
 sg13g2_nor2b_1 _17208_ (.A(_02866_),
    .B_N(_02934_),
    .Y(_02948_));
 sg13g2_nand2b_2 _17209_ (.Y(_02949_),
    .B(_02934_),
    .A_N(_02866_));
 sg13g2_a221oi_1 _17210_ (.B2(_02937_),
    .C1(_02933_),
    .B1(net4435),
    .A1(_02943_),
    .Y(_02950_),
    .A2(net4211));
 sg13g2_nand4_1 _17211_ (.B(_02895_),
    .C(_02942_),
    .A(_02868_),
    .Y(_02951_),
    .D(_02950_));
 sg13g2_o21ai_1 _17212_ (.B1(_02673_),
    .Y(_02952_),
    .A1(_02865_),
    .A2(_02951_));
 sg13g2_o21ai_1 _17213_ (.B1(_02952_),
    .Y(_01386_),
    .A1(_05478_),
    .A2(net4746));
 sg13g2_nor2_2 _17214_ (.A(net4865),
    .B(_02669_),
    .Y(_02953_));
 sg13g2_inv_2 _17215_ (.Y(_02954_),
    .A(_02953_));
 sg13g2_mux4_1 _17216_ (.S0(net4841),
    .A0(\soc_inst.cpu_core.alu.a[21] ),
    .A1(\soc_inst.cpu_core.alu.a[22] ),
    .A2(net4859),
    .A3(\soc_inst.cpu_core.alu.a[24] ),
    .S1(net4826),
    .X(_02955_));
 sg13g2_nand2_1 _17217_ (.Y(_02956_),
    .A(net4862),
    .B(net4845));
 sg13g2_o21ai_1 _17218_ (.B1(_02956_),
    .Y(_02957_),
    .A1(_05806_),
    .A2(net4840));
 sg13g2_nand2_1 _17219_ (.Y(_02958_),
    .A(net4860),
    .B(net4839));
 sg13g2_o21ai_1 _17220_ (.B1(_02958_),
    .Y(_02959_),
    .A1(_05802_),
    .A2(net4839));
 sg13g2_mux2_1 _17221_ (.A0(_02957_),
    .A1(_02959_),
    .S(net4827),
    .X(_02960_));
 sg13g2_mux2_1 _17222_ (.A0(_02955_),
    .A1(_02960_),
    .S(net4718),
    .X(_02961_));
 sg13g2_nand2_1 _17223_ (.Y(_02962_),
    .A(net4729),
    .B(_02961_));
 sg13g2_nor2b_1 _17224_ (.A(net4843),
    .B_N(\soc_inst.cpu_core.alu.a[27] ),
    .Y(_02963_));
 sg13g2_and2_1 _17225_ (.A(net4855),
    .B(net4843),
    .X(_02964_));
 sg13g2_mux4_1 _17226_ (.S0(net4842),
    .A0(net4858),
    .A1(net4856),
    .A2(\soc_inst.cpu_core.alu.a[27] ),
    .A3(net4855),
    .S1(net4824),
    .X(_02965_));
 sg13g2_and2_1 _17227_ (.A(net4718),
    .B(_02965_),
    .X(_02966_));
 sg13g2_nor2b_1 _17228_ (.A(net4842),
    .B_N(net4854),
    .Y(_02967_));
 sg13g2_nor2b_1 _17229_ (.A(net4843),
    .B_N(\soc_inst.cpu_core.alu.a[29] ),
    .Y(_02968_));
 sg13g2_a21oi_1 _17230_ (.A1(\soc_inst.cpu_core.alu.a[30] ),
    .A2(net4842),
    .Y(_02969_),
    .B1(_02968_));
 sg13g2_nor2_1 _17231_ (.A(net4829),
    .B(_02969_),
    .Y(_02970_));
 sg13g2_a21o_1 _17232_ (.A2(_02967_),
    .A1(net4829),
    .B1(_02970_),
    .X(_02971_));
 sg13g2_a21oi_1 _17233_ (.A1(net4817),
    .A2(_02971_),
    .Y(_02972_),
    .B1(_02966_));
 sg13g2_o21ai_1 _17234_ (.B1(_02962_),
    .Y(_02973_),
    .A1(net4729),
    .A2(_02972_));
 sg13g2_and2_1 _17235_ (.A(net4865),
    .B(_02668_),
    .X(_02974_));
 sg13g2_nand3_1 _17236_ (.B(net4817),
    .C(net4824),
    .A(net4853),
    .Y(_02975_));
 sg13g2_a21o_1 _17237_ (.A2(net4829),
    .A1(net4853),
    .B1(_02970_),
    .X(_02976_));
 sg13g2_a21oi_1 _17238_ (.A1(net4817),
    .A2(_02976_),
    .Y(_02977_),
    .B1(_02966_));
 sg13g2_o21ai_1 _17239_ (.B1(_02962_),
    .Y(_02978_),
    .A1(net4729),
    .A2(_02977_));
 sg13g2_a22oi_1 _17240_ (.Y(_02979_),
    .B1(_02974_),
    .B2(_02978_),
    .A2(_02973_),
    .A1(_02953_));
 sg13g2_inv_1 _17241_ (.Y(_02980_),
    .A(_02979_));
 sg13g2_nand2_1 _17242_ (.Y(_02981_),
    .A(\soc_inst.cpu_core.alu.a[6] ),
    .B(net4852));
 sg13g2_o21ai_1 _17243_ (.B1(_02981_),
    .Y(_02982_),
    .A1(_05830_),
    .A2(net4852));
 sg13g2_nor2_1 _17244_ (.A(net4833),
    .B(_02982_),
    .Y(_02983_));
 sg13g2_nor2b_1 _17245_ (.A(net4852),
    .B_N(\soc_inst.cpu_core.alu.a[7] ),
    .Y(_02984_));
 sg13g2_a21oi_1 _17246_ (.A1(\soc_inst.cpu_core.alu.a[8] ),
    .A2(net4850),
    .Y(_02985_),
    .B1(_02984_));
 sg13g2_a21oi_1 _17247_ (.A1(net4833),
    .A2(_02985_),
    .Y(_02986_),
    .B1(_02983_));
 sg13g2_nor2b_1 _17248_ (.A(net4848),
    .B_N(\soc_inst.cpu_core.alu.a[1] ),
    .Y(_02987_));
 sg13g2_a21oi_1 _17249_ (.A1(net4864),
    .A2(net4848),
    .Y(_02988_),
    .B1(_02987_));
 sg13g2_nand2_1 _17250_ (.Y(_02989_),
    .A(\soc_inst.cpu_core.alu.a[4] ),
    .B(net4850));
 sg13g2_nor2b_1 _17251_ (.A(net4849),
    .B_N(\soc_inst.cpu_core.alu.a[3] ),
    .Y(_02990_));
 sg13g2_a21oi_1 _17252_ (.A1(\soc_inst.cpu_core.alu.a[4] ),
    .A2(net4849),
    .Y(_02991_),
    .B1(_02990_));
 sg13g2_a22oi_1 _17253_ (.Y(_02992_),
    .B1(_02991_),
    .B2(_02923_),
    .A2(_02988_),
    .A1(_02924_));
 sg13g2_o21ai_1 _17254_ (.B1(_02992_),
    .Y(_02993_),
    .A1(net4725),
    .A2(_02986_));
 sg13g2_nand2_1 _17255_ (.Y(_02994_),
    .A(\soc_inst.cpu_core.alu.a[14] ),
    .B(net4847));
 sg13g2_o21ai_1 _17256_ (.B1(_02994_),
    .Y(_02995_),
    .A1(_05814_),
    .A2(net4852));
 sg13g2_nand2_1 _17257_ (.Y(_02996_),
    .A(\soc_inst.cpu_core.alu.a[16] ),
    .B(net4845));
 sg13g2_o21ai_1 _17258_ (.B1(_02996_),
    .Y(_02997_),
    .A1(_05810_),
    .A2(net4845));
 sg13g2_mux2_1 _17259_ (.A0(_02995_),
    .A1(_02997_),
    .S(net4832),
    .X(_02998_));
 sg13g2_nand2_1 _17260_ (.Y(_02999_),
    .A(\soc_inst.cpu_core.alu.a[9] ),
    .B(_05839_));
 sg13g2_o21ai_1 _17261_ (.B1(_02999_),
    .Y(_03000_),
    .A1(_05820_),
    .A2(_05839_));
 sg13g2_nor2_1 _17262_ (.A(net4834),
    .B(_03000_),
    .Y(_03001_));
 sg13g2_nor2b_1 _17263_ (.A(net4851),
    .B_N(\soc_inst.cpu_core.alu.a[11] ),
    .Y(_03002_));
 sg13g2_a21oi_1 _17264_ (.A1(\soc_inst.cpu_core.alu.a[12] ),
    .A2(net4851),
    .Y(_03003_),
    .B1(_03002_));
 sg13g2_a21oi_1 _17265_ (.A1(net4833),
    .A2(_03003_),
    .Y(_03004_),
    .B1(_03001_));
 sg13g2_mux2_1 _17266_ (.A0(_02998_),
    .A1(_03004_),
    .S(net4726),
    .X(_03005_));
 sg13g2_nor2_1 _17267_ (.A(net4732),
    .B(_03005_),
    .Y(_03006_));
 sg13g2_a21oi_1 _17268_ (.A1(net4732),
    .A2(_02993_),
    .Y(_03007_),
    .B1(_03006_));
 sg13g2_xnor2_1 _17269_ (.Y(_03008_),
    .A(_02737_),
    .B(_02738_));
 sg13g2_o21ai_1 _17270_ (.B1(net4742),
    .Y(_03009_),
    .A1(_02736_),
    .A2(net4433));
 sg13g2_and2_1 _17271_ (.A(_02665_),
    .B(_02934_),
    .X(_03010_));
 sg13g2_nand2_2 _17272_ (.Y(_03011_),
    .A(_02665_),
    .B(_02934_));
 sg13g2_o21ai_1 _17273_ (.B1(net4439),
    .Y(_03012_),
    .A1(net4830),
    .A2(\soc_inst.cpu_core.alu.a[1] ));
 sg13g2_o21ai_1 _17274_ (.B1(_03012_),
    .Y(_03013_),
    .A1(_02737_),
    .A2(_03011_));
 sg13g2_and2_1 _17275_ (.A(_02665_),
    .B(_02862_),
    .X(_03014_));
 sg13g2_nand2_2 _17276_ (.Y(_03015_),
    .A(_02665_),
    .B(_02862_));
 sg13g2_xnor2_1 _17277_ (.Y(_03016_),
    .A(_02737_),
    .B(_02937_));
 sg13g2_nor2_2 _17278_ (.A(net4812),
    .B(_02945_),
    .Y(_03017_));
 sg13g2_or2_1 _17279_ (.X(_03018_),
    .B(_02987_),
    .A(_02937_));
 sg13g2_nand3_1 _17280_ (.B(net4210),
    .C(_03018_),
    .A(_02924_),
    .Y(_03019_));
 sg13g2_nor2_1 _17281_ (.A(net4804),
    .B(_03019_),
    .Y(_03020_));
 sg13g2_nor3_1 _17282_ (.A(_03009_),
    .B(_03013_),
    .C(_03020_),
    .Y(_03021_));
 sg13g2_a22oi_1 _17283_ (.Y(_03022_),
    .B1(net4426),
    .B2(_03016_),
    .A2(_03007_),
    .A1(net4214));
 sg13g2_o21ai_1 _17284_ (.B1(_03021_),
    .Y(_03023_),
    .A1(net4445),
    .A2(_03008_));
 sg13g2_a21oi_1 _17285_ (.A1(net4804),
    .A2(_02980_),
    .Y(_03024_),
    .B1(_03023_));
 sg13g2_a22oi_1 _17286_ (.Y(_01387_),
    .B1(_03022_),
    .B2(_03024_),
    .A2(net4885),
    .A1(_05477_));
 sg13g2_nand2_1 _17287_ (.Y(_03025_),
    .A(net4827),
    .B(_02870_));
 sg13g2_o21ai_1 _17288_ (.B1(_03025_),
    .Y(_03026_),
    .A1(net4827),
    .A2(_02877_));
 sg13g2_nor2_1 _17289_ (.A(net4826),
    .B(_02872_),
    .Y(_03027_));
 sg13g2_a21oi_1 _17290_ (.A1(net4826),
    .A2(_02888_),
    .Y(_03028_),
    .B1(_03027_));
 sg13g2_mux2_1 _17291_ (.A0(_03026_),
    .A1(_03028_),
    .S(net4818),
    .X(_03029_));
 sg13g2_nand2_1 _17292_ (.Y(_03030_),
    .A(net4728),
    .B(_03029_));
 sg13g2_nor2_2 _17293_ (.A(net4726),
    .B(net4829),
    .Y(_03031_));
 sg13g2_nor2_1 _17294_ (.A(net4824),
    .B(_02889_),
    .Y(_03032_));
 sg13g2_a21oi_1 _17295_ (.A1(net4824),
    .A2(_02882_),
    .Y(_03033_),
    .B1(_03032_));
 sg13g2_a22oi_1 _17296_ (.Y(_03034_),
    .B1(_03033_),
    .B2(net4718),
    .A2(_03031_),
    .A1(_02884_));
 sg13g2_inv_1 _17297_ (.Y(_03035_),
    .A(_03034_));
 sg13g2_o21ai_1 _17298_ (.B1(_03030_),
    .Y(_03036_),
    .A1(net4728),
    .A2(_03034_));
 sg13g2_nand2_1 _17299_ (.Y(_03037_),
    .A(_02975_),
    .B(_03034_));
 sg13g2_nand2_1 _17300_ (.Y(_03038_),
    .A(net4808),
    .B(_03037_));
 sg13g2_nand2_1 _17301_ (.Y(_03039_),
    .A(_03030_),
    .B(_03038_));
 sg13g2_a22oi_1 _17302_ (.Y(_03040_),
    .B1(_03039_),
    .B2(_02974_),
    .A2(_03036_),
    .A1(_02953_));
 sg13g2_inv_1 _17303_ (.Y(_03041_),
    .A(_03040_));
 sg13g2_nand2_1 _17304_ (.Y(_03042_),
    .A(net4836),
    .B(_02903_));
 sg13g2_o21ai_1 _17305_ (.B1(_03042_),
    .Y(_03043_),
    .A1(net4836),
    .A2(_02918_));
 sg13g2_inv_1 _17306_ (.Y(_03044_),
    .A(_03043_));
 sg13g2_a22oi_1 _17307_ (.Y(_03045_),
    .B1(_03044_),
    .B2(net4821),
    .A2(_02923_),
    .A1(_02914_));
 sg13g2_o21ai_1 _17308_ (.B1(_03045_),
    .Y(_03046_),
    .A1(_02922_),
    .A2(net4659));
 sg13g2_nor2_1 _17309_ (.A(net4831),
    .B(_02899_),
    .Y(_03047_));
 sg13g2_a21oi_1 _17310_ (.A1(net4831),
    .A2(_02875_),
    .Y(_03048_),
    .B1(_03047_));
 sg13g2_nand2_1 _17311_ (.Y(_03049_),
    .A(net4830),
    .B(_02897_));
 sg13g2_o21ai_1 _17312_ (.B1(_03049_),
    .Y(_03050_),
    .A1(net4830),
    .A2(_02906_));
 sg13g2_mux2_1 _17313_ (.A0(_03048_),
    .A1(_03050_),
    .S(net4721),
    .X(_03051_));
 sg13g2_a21oi_1 _17314_ (.A1(net4732),
    .A2(_03046_),
    .Y(_03052_),
    .B1(_02911_));
 sg13g2_o21ai_1 _17315_ (.B1(_03052_),
    .Y(_03053_),
    .A1(net4732),
    .A2(_03051_));
 sg13g2_o21ai_1 _17316_ (.B1(_02736_),
    .Y(_03054_),
    .A1(_02737_),
    .A2(_02938_));
 sg13g2_xnor2_1 _17317_ (.Y(_03055_),
    .A(_02734_),
    .B(_03054_));
 sg13g2_o21ai_1 _17318_ (.B1(net4440),
    .Y(_03056_),
    .A1(net4823),
    .A2(net4864));
 sg13g2_a221oi_1 _17319_ (.B2(_02733_),
    .C1(net4886),
    .B1(net4429),
    .A1(_02732_),
    .Y(_03057_),
    .A2(net4435));
 sg13g2_nand2_1 _17320_ (.Y(_03058_),
    .A(_02920_),
    .B(_02929_));
 sg13g2_nand2_1 _17321_ (.Y(_03059_),
    .A(net4830),
    .B(_02927_));
 sg13g2_o21ai_1 _17322_ (.B1(_03059_),
    .Y(_03060_),
    .A1(net4830),
    .A2(_03058_));
 sg13g2_nand2b_1 _17323_ (.Y(_03061_),
    .B(net4723),
    .A_N(_03060_));
 sg13g2_nor2_2 _17324_ (.A(net4814),
    .B(_03061_),
    .Y(_03062_));
 sg13g2_a21oi_1 _17325_ (.A1(_02734_),
    .A2(_02739_),
    .Y(_03063_),
    .B1(net4445));
 sg13g2_o21ai_1 _17326_ (.B1(_03063_),
    .Y(_03064_),
    .A1(_02734_),
    .A2(_02739_));
 sg13g2_a22oi_1 _17327_ (.Y(_03065_),
    .B1(_03062_),
    .B2(net4211),
    .A2(_03055_),
    .A1(net4426));
 sg13g2_nand4_1 _17328_ (.B(_03057_),
    .C(_03064_),
    .A(_03056_),
    .Y(_03066_),
    .D(_03065_));
 sg13g2_a21oi_1 _17329_ (.A1(net4807),
    .A2(_03041_),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_a22oi_1 _17330_ (.Y(_01388_),
    .B1(_03053_),
    .B2(_03067_),
    .A2(_05758_),
    .A1(net4887));
 sg13g2_mux4_1 _17331_ (.S0(net4841),
    .A0(net4859),
    .A1(\soc_inst.cpu_core.alu.a[24] ),
    .A2(net4858),
    .A3(net4856),
    .S1(net4826),
    .X(_03068_));
 sg13g2_mux4_1 _17332_ (.S0(net4840),
    .A0(net4861),
    .A1(net4860),
    .A2(\soc_inst.cpu_core.alu.a[21] ),
    .A3(\soc_inst.cpu_core.alu.a[22] ),
    .S1(net4827),
    .X(_03069_));
 sg13g2_mux2_1 _17333_ (.A0(_03068_),
    .A1(_03069_),
    .S(net4718),
    .X(_03070_));
 sg13g2_nand2_1 _17334_ (.Y(_03071_),
    .A(net4729),
    .B(_03070_));
 sg13g2_nor3_1 _17335_ (.A(net4829),
    .B(_02963_),
    .C(_02964_),
    .Y(_03072_));
 sg13g2_a21oi_1 _17336_ (.A1(net4829),
    .A2(_02969_),
    .Y(_03073_),
    .B1(_03072_));
 sg13g2_and2_1 _17337_ (.A(net4719),
    .B(_03073_),
    .X(_03074_));
 sg13g2_a21o_1 _17338_ (.A2(_03031_),
    .A1(_02967_),
    .B1(_03074_),
    .X(_03075_));
 sg13g2_nand2_1 _17339_ (.Y(_03076_),
    .A(net4810),
    .B(_03075_));
 sg13g2_nand2_1 _17340_ (.Y(_03077_),
    .A(_03071_),
    .B(_03076_));
 sg13g2_a21oi_1 _17341_ (.A1(net4853),
    .A2(net4817),
    .Y(_03078_),
    .B1(_03074_));
 sg13g2_inv_1 _17342_ (.Y(_03079_),
    .A(_03078_));
 sg13g2_o21ai_1 _17343_ (.B1(_03071_),
    .Y(_03080_),
    .A1(net4728),
    .A2(_03078_));
 sg13g2_a22oi_1 _17344_ (.Y(_03081_),
    .B1(_03080_),
    .B2(_02974_),
    .A2(_03077_),
    .A1(_02953_));
 sg13g2_nand2b_1 _17345_ (.Y(_03082_),
    .B(net4807),
    .A_N(_03081_));
 sg13g2_a21oi_1 _17346_ (.A1(_02733_),
    .A2(_03054_),
    .Y(_03083_),
    .B1(_02732_));
 sg13g2_xor2_1 _17347_ (.B(_03083_),
    .A(_02730_),
    .X(_03084_));
 sg13g2_xor2_1 _17348_ (.B(_02740_),
    .A(_02730_),
    .X(_03085_));
 sg13g2_mux2_1 _17349_ (.A0(_02997_),
    .A1(_02957_),
    .S(net4828),
    .X(_03086_));
 sg13g2_nand2_1 _17350_ (.Y(_03087_),
    .A(net4833),
    .B(_02995_));
 sg13g2_o21ai_1 _17351_ (.B1(_03087_),
    .Y(_03088_),
    .A1(net4833),
    .A2(_03003_));
 sg13g2_mux2_1 _17352_ (.A0(_03086_),
    .A1(_03088_),
    .S(net4726),
    .X(_03089_));
 sg13g2_inv_1 _17353_ (.Y(_03090_),
    .A(_03089_));
 sg13g2_nand2_1 _17354_ (.Y(_03091_),
    .A(net4833),
    .B(_03000_));
 sg13g2_o21ai_1 _17355_ (.B1(_03091_),
    .Y(_03092_),
    .A1(net4833),
    .A2(_02985_));
 sg13g2_o21ai_1 _17356_ (.B1(net4732),
    .Y(_03093_),
    .A1(_02925_),
    .A2(_02991_));
 sg13g2_a221oi_1 _17357_ (.B2(net4821),
    .C1(_03093_),
    .B1(_03092_),
    .A1(_02923_),
    .Y(_03094_),
    .A2(_02982_));
 sg13g2_a21oi_1 _17358_ (.A1(net4815),
    .A2(_03090_),
    .Y(_03095_),
    .B1(_03094_));
 sg13g2_a21oi_1 _17359_ (.A1(net4864),
    .A2(net4849),
    .Y(_03096_),
    .B1(_02990_));
 sg13g2_nand2_1 _17360_ (.Y(_03097_),
    .A(net4837),
    .B(_03018_));
 sg13g2_o21ai_1 _17361_ (.B1(_03097_),
    .Y(_03098_),
    .A1(net4835),
    .A2(_03096_));
 sg13g2_nand2_2 _17362_ (.Y(_03099_),
    .A(net4724),
    .B(_03098_));
 sg13g2_nor2_1 _17363_ (.A(net4816),
    .B(_03099_),
    .Y(_03100_));
 sg13g2_a221oi_1 _17364_ (.B2(_02730_),
    .C1(net4880),
    .B1(net4430),
    .A1(_02727_),
    .Y(_03101_),
    .A2(net4436));
 sg13g2_o21ai_1 _17365_ (.B1(_03101_),
    .Y(_03102_),
    .A1(_02729_),
    .A2(_02936_));
 sg13g2_a221oi_1 _17366_ (.B2(net4212),
    .C1(_03102_),
    .B1(_03100_),
    .A1(net4214),
    .Y(_03103_),
    .A2(_03095_));
 sg13g2_o21ai_1 _17367_ (.B1(_03103_),
    .Y(_03104_),
    .A1(_03015_),
    .A2(_03084_));
 sg13g2_a21oi_1 _17368_ (.A1(net4447),
    .A2(_03085_),
    .Y(_03105_),
    .B1(_03104_));
 sg13g2_a22oi_1 _17369_ (.Y(_01389_),
    .B1(_03082_),
    .B2(_03105_),
    .A2(_05759_),
    .A1(net4885));
 sg13g2_o21ai_1 _17370_ (.B1(_02728_),
    .Y(_03106_),
    .A1(_02729_),
    .A2(_03083_));
 sg13g2_nand2b_1 _17371_ (.Y(_03107_),
    .B(_02725_),
    .A_N(_03106_));
 sg13g2_nand2b_1 _17372_ (.Y(_03108_),
    .B(_03106_),
    .A_N(_02725_));
 sg13g2_nand3_1 _17373_ (.B(_03107_),
    .C(_03108_),
    .A(net4426),
    .Y(_03109_));
 sg13g2_xnor2_1 _17374_ (.Y(_03110_),
    .A(_02725_),
    .B(_02741_));
 sg13g2_o21ai_1 _17375_ (.B1(_03109_),
    .Y(_03111_),
    .A1(net4444),
    .A2(_03110_));
 sg13g2_mux2_1 _17376_ (.A0(_02873_),
    .A1(_02891_),
    .S(net4819),
    .X(_03112_));
 sg13g2_inv_1 _17377_ (.Y(_03113_),
    .A(_03112_));
 sg13g2_nor2_1 _17378_ (.A(net4809),
    .B(_03113_),
    .Y(_03114_));
 sg13g2_and2_1 _17379_ (.A(net4718),
    .B(_02886_),
    .X(_03115_));
 sg13g2_a21o_1 _17380_ (.A2(_03115_),
    .A1(net4809),
    .B1(_03114_),
    .X(_03116_));
 sg13g2_a21o_1 _17381_ (.A2(net4819),
    .A1(net4853),
    .B1(_03115_),
    .X(_03117_));
 sg13g2_a21o_1 _17382_ (.A2(_03117_),
    .A1(net4809),
    .B1(_03114_),
    .X(_03118_));
 sg13g2_a22oi_1 _17383_ (.Y(_03119_),
    .B1(_03118_),
    .B2(_02974_),
    .A2(_03116_),
    .A1(_02953_));
 sg13g2_nor2_1 _17384_ (.A(net4735),
    .B(_03119_),
    .Y(_03120_));
 sg13g2_mux2_1 _17385_ (.A0(_02878_),
    .A1(_02900_),
    .S(net4721),
    .X(_03121_));
 sg13g2_a21oi_1 _17386_ (.A1(net4821),
    .A2(_02908_),
    .Y(_03122_),
    .B1(net4814));
 sg13g2_o21ai_1 _17387_ (.B1(_03122_),
    .Y(_03123_),
    .A1(net4822),
    .A2(_02919_));
 sg13g2_nand2_1 _17388_ (.Y(_03124_),
    .A(net4811),
    .B(_03121_));
 sg13g2_a21oi_1 _17389_ (.A1(_03123_),
    .A2(_03124_),
    .Y(_03125_),
    .B1(_02911_));
 sg13g2_o21ai_1 _17390_ (.B1(_02921_),
    .Y(_03126_),
    .A1(_05832_),
    .A2(net4849));
 sg13g2_mux2_1 _17391_ (.A0(_03126_),
    .A1(_03058_),
    .S(net4835),
    .X(_03127_));
 sg13g2_a22oi_1 _17392_ (.Y(_03128_),
    .B1(_03127_),
    .B2(net4723),
    .A2(_03031_),
    .A1(_02926_));
 sg13g2_or2_1 _17393_ (.X(_03129_),
    .B(_03128_),
    .A(net4811));
 sg13g2_o21ai_1 _17394_ (.B1(_02936_),
    .Y(_03130_),
    .A1(_02724_),
    .A2(_03011_));
 sg13g2_a221oi_1 _17395_ (.B2(_02723_),
    .C1(net4881),
    .B1(_03130_),
    .A1(_02724_),
    .Y(_03131_),
    .A2(net4435));
 sg13g2_o21ai_1 _17396_ (.B1(_03131_),
    .Y(_03132_),
    .A1(_02947_),
    .A2(_03129_));
 sg13g2_nor4_2 _17397_ (.A(_03111_),
    .B(_03120_),
    .C(_03125_),
    .Y(_03133_),
    .D(_03132_));
 sg13g2_a21oi_1 _17398_ (.A1(net4908),
    .A2(_05760_),
    .Y(_01390_),
    .B1(_03133_));
 sg13g2_a21oi_1 _17399_ (.A1(_02719_),
    .A2(_02742_),
    .Y(_03134_),
    .B1(net4445));
 sg13g2_o21ai_1 _17400_ (.B1(_03134_),
    .Y(_03135_),
    .A1(_02719_),
    .A2(_02742_));
 sg13g2_a21oi_2 _17401_ (.B1(_02724_),
    .Y(_03136_),
    .A2(_03106_),
    .A1(_02723_));
 sg13g2_xnor2_1 _17402_ (.Y(_03137_),
    .A(_02719_),
    .B(_03136_));
 sg13g2_mux2_1 _17403_ (.A0(_02955_),
    .A1(_02965_),
    .S(net4818),
    .X(_03138_));
 sg13g2_and2_1 _17404_ (.A(net4728),
    .B(_03138_),
    .X(_03139_));
 sg13g2_and2_1 _17405_ (.A(net4718),
    .B(_02971_),
    .X(_03140_));
 sg13g2_a21oi_1 _17406_ (.A1(net4808),
    .A2(_03140_),
    .Y(_03141_),
    .B1(_03139_));
 sg13g2_nand2_1 _17407_ (.Y(_03142_),
    .A(net4853),
    .B(net4659));
 sg13g2_o21ai_1 _17408_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net4659),
    .A2(_02969_));
 sg13g2_a21oi_1 _17409_ (.A1(net4809),
    .A2(_03143_),
    .Y(_03144_),
    .B1(_03139_));
 sg13g2_nand2b_1 _17410_ (.Y(_03145_),
    .B(_02974_),
    .A_N(_03144_));
 sg13g2_o21ai_1 _17411_ (.B1(_03145_),
    .Y(_03146_),
    .A1(_02954_),
    .A2(_03141_));
 sg13g2_and2_1 _17412_ (.A(net4818),
    .B(_02960_),
    .X(_03147_));
 sg13g2_a21oi_1 _17413_ (.A1(net4720),
    .A2(_02998_),
    .Y(_03148_),
    .B1(_03147_));
 sg13g2_nand2_1 _17414_ (.Y(_03149_),
    .A(net4726),
    .B(_02986_));
 sg13g2_a21oi_1 _17415_ (.A1(net4821),
    .A2(_03004_),
    .Y(_03150_),
    .B1(net4815));
 sg13g2_a22oi_1 _17416_ (.Y(_03151_),
    .B1(_03149_),
    .B2(_03150_),
    .A2(_03148_),
    .A1(net4815));
 sg13g2_nand2b_1 _17417_ (.Y(_03152_),
    .B(net4435),
    .A_N(_02718_));
 sg13g2_a22oi_1 _17418_ (.Y(_03153_),
    .B1(net4429),
    .B2(_02719_),
    .A2(net4439),
    .A1(_02717_));
 sg13g2_o21ai_1 _17419_ (.B1(_02989_),
    .Y(_03154_),
    .A1(_05830_),
    .A2(net4850));
 sg13g2_nor2_1 _17420_ (.A(net4836),
    .B(_03154_),
    .Y(_03155_));
 sg13g2_a21oi_1 _17421_ (.A1(net4835),
    .A2(_03096_),
    .Y(_03156_),
    .B1(_03155_));
 sg13g2_a22oi_1 _17422_ (.Y(_03157_),
    .B1(_03156_),
    .B2(net4723),
    .A2(_03031_),
    .A1(_03018_));
 sg13g2_nor2_2 _17423_ (.A(net4814),
    .B(_03157_),
    .Y(_03158_));
 sg13g2_a22oi_1 _17424_ (.Y(_03159_),
    .B1(_03158_),
    .B2(net4211),
    .A2(_03151_),
    .A1(net4213));
 sg13g2_nand4_1 _17425_ (.B(_03152_),
    .C(_03153_),
    .A(net4742),
    .Y(_03160_),
    .D(_03159_));
 sg13g2_a221oi_1 _17426_ (.B2(net4806),
    .C1(_03160_),
    .B1(_03146_),
    .A1(net4426),
    .Y(_03161_),
    .A2(_03137_));
 sg13g2_a22oi_1 _17427_ (.Y(_01391_),
    .B1(_03135_),
    .B2(_03161_),
    .A2(_05761_),
    .A1(net4889));
 sg13g2_o21ai_1 _17428_ (.B1(_02718_),
    .Y(_03162_),
    .A1(_02720_),
    .A2(_03136_));
 sg13g2_o21ai_1 _17429_ (.B1(net4426),
    .Y(_03163_),
    .A1(_02714_),
    .A2(_03162_));
 sg13g2_a21o_1 _17430_ (.A2(_03162_),
    .A1(_02714_),
    .B1(_03163_),
    .X(_03164_));
 sg13g2_xnor2_1 _17431_ (.Y(_03165_),
    .A(_02714_),
    .B(_02743_));
 sg13g2_mux2_1 _17432_ (.A0(_03028_),
    .A1(_03033_),
    .S(net4818),
    .X(_03166_));
 sg13g2_inv_1 _17433_ (.Y(_03167_),
    .A(_03166_));
 sg13g2_nand2_1 _17434_ (.Y(_03168_),
    .A(net4728),
    .B(_03166_));
 sg13g2_and2_1 _17435_ (.A(_02884_),
    .B(_02924_),
    .X(_03169_));
 sg13g2_nand2_1 _17436_ (.Y(_03170_),
    .A(net4808),
    .B(_03169_));
 sg13g2_nand2_1 _17437_ (.Y(_03171_),
    .A(_03168_),
    .B(_03170_));
 sg13g2_a21oi_1 _17438_ (.A1(net4853),
    .A2(net4659),
    .Y(_03172_),
    .B1(_03169_));
 sg13g2_o21ai_1 _17439_ (.B1(_03168_),
    .Y(_03173_),
    .A1(net4728),
    .A2(_03172_));
 sg13g2_a22oi_1 _17440_ (.Y(_03174_),
    .B1(_03173_),
    .B2(_02974_),
    .A2(_03171_),
    .A1(_02953_));
 sg13g2_nand2b_1 _17441_ (.Y(_03175_),
    .B(net4806),
    .A_N(_03174_));
 sg13g2_nand2_1 _17442_ (.Y(_03176_),
    .A(net4820),
    .B(_03050_));
 sg13g2_a21oi_1 _17443_ (.A1(net4725),
    .A2(_03043_),
    .Y(_03177_),
    .B1(net4815));
 sg13g2_mux2_1 _17444_ (.A0(_03026_),
    .A1(_03048_),
    .S(net4719),
    .X(_03178_));
 sg13g2_nor2_1 _17445_ (.A(net4730),
    .B(_03178_),
    .Y(_03179_));
 sg13g2_a21oi_1 _17446_ (.A1(_03176_),
    .A2(_03177_),
    .Y(_03180_),
    .B1(_03179_));
 sg13g2_a22oi_1 _17447_ (.Y(_03181_),
    .B1(net4429),
    .B2(_02714_),
    .A2(net4439),
    .A1(_02711_));
 sg13g2_a21oi_1 _17448_ (.A1(_02713_),
    .A2(net4435),
    .Y(_03182_),
    .B1(net4880));
 sg13g2_nor2_1 _17449_ (.A(net4723),
    .B(_03060_),
    .Y(_03183_));
 sg13g2_a21oi_1 _17450_ (.A1(\soc_inst.cpu_core.alu.a[5] ),
    .A2(net4850),
    .Y(_03184_),
    .B1(_02916_));
 sg13g2_nand2_1 _17451_ (.Y(_03185_),
    .A(net4835),
    .B(_03126_));
 sg13g2_o21ai_1 _17452_ (.B1(_03185_),
    .Y(_03186_),
    .A1(net4835),
    .A2(_03184_));
 sg13g2_a21oi_1 _17453_ (.A1(net4723),
    .A2(_03186_),
    .Y(_03187_),
    .B1(_03183_));
 sg13g2_nor2_1 _17454_ (.A(net4811),
    .B(_03187_),
    .Y(_03188_));
 sg13g2_a22oi_1 _17455_ (.Y(_03189_),
    .B1(_03188_),
    .B2(net4212),
    .A2(_03180_),
    .A1(net4213));
 sg13g2_nand4_1 _17456_ (.B(_03181_),
    .C(_03182_),
    .A(_03175_),
    .Y(_03190_),
    .D(_03189_));
 sg13g2_a21oi_1 _17457_ (.A1(net4447),
    .A2(_03165_),
    .Y(_03191_),
    .B1(_03190_));
 sg13g2_a22oi_1 _17458_ (.Y(_01392_),
    .B1(_03164_),
    .B2(_03191_),
    .A2(_05762_),
    .A1(net4890));
 sg13g2_o21ai_1 _17459_ (.B1(net4447),
    .Y(_03192_),
    .A1(_02709_),
    .A2(_02744_));
 sg13g2_a21o_1 _17460_ (.A2(_02744_),
    .A1(_02709_),
    .B1(_03192_),
    .X(_03193_));
 sg13g2_a21o_2 _17461_ (.A2(_03162_),
    .A1(_02714_),
    .B1(_02713_),
    .X(_03194_));
 sg13g2_o21ai_1 _17462_ (.B1(net4426),
    .Y(_03195_),
    .A1(_02709_),
    .A2(_03194_));
 sg13g2_a21oi_1 _17463_ (.A1(_02709_),
    .A2(_03194_),
    .Y(_03196_),
    .B1(_03195_));
 sg13g2_nand2_1 _17464_ (.Y(_03197_),
    .A(net4821),
    .B(_03088_));
 sg13g2_a21oi_1 _17465_ (.A1(net4726),
    .A2(_03092_),
    .Y(_03198_),
    .B1(net4815));
 sg13g2_mux2_1 _17466_ (.A0(_03069_),
    .A1(_03086_),
    .S(net4718),
    .X(_03199_));
 sg13g2_nor2_1 _17467_ (.A(net4729),
    .B(_03199_),
    .Y(_03200_));
 sg13g2_a21oi_1 _17468_ (.A1(_03197_),
    .A2(_03198_),
    .Y(_03201_),
    .B1(_03200_));
 sg13g2_a21oi_1 _17469_ (.A1(\soc_inst.cpu_core.alu.a[6] ),
    .A2(net4850),
    .Y(_03202_),
    .B1(_02984_));
 sg13g2_nand2_1 _17470_ (.Y(_03203_),
    .A(net4837),
    .B(_03154_));
 sg13g2_o21ai_1 _17471_ (.B1(_03203_),
    .Y(_03204_),
    .A1(net4837),
    .A2(_03202_));
 sg13g2_mux2_1 _17472_ (.A0(_03098_),
    .A1(_03204_),
    .S(net4724),
    .X(_03205_));
 sg13g2_and2_1 _17473_ (.A(net4734),
    .B(_03205_),
    .X(_03206_));
 sg13g2_a221oi_1 _17474_ (.B2(_02709_),
    .C1(net4880),
    .B1(net4429),
    .A1(_02706_),
    .Y(_03207_),
    .A2(net4439));
 sg13g2_o21ai_1 _17475_ (.B1(_03207_),
    .Y(_03208_),
    .A1(_02707_),
    .A2(net4432));
 sg13g2_a221oi_1 _17476_ (.B2(net4211),
    .C1(_03208_),
    .B1(_03206_),
    .A1(net4213),
    .Y(_03209_),
    .A2(_03201_));
 sg13g2_mux2_1 _17477_ (.A0(_03068_),
    .A1(_03073_),
    .S(net4818),
    .X(_03210_));
 sg13g2_nor2_1 _17478_ (.A(net4808),
    .B(_03210_),
    .Y(_03211_));
 sg13g2_and2_1 _17479_ (.A(net4853),
    .B(_02974_),
    .X(_03212_));
 sg13g2_and2_1 _17480_ (.A(net4728),
    .B(_02974_),
    .X(_03213_));
 sg13g2_nor2_1 _17481_ (.A(_03212_),
    .B(_03213_),
    .Y(_03214_));
 sg13g2_nand2_1 _17482_ (.Y(_03215_),
    .A(_02924_),
    .B(_02967_));
 sg13g2_a21o_1 _17483_ (.A2(_03215_),
    .A1(net4809),
    .B1(_02954_),
    .X(_03216_));
 sg13g2_and2_1 _17484_ (.A(net4808),
    .B(_03212_),
    .X(_03217_));
 sg13g2_a21oi_2 _17485_ (.B1(_03211_),
    .Y(_03218_),
    .A2(_03216_),
    .A1(_03214_));
 sg13g2_a21oi_1 _17486_ (.A1(net4806),
    .A2(_03218_),
    .Y(_03219_),
    .B1(_03196_));
 sg13g2_and2_1 _17487_ (.A(_03209_),
    .B(_03219_),
    .X(_03220_));
 sg13g2_a22oi_1 _17488_ (.Y(_01393_),
    .B1(_03193_),
    .B2(_03220_),
    .A2(_05764_),
    .A1(net4886));
 sg13g2_a21o_2 _17489_ (.A2(_03194_),
    .A1(_02709_),
    .B1(_02708_),
    .X(_03221_));
 sg13g2_nand2b_1 _17490_ (.Y(_03222_),
    .B(_02749_),
    .A_N(_03221_));
 sg13g2_nand2_1 _17491_ (.Y(_03223_),
    .A(_02748_),
    .B(_03221_));
 sg13g2_nand3_1 _17492_ (.B(_03222_),
    .C(_03223_),
    .A(net4427),
    .Y(_03224_));
 sg13g2_nor2_1 _17493_ (.A(net4445),
    .B(_02751_),
    .Y(_03225_));
 sg13g2_o21ai_1 _17494_ (.B1(_03225_),
    .Y(_03226_),
    .A1(_02745_),
    .A2(_02749_));
 sg13g2_nor2_1 _17495_ (.A(net4733),
    .B(_02945_),
    .Y(_03227_));
 sg13g2_nand2_1 _17496_ (.Y(_03228_),
    .A(_02902_),
    .B(_02917_));
 sg13g2_nor2_1 _17497_ (.A(net4836),
    .B(_03228_),
    .Y(_03229_));
 sg13g2_a21oi_1 _17498_ (.A1(net4835),
    .A2(_03184_),
    .Y(_03230_),
    .B1(_03229_));
 sg13g2_mux2_1 _17499_ (.A0(_03127_),
    .A1(_03230_),
    .S(net4723),
    .X(_03231_));
 sg13g2_a22oi_1 _17500_ (.Y(_03232_),
    .B1(_03231_),
    .B2(net4210),
    .A2(net4209),
    .A1(_02928_));
 sg13g2_a21oi_1 _17501_ (.A1(net4811),
    .A2(_02880_),
    .Y(_03233_),
    .B1(_02669_));
 sg13g2_o21ai_1 _17502_ (.B1(_03233_),
    .Y(_03234_),
    .A1(net4812),
    .A2(_02909_));
 sg13g2_a21oi_1 _17503_ (.A1(_03232_),
    .A2(_03234_),
    .Y(_03235_),
    .B1(net4806));
 sg13g2_a21oi_1 _17504_ (.A1(net4730),
    .A2(_02892_),
    .Y(_03236_),
    .B1(_03217_));
 sg13g2_nor3_1 _17505_ (.A(net4735),
    .B(_02669_),
    .C(_03236_),
    .Y(_03237_));
 sg13g2_a22oi_1 _17506_ (.Y(_03238_),
    .B1(net4430),
    .B2(_02748_),
    .A2(net4440),
    .A1(_02746_));
 sg13g2_o21ai_1 _17507_ (.B1(_03238_),
    .Y(_03239_),
    .A1(_02747_),
    .A2(net4433));
 sg13g2_nor4_1 _17508_ (.A(net4881),
    .B(_03235_),
    .C(_03237_),
    .D(_03239_),
    .Y(_03240_));
 sg13g2_and2_1 _17509_ (.A(_03224_),
    .B(_03240_),
    .X(_03241_));
 sg13g2_a22oi_1 _17510_ (.Y(_01394_),
    .B1(_03226_),
    .B2(_03241_),
    .A2(_05765_),
    .A1(net4886));
 sg13g2_nand3_1 _17511_ (.B(_02747_),
    .C(_03223_),
    .A(_02701_),
    .Y(_03242_));
 sg13g2_nor2_1 _17512_ (.A(_02701_),
    .B(_02749_),
    .Y(_03243_));
 sg13g2_nand2_1 _17513_ (.Y(_03244_),
    .A(_03221_),
    .B(_03243_));
 sg13g2_or2_1 _17514_ (.X(_03245_),
    .B(_02747_),
    .A(_02701_));
 sg13g2_nand4_1 _17515_ (.B(_03242_),
    .C(_03244_),
    .A(net4427),
    .Y(_03246_),
    .D(_03245_));
 sg13g2_nand3_1 _17516_ (.B(_02702_),
    .C(_02750_),
    .A(_02700_),
    .Y(_03247_));
 sg13g2_nand4_1 _17517_ (.B(_02703_),
    .C(_02752_),
    .A(_02670_),
    .Y(_03248_),
    .D(_03247_));
 sg13g2_o21ai_1 _17518_ (.B1(_02999_),
    .Y(_03249_),
    .A1(_05824_),
    .A2(_05839_));
 sg13g2_nor2_1 _17519_ (.A(net4836),
    .B(_03249_),
    .Y(_03250_));
 sg13g2_a21oi_1 _17520_ (.A1(net4835),
    .A2(_03202_),
    .Y(_03251_),
    .B1(_03250_));
 sg13g2_mux2_1 _17521_ (.A0(_03156_),
    .A1(_03251_),
    .S(net4724),
    .X(_03252_));
 sg13g2_nor2_1 _17522_ (.A(net4814),
    .B(_03252_),
    .Y(_03253_));
 sg13g2_a21oi_1 _17523_ (.A1(_02924_),
    .A2(_03018_),
    .Y(_03254_),
    .B1(net4734));
 sg13g2_nor2_1 _17524_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sg13g2_mux2_1 _17525_ (.A0(_02961_),
    .A1(_03005_),
    .S(net4732),
    .X(_03256_));
 sg13g2_a221oi_1 _17526_ (.B2(_02700_),
    .C1(net4880),
    .B1(net4429),
    .A1(_02698_),
    .Y(_03257_),
    .A2(net4439));
 sg13g2_o21ai_1 _17527_ (.B1(_03257_),
    .Y(_03258_),
    .A1(_02699_),
    .A2(net4432));
 sg13g2_nand2b_1 _17528_ (.Y(_03259_),
    .B(_03213_),
    .A_N(_02977_));
 sg13g2_nor2_2 _17529_ (.A(net4808),
    .B(_02954_),
    .Y(_03260_));
 sg13g2_nand2b_1 _17530_ (.Y(_03261_),
    .B(_03260_),
    .A_N(_02972_));
 sg13g2_nand3b_1 _17531_ (.B(_03259_),
    .C(_03261_),
    .Y(_03262_),
    .A_N(_03217_));
 sg13g2_a221oi_1 _17532_ (.B2(net4806),
    .C1(_03258_),
    .B1(_03262_),
    .A1(net4211),
    .Y(_03263_),
    .A2(_03255_));
 sg13g2_nand2_1 _17533_ (.Y(_03264_),
    .A(_03248_),
    .B(_03263_));
 sg13g2_a21oi_1 _17534_ (.A1(net4213),
    .A2(_03256_),
    .Y(_03265_),
    .B1(_03264_));
 sg13g2_a22oi_1 _17535_ (.Y(_01395_),
    .B1(_03246_),
    .B2(_03265_),
    .A2(_05766_),
    .A1(net4886));
 sg13g2_nand2_1 _17536_ (.Y(_03266_),
    .A(_02699_),
    .B(_03245_));
 sg13g2_a21oi_1 _17537_ (.A1(_03221_),
    .A2(_03243_),
    .Y(_03267_),
    .B1(_03266_));
 sg13g2_nand2b_1 _17538_ (.Y(_03268_),
    .B(_02695_),
    .A_N(_03267_));
 sg13g2_a21oi_1 _17539_ (.A1(_02696_),
    .A2(_03267_),
    .Y(_03269_),
    .B1(_03015_));
 sg13g2_nor2_1 _17540_ (.A(_02695_),
    .B(_02753_),
    .Y(_03270_));
 sg13g2_xnor2_1 _17541_ (.Y(_03271_),
    .A(_02696_),
    .B(_02753_));
 sg13g2_nor2_1 _17542_ (.A(net4811),
    .B(_03051_),
    .Y(_03272_));
 sg13g2_o21ai_1 _17543_ (.B1(net4213),
    .Y(_03273_),
    .A1(net4730),
    .A2(_03029_));
 sg13g2_a21o_1 _17544_ (.A2(net4849),
    .A1(\soc_inst.cpu_core.alu.a[9] ),
    .B1(_02905_),
    .X(_03274_));
 sg13g2_mux2_1 _17545_ (.A0(_03274_),
    .A1(_03228_),
    .S(net4835),
    .X(_03275_));
 sg13g2_mux2_1 _17546_ (.A0(_03186_),
    .A1(_03275_),
    .S(net4722),
    .X(_03276_));
 sg13g2_nor2_1 _17547_ (.A(net4812),
    .B(_03276_),
    .Y(_03277_));
 sg13g2_a21oi_1 _17548_ (.A1(net4812),
    .A2(_03061_),
    .Y(_03278_),
    .B1(_03277_));
 sg13g2_a221oi_1 _17549_ (.B2(_02695_),
    .C1(net4886),
    .B1(net4430),
    .A1(_02693_),
    .Y(_03279_),
    .A2(net4440));
 sg13g2_o21ai_1 _17550_ (.B1(_03279_),
    .Y(_03280_),
    .A1(_02694_),
    .A2(net4433));
 sg13g2_a221oi_1 _17551_ (.B2(_03035_),
    .C1(_03217_),
    .B1(_03260_),
    .A1(_03037_),
    .Y(_03281_),
    .A2(_03213_));
 sg13g2_inv_1 _17552_ (.Y(_03282_),
    .A(_03281_));
 sg13g2_a221oi_1 _17553_ (.B2(net4803),
    .C1(_03280_),
    .B1(_03282_),
    .A1(net4212),
    .Y(_03283_),
    .A2(_03278_));
 sg13g2_o21ai_1 _17554_ (.B1(_03283_),
    .Y(_03284_),
    .A1(_03272_),
    .A2(_03273_));
 sg13g2_a221oi_1 _17555_ (.B2(net4447),
    .C1(_03284_),
    .B1(_03271_),
    .A1(_03268_),
    .Y(_03285_),
    .A2(_03269_));
 sg13g2_a21oi_1 _17556_ (.A1(net4907),
    .A2(_05767_),
    .Y(_01396_),
    .B1(_03285_));
 sg13g2_nor2_1 _17557_ (.A(_02755_),
    .B(_03270_),
    .Y(_03286_));
 sg13g2_xor2_1 _17558_ (.B(_03286_),
    .A(_02691_),
    .X(_03287_));
 sg13g2_nand2_1 _17559_ (.Y(_03288_),
    .A(_02694_),
    .B(_03268_));
 sg13g2_a21oi_1 _17560_ (.A1(_02691_),
    .A2(_03288_),
    .Y(_03289_),
    .B1(_03015_));
 sg13g2_o21ai_1 _17561_ (.B1(_03289_),
    .Y(_03290_),
    .A1(_02691_),
    .A2(_03288_));
 sg13g2_a221oi_1 _17562_ (.B2(_03075_),
    .C1(_03217_),
    .B1(_03260_),
    .A1(_03079_),
    .Y(_03291_),
    .A2(_03213_));
 sg13g2_nor2_1 _17563_ (.A(net4729),
    .B(_03070_),
    .Y(_03292_));
 sg13g2_a21oi_1 _17564_ (.A1(net4732),
    .A2(_03090_),
    .Y(_03293_),
    .B1(_03292_));
 sg13g2_a21o_1 _17565_ (.A2(net4851),
    .A1(\soc_inst.cpu_core.alu.a[10] ),
    .B1(_03002_),
    .X(_03294_));
 sg13g2_mux2_1 _17566_ (.A0(_03294_),
    .A1(_03249_),
    .S(net4838),
    .X(_03295_));
 sg13g2_mux2_1 _17567_ (.A0(_03204_),
    .A1(_03295_),
    .S(net4724),
    .X(_03296_));
 sg13g2_nor2_1 _17568_ (.A(net4814),
    .B(_03296_),
    .Y(_03297_));
 sg13g2_a21oi_1 _17569_ (.A1(net4814),
    .A2(_03099_),
    .Y(_03298_),
    .B1(_03297_));
 sg13g2_a221oi_1 _17570_ (.B2(_02691_),
    .C1(net4886),
    .B1(net4430),
    .A1(_02689_),
    .Y(_03299_),
    .A2(net4440));
 sg13g2_o21ai_1 _17571_ (.B1(_03299_),
    .Y(_03300_),
    .A1(_02690_),
    .A2(net4433));
 sg13g2_a221oi_1 _17572_ (.B2(net4211),
    .C1(_03300_),
    .B1(_03298_),
    .A1(net4214),
    .Y(_03301_),
    .A2(_03293_));
 sg13g2_o21ai_1 _17573_ (.B1(_03301_),
    .Y(_03302_),
    .A1(net4736),
    .A2(_03291_));
 sg13g2_a21oi_1 _17574_ (.A1(net4447),
    .A2(_03287_),
    .Y(_03303_),
    .B1(_03302_));
 sg13g2_a22oi_1 _17575_ (.Y(_01397_),
    .B1(_03290_),
    .B2(_03303_),
    .A2(_05768_),
    .A1(net4886));
 sg13g2_a21oi_1 _17576_ (.A1(_02690_),
    .A2(_02692_),
    .Y(_03304_),
    .B1(_02688_));
 sg13g2_nand2_1 _17577_ (.Y(_03305_),
    .A(_02690_),
    .B(_02694_));
 sg13g2_a221oi_1 _17578_ (.B2(_02689_),
    .C1(_03266_),
    .B1(_03305_),
    .A1(_03221_),
    .Y(_03306_),
    .A2(_03243_));
 sg13g2_nand2b_1 _17579_ (.Y(_03307_),
    .B(_03304_),
    .A_N(_03306_));
 sg13g2_or2_1 _17580_ (.X(_03308_),
    .B(_03307_),
    .A(_02761_));
 sg13g2_a21oi_1 _17581_ (.A1(_02761_),
    .A2(_03307_),
    .Y(_03309_),
    .B1(net4424));
 sg13g2_mux2_1 _17582_ (.A0(\soc_inst.cpu_core.alu.a[12] ),
    .A1(\soc_inst.cpu_core.alu.a[11] ),
    .S(net4851),
    .X(_03310_));
 sg13g2_mux2_1 _17583_ (.A0(_03310_),
    .A1(_03274_),
    .S(net4830),
    .X(_03311_));
 sg13g2_mux2_1 _17584_ (.A0(_03230_),
    .A1(_03311_),
    .S(net4723),
    .X(_03312_));
 sg13g2_nor2_1 _17585_ (.A(net4811),
    .B(_03312_),
    .Y(_03313_));
 sg13g2_a21oi_1 _17586_ (.A1(net4811),
    .A2(_03128_),
    .Y(_03314_),
    .B1(_03313_));
 sg13g2_o21ai_1 _17587_ (.B1(net4213),
    .Y(_03315_),
    .A1(net4813),
    .A2(_03121_));
 sg13g2_a21oi_1 _17588_ (.A1(net4813),
    .A2(_03113_),
    .Y(_03316_),
    .B1(_03315_));
 sg13g2_a21oi_1 _17589_ (.A1(net4212),
    .A2(_03314_),
    .Y(_03317_),
    .B1(_03316_));
 sg13g2_a221oi_1 _17590_ (.B2(_03115_),
    .C1(_03217_),
    .B1(_03260_),
    .A1(_03117_),
    .Y(_03318_),
    .A2(_03213_));
 sg13g2_o21ai_1 _17591_ (.B1(net4438),
    .Y(_03319_),
    .A1(net1895),
    .A2(\soc_inst.cpu_core.alu.a[12] ));
 sg13g2_nor2_1 _17592_ (.A(_02760_),
    .B(net4432),
    .Y(_03320_));
 sg13g2_o21ai_1 _17593_ (.B1(_03319_),
    .Y(_03321_),
    .A1(_02761_),
    .A2(_03011_));
 sg13g2_o21ai_1 _17594_ (.B1(_03317_),
    .Y(_03322_),
    .A1(net4735),
    .A2(_03318_));
 sg13g2_nor4_1 _17595_ (.A(net4883),
    .B(_03320_),
    .C(_03321_),
    .D(_03322_),
    .Y(_03323_));
 sg13g2_nor2_1 _17596_ (.A(_02759_),
    .B(_02761_),
    .Y(_03324_));
 sg13g2_nor2_1 _17597_ (.A(net4444),
    .B(_03324_),
    .Y(_03325_));
 sg13g2_a22oi_1 _17598_ (.Y(_03326_),
    .B1(_03325_),
    .B2(_02762_),
    .A2(_03309_),
    .A1(_03308_));
 sg13g2_a22oi_1 _17599_ (.Y(_01398_),
    .B1(_03323_),
    .B2(_03326_),
    .A2(_05769_),
    .A1(net4884));
 sg13g2_nor2_1 _17600_ (.A(_02687_),
    .B(_03308_),
    .Y(_03327_));
 sg13g2_nor2_1 _17601_ (.A(_02687_),
    .B(_02760_),
    .Y(_03328_));
 sg13g2_and3_1 _17602_ (.X(_03329_),
    .A(_02687_),
    .B(_02760_),
    .C(_03308_));
 sg13g2_nor4_1 _17603_ (.A(net4424),
    .B(_03327_),
    .C(_03328_),
    .D(_03329_),
    .Y(_03330_));
 sg13g2_nand3_1 _17604_ (.B(_02762_),
    .C(_02764_),
    .A(_02686_),
    .Y(_03331_));
 sg13g2_nand4_1 _17605_ (.B(_02763_),
    .C(_02766_),
    .A(net4446),
    .Y(_03332_),
    .D(_03331_));
 sg13g2_mux2_1 _17606_ (.A0(\soc_inst.cpu_core.alu.a[13] ),
    .A1(\soc_inst.cpu_core.alu.a[12] ),
    .S(net4847),
    .X(_03333_));
 sg13g2_mux2_1 _17607_ (.A0(_03333_),
    .A1(_03294_),
    .S(net4832),
    .X(_03334_));
 sg13g2_mux2_1 _17608_ (.A0(_03251_),
    .A1(_03334_),
    .S(net4723),
    .X(_03335_));
 sg13g2_nand2_1 _17609_ (.Y(_03336_),
    .A(net4812),
    .B(_03157_));
 sg13g2_o21ai_1 _17610_ (.B1(_03336_),
    .Y(_03337_),
    .A1(net4812),
    .A2(_03335_));
 sg13g2_nor2_1 _17611_ (.A(_02947_),
    .B(_03337_),
    .Y(_03338_));
 sg13g2_a221oi_1 _17612_ (.B2(_03140_),
    .C1(_03217_),
    .B1(_03260_),
    .A1(_03143_),
    .Y(_03339_),
    .A2(_03213_));
 sg13g2_nand2b_1 _17613_ (.Y(_03340_),
    .B(net4802),
    .A_N(_03339_));
 sg13g2_o21ai_1 _17614_ (.B1(net4437),
    .Y(_03341_),
    .A1(net2621),
    .A2(net4863));
 sg13g2_nand3_1 _17615_ (.B(net4863),
    .C(net4434),
    .A(net2621),
    .Y(_03342_));
 sg13g2_a21oi_1 _17616_ (.A1(_02686_),
    .A2(net4428),
    .Y(_03343_),
    .B1(net4883));
 sg13g2_nand4_1 _17617_ (.B(_03341_),
    .C(_03342_),
    .A(_03340_),
    .Y(_03344_),
    .D(_03343_));
 sg13g2_o21ai_1 _17618_ (.B1(net4213),
    .Y(_03345_),
    .A1(net4729),
    .A2(_03138_));
 sg13g2_a21oi_1 _17619_ (.A1(net4731),
    .A2(_03148_),
    .Y(_03346_),
    .B1(_03345_));
 sg13g2_nor4_1 _17620_ (.A(_03330_),
    .B(_03338_),
    .C(_03344_),
    .D(_03346_),
    .Y(_03347_));
 sg13g2_a22oi_1 _17621_ (.Y(_01399_),
    .B1(_03332_),
    .B2(_03347_),
    .A2(_05770_),
    .A1(net4884));
 sg13g2_and2_1 _17622_ (.A(_02763_),
    .B(_02767_),
    .X(_03348_));
 sg13g2_xnor2_1 _17623_ (.Y(_03349_),
    .A(_02684_),
    .B(_03348_));
 sg13g2_o21ai_1 _17624_ (.B1(_02896_),
    .Y(_03350_),
    .A1(_05812_),
    .A2(net4846));
 sg13g2_mux2_1 _17625_ (.A0(_03350_),
    .A1(_03310_),
    .S(net4832),
    .X(_03351_));
 sg13g2_mux2_1 _17626_ (.A0(_03275_),
    .A1(_03351_),
    .S(net4722),
    .X(_03352_));
 sg13g2_nor2_1 _17627_ (.A(net4813),
    .B(_03352_),
    .Y(_03353_));
 sg13g2_a21oi_1 _17628_ (.A1(net4811),
    .A2(_03187_),
    .Y(_03354_),
    .B1(_03353_));
 sg13g2_a21oi_1 _17629_ (.A1(net4728),
    .A2(_03172_),
    .Y(_03355_),
    .B1(_03214_));
 sg13g2_a21o_2 _17630_ (.A2(_03260_),
    .A1(_03169_),
    .B1(_03355_),
    .X(_03356_));
 sg13g2_a22oi_1 _17631_ (.Y(_03357_),
    .B1(net4431),
    .B2(_02683_),
    .A2(net4437),
    .A1(_02682_));
 sg13g2_a21oi_1 _17632_ (.A1(_02681_),
    .A2(net4434),
    .Y(_03358_),
    .B1(net4883));
 sg13g2_a21oi_1 _17633_ (.A1(net4809),
    .A2(_03167_),
    .Y(_03359_),
    .B1(_02911_));
 sg13g2_o21ai_1 _17634_ (.B1(_03359_),
    .Y(_03360_),
    .A1(net4809),
    .A2(_03178_));
 sg13g2_a22oi_1 _17635_ (.Y(_03361_),
    .B1(_03356_),
    .B2(net4802),
    .A2(_03354_),
    .A1(net4212));
 sg13g2_nand4_1 _17636_ (.B(_03358_),
    .C(_03360_),
    .A(_03357_),
    .Y(_03362_),
    .D(_03361_));
 sg13g2_a21o_1 _17637_ (.A2(net4863),
    .A1(\soc_inst.cpu_core.alu.b[13] ),
    .B1(_03328_),
    .X(_03363_));
 sg13g2_nor2_1 _17638_ (.A(_03327_),
    .B(_03363_),
    .Y(_03364_));
 sg13g2_nor2_1 _17639_ (.A(_02684_),
    .B(_03364_),
    .Y(_03365_));
 sg13g2_xnor2_1 _17640_ (.Y(_03366_),
    .A(_02683_),
    .B(_03364_));
 sg13g2_a221oi_1 _17641_ (.B2(net4427),
    .C1(_03362_),
    .B1(_03366_),
    .A1(net4446),
    .Y(_03367_),
    .A2(_03349_));
 sg13g2_a21oi_1 _17642_ (.A1(net4883),
    .A2(_05771_),
    .Y(_01400_),
    .B1(_03367_));
 sg13g2_o21ai_1 _17643_ (.B1(_02685_),
    .Y(_03368_),
    .A1(_02683_),
    .A2(_03348_));
 sg13g2_xnor2_1 _17644_ (.Y(_03369_),
    .A(_02679_),
    .B(_03368_));
 sg13g2_nor2_1 _17645_ (.A(_02681_),
    .B(_03365_),
    .Y(_03370_));
 sg13g2_a21oi_1 _17646_ (.A1(_02680_),
    .A2(_03370_),
    .Y(_03371_),
    .B1(net4424));
 sg13g2_o21ai_1 _17647_ (.B1(_03371_),
    .Y(_03372_),
    .A1(_02680_),
    .A2(_03370_));
 sg13g2_o21ai_1 _17648_ (.B1(_02994_),
    .Y(_03373_),
    .A1(_05810_),
    .A2(net4846));
 sg13g2_mux2_1 _17649_ (.A0(_03373_),
    .A1(_03333_),
    .S(net4830),
    .X(_03374_));
 sg13g2_mux2_1 _17650_ (.A0(_03295_),
    .A1(_03374_),
    .S(net4722),
    .X(_03375_));
 sg13g2_mux2_1 _17651_ (.A0(_03205_),
    .A1(_03375_),
    .S(net4733),
    .X(_03376_));
 sg13g2_mux2_1 _17652_ (.A0(_03199_),
    .A1(_03210_),
    .S(net4808),
    .X(_03377_));
 sg13g2_and2_1 _17653_ (.A(net4803),
    .B(_03212_),
    .X(_03378_));
 sg13g2_nand2_2 _17654_ (.Y(_03379_),
    .A(net4802),
    .B(_03212_));
 sg13g2_a22oi_1 _17655_ (.Y(_03380_),
    .B1(net4428),
    .B2(_02679_),
    .A2(net4438),
    .A1(_02677_));
 sg13g2_a21oi_1 _17656_ (.A1(_02678_),
    .A2(net4434),
    .Y(_03381_),
    .B1(net4883));
 sg13g2_nor3_2 _17657_ (.A(net4808),
    .B(_02954_),
    .C(_03215_),
    .Y(_03382_));
 sg13g2_a22oi_1 _17658_ (.Y(_03383_),
    .B1(_03382_),
    .B2(net4804),
    .A2(_03376_),
    .A1(net4212));
 sg13g2_nand4_1 _17659_ (.B(_03380_),
    .C(_03381_),
    .A(_03379_),
    .Y(_03384_),
    .D(_03383_));
 sg13g2_a221oi_1 _17660_ (.B2(net4214),
    .C1(_03384_),
    .B1(_03377_),
    .A1(net4446),
    .Y(_03385_),
    .A2(_03369_));
 sg13g2_a22oi_1 _17661_ (.Y(_01401_),
    .B1(_03372_),
    .B2(_03385_),
    .A2(_05772_),
    .A1(net4883));
 sg13g2_nor4_1 _17662_ (.A(_02680_),
    .B(_02684_),
    .C(_02687_),
    .D(_02761_),
    .Y(_03386_));
 sg13g2_nand3b_1 _17663_ (.B(_03386_),
    .C(_03304_),
    .Y(_03387_),
    .A_N(_03306_));
 sg13g2_nand3_1 _17664_ (.B(_02683_),
    .C(_03363_),
    .A(_02679_),
    .Y(_03388_));
 sg13g2_a21oi_1 _17665_ (.A1(_02677_),
    .A2(_02681_),
    .Y(_03389_),
    .B1(_02678_));
 sg13g2_nand2_1 _17666_ (.Y(_03390_),
    .A(_03388_),
    .B(_03389_));
 sg13g2_inv_1 _17667_ (.Y(_03391_),
    .A(_03390_));
 sg13g2_and2_1 _17668_ (.A(_03387_),
    .B(_03391_),
    .X(_03392_));
 sg13g2_nor2b_1 _17669_ (.A(_03392_),
    .B_N(net4443),
    .Y(_03393_));
 sg13g2_xnor2_1 _17670_ (.Y(_03394_),
    .A(net4443),
    .B(_03392_));
 sg13g2_or2_1 _17671_ (.X(_03395_),
    .B(net4443),
    .A(_02771_));
 sg13g2_a21oi_1 _17672_ (.A1(_02771_),
    .A2(net4443),
    .Y(_03396_),
    .B1(net4444));
 sg13g2_mux2_1 _17673_ (.A0(\soc_inst.cpu_core.alu.a[16] ),
    .A1(\soc_inst.cpu_core.alu.a[15] ),
    .S(net4846),
    .X(_03397_));
 sg13g2_mux2_1 _17674_ (.A0(_03397_),
    .A1(_03350_),
    .S(net4831),
    .X(_03398_));
 sg13g2_and2_1 _17675_ (.A(net4721),
    .B(_03398_),
    .X(_03399_));
 sg13g2_a21oi_1 _17676_ (.A1(net4820),
    .A2(_03311_),
    .Y(_03400_),
    .B1(_03399_));
 sg13g2_a21oi_1 _17677_ (.A1(net4733),
    .A2(_03400_),
    .Y(_03401_),
    .B1(_02947_));
 sg13g2_o21ai_1 _17678_ (.B1(_03401_),
    .Y(_03402_),
    .A1(net4733),
    .A2(_03231_));
 sg13g2_nor2_1 _17679_ (.A(_02776_),
    .B(net4432),
    .Y(_03403_));
 sg13g2_a21oi_1 _17680_ (.A1(_02777_),
    .A2(net4431),
    .Y(_03404_),
    .B1(_03403_));
 sg13g2_o21ai_1 _17681_ (.B1(_03404_),
    .Y(_03405_),
    .A1(_02775_),
    .A2(_02936_));
 sg13g2_nor2_2 _17682_ (.A(net4736),
    .B(_02945_),
    .Y(_03406_));
 sg13g2_nand2_1 _17683_ (.Y(_03407_),
    .A(net4805),
    .B(_02944_));
 sg13g2_nand2b_1 _17684_ (.Y(_03408_),
    .B(net4067),
    .A_N(_03405_));
 sg13g2_a221oi_1 _17685_ (.B2(net4208),
    .C1(_03408_),
    .B1(_02943_),
    .A1(_02894_),
    .Y(_03409_),
    .A2(net4214));
 sg13g2_nand2_1 _17686_ (.Y(_03410_),
    .A(_03402_),
    .B(_03409_));
 sg13g2_a221oi_1 _17687_ (.B2(_03396_),
    .C1(_03410_),
    .B1(_03395_),
    .A1(net4425),
    .Y(_03411_),
    .A2(_03394_));
 sg13g2_nand2_1 _17688_ (.Y(_03412_),
    .A(net4917),
    .B(net1109));
 sg13g2_o21ai_1 _17689_ (.B1(_03412_),
    .Y(_01402_),
    .A1(net4111),
    .A2(_03411_));
 sg13g2_nand2_1 _17690_ (.Y(_03413_),
    .A(net4914),
    .B(net1996));
 sg13g2_o21ai_1 _17691_ (.B1(_02776_),
    .Y(_03414_),
    .A1(_02775_),
    .A2(_03392_));
 sg13g2_xor2_1 _17692_ (.B(_03414_),
    .A(net4215),
    .X(_03415_));
 sg13g2_nand3_1 _17693_ (.B(_02808_),
    .C(_03395_),
    .A(net4215),
    .Y(_03416_));
 sg13g2_o21ai_1 _17694_ (.B1(net4447),
    .Y(_03417_),
    .A1(net4215),
    .A2(_02808_));
 sg13g2_nor2_1 _17695_ (.A(_02778_),
    .B(_03417_),
    .Y(_03418_));
 sg13g2_o21ai_1 _17696_ (.B1(_02996_),
    .Y(_03419_),
    .A1(_05806_),
    .A2(net4845));
 sg13g2_mux2_1 _17697_ (.A0(_03419_),
    .A1(_03373_),
    .S(net4830),
    .X(_03420_));
 sg13g2_mux2_1 _17698_ (.A0(_03334_),
    .A1(_03420_),
    .S(net4722),
    .X(_03421_));
 sg13g2_a22oi_1 _17699_ (.Y(_03422_),
    .B1(_03421_),
    .B2(_03017_),
    .A2(_03252_),
    .A1(net4209));
 sg13g2_a21o_1 _17700_ (.A2(_03422_),
    .A1(_02979_),
    .B1(net4804),
    .X(_03423_));
 sg13g2_nor2_1 _17701_ (.A(_02773_),
    .B(net4432),
    .Y(_03424_));
 sg13g2_a221oi_1 _17702_ (.B2(net4215),
    .C1(_03424_),
    .B1(net4428),
    .A1(_02772_),
    .Y(_03425_),
    .A2(net4438));
 sg13g2_or2_1 _17703_ (.X(_03426_),
    .B(_03019_),
    .A(net4736));
 sg13g2_nand4_1 _17704_ (.B(_03423_),
    .C(_03425_),
    .A(net4067),
    .Y(_03427_),
    .D(_03426_));
 sg13g2_a221oi_1 _17705_ (.B2(_03418_),
    .C1(_03427_),
    .B1(_03416_),
    .A1(net4425),
    .Y(_03428_),
    .A2(_03415_));
 sg13g2_o21ai_1 _17706_ (.B1(_03413_),
    .Y(_01403_),
    .A1(net4111),
    .A2(_03428_));
 sg13g2_nand2_1 _17707_ (.Y(_03429_),
    .A(_02773_),
    .B(_02776_));
 sg13g2_nand2_1 _17708_ (.Y(_03430_),
    .A(_02772_),
    .B(_03429_));
 sg13g2_o21ai_1 _17709_ (.B1(_02772_),
    .Y(_03431_),
    .A1(_03393_),
    .A2(_03429_));
 sg13g2_or2_1 _17710_ (.X(_03432_),
    .B(_03431_),
    .A(_02799_));
 sg13g2_a21oi_1 _17711_ (.A1(_02799_),
    .A2(_03431_),
    .Y(_03433_),
    .B1(net4424));
 sg13g2_nor2_1 _17712_ (.A(_02778_),
    .B(_02810_),
    .Y(_03434_));
 sg13g2_nor2_1 _17713_ (.A(_02798_),
    .B(_03434_),
    .Y(_03435_));
 sg13g2_xnor2_1 _17714_ (.Y(_03436_),
    .A(_02799_),
    .B(_03434_));
 sg13g2_mux2_1 _17715_ (.A0(net4862),
    .A1(\soc_inst.cpu_core.alu.a[17] ),
    .S(net4845),
    .X(_03437_));
 sg13g2_mux2_1 _17716_ (.A0(_03437_),
    .A1(_03397_),
    .S(net4831),
    .X(_03438_));
 sg13g2_mux2_1 _17717_ (.A0(_03351_),
    .A1(_03438_),
    .S(net4721),
    .X(_03439_));
 sg13g2_a22oi_1 _17718_ (.Y(_03440_),
    .B1(_03439_),
    .B2(net4210),
    .A2(_03276_),
    .A1(net4209));
 sg13g2_a21oi_1 _17719_ (.A1(_03040_),
    .A2(_03440_),
    .Y(_03441_),
    .B1(net4804));
 sg13g2_o21ai_1 _17720_ (.B1(net4438),
    .Y(_03442_),
    .A1(\soc_inst.cpu_core.alu.b[18] ),
    .A2(\soc_inst.cpu_core.alu.a[18] ));
 sg13g2_o21ai_1 _17721_ (.B1(_03442_),
    .Y(_03443_),
    .A1(_02797_),
    .A2(net4432));
 sg13g2_nand2b_1 _17722_ (.Y(_03444_),
    .B(_03379_),
    .A_N(_03443_));
 sg13g2_a221oi_1 _17723_ (.B2(net4208),
    .C1(_03444_),
    .B1(_03062_),
    .A1(_02798_),
    .Y(_03445_),
    .A2(net4428));
 sg13g2_nand2b_1 _17724_ (.Y(_03446_),
    .B(_03445_),
    .A_N(_03441_));
 sg13g2_a221oi_1 _17725_ (.B2(net4446),
    .C1(_03446_),
    .B1(_03436_),
    .A1(_03432_),
    .Y(_03447_),
    .A2(_03433_));
 sg13g2_nand2_1 _17726_ (.Y(_03448_),
    .A(net4914),
    .B(net1128));
 sg13g2_o21ai_1 _17727_ (.B1(_03448_),
    .Y(_01404_),
    .A1(net4111),
    .A2(_03447_));
 sg13g2_a21oi_1 _17728_ (.A1(_02797_),
    .A2(_03432_),
    .Y(_03449_),
    .B1(_02796_));
 sg13g2_nand3_1 _17729_ (.B(_02797_),
    .C(_03432_),
    .A(_02796_),
    .Y(_03450_));
 sg13g2_nor2_1 _17730_ (.A(net4424),
    .B(_03449_),
    .Y(_03451_));
 sg13g2_nor3_1 _17731_ (.A(_02796_),
    .B(_02807_),
    .C(_03435_),
    .Y(_03452_));
 sg13g2_o21ai_1 _17732_ (.B1(_02796_),
    .Y(_03453_),
    .A1(_02807_),
    .A2(_03435_));
 sg13g2_nor2_1 _17733_ (.A(net4444),
    .B(_03452_),
    .Y(_03454_));
 sg13g2_o21ai_1 _17734_ (.B1(_02956_),
    .Y(_03455_),
    .A1(_05802_),
    .A2(net4845));
 sg13g2_mux2_1 _17735_ (.A0(_03455_),
    .A1(_03419_),
    .S(net4831),
    .X(_03456_));
 sg13g2_mux2_1 _17736_ (.A0(_03374_),
    .A1(_03456_),
    .S(net4727),
    .X(_03457_));
 sg13g2_a22oi_1 _17737_ (.Y(_03458_),
    .B1(_03457_),
    .B2(_03017_),
    .A2(_03296_),
    .A1(_03227_));
 sg13g2_a21oi_1 _17738_ (.A1(_03081_),
    .A2(_03458_),
    .Y(_03459_),
    .B1(net4804));
 sg13g2_nor3_1 _17739_ (.A(net4812),
    .B(_03099_),
    .C(_03407_),
    .Y(_03460_));
 sg13g2_nand3_1 _17740_ (.B(\soc_inst.cpu_core.alu.a[19] ),
    .C(net4434),
    .A(\soc_inst.cpu_core.alu.b[19] ),
    .Y(_03461_));
 sg13g2_o21ai_1 _17741_ (.B1(_03461_),
    .Y(_03462_),
    .A1(_02794_),
    .A2(_02936_));
 sg13g2_nor4_1 _17742_ (.A(_03378_),
    .B(_03459_),
    .C(_03460_),
    .D(_03462_),
    .Y(_03463_));
 sg13g2_o21ai_1 _17743_ (.B1(_03463_),
    .Y(_03464_),
    .A1(_02796_),
    .A2(_03011_));
 sg13g2_a221oi_1 _17744_ (.B2(_03454_),
    .C1(_03464_),
    .B1(_03453_),
    .A1(_03450_),
    .Y(_03465_),
    .A2(_03451_));
 sg13g2_nand2_1 _17745_ (.Y(_03466_),
    .A(net4913),
    .B(net898));
 sg13g2_o21ai_1 _17746_ (.B1(_03466_),
    .Y(_01405_),
    .A1(net4111),
    .A2(_03465_));
 sg13g2_nor4_1 _17747_ (.A(_02771_),
    .B(net4215),
    .C(net4443),
    .D(_02800_),
    .Y(_03467_));
 sg13g2_o21ai_1 _17748_ (.B1(_02793_),
    .Y(_03468_),
    .A1(_02814_),
    .A2(_03467_));
 sg13g2_nor3_1 _17749_ (.A(_02793_),
    .B(_02814_),
    .C(_03467_),
    .Y(_03469_));
 sg13g2_nor2_1 _17750_ (.A(net4444),
    .B(_03469_),
    .Y(_03470_));
 sg13g2_nand2_1 _17751_ (.Y(_03471_),
    .A(_02795_),
    .B(_02798_));
 sg13g2_nand4_1 _17752_ (.B(net4443),
    .C(_02795_),
    .A(_02774_),
    .Y(_03472_),
    .D(_02798_));
 sg13g2_a21oi_1 _17753_ (.A1(_03387_),
    .A2(_03391_),
    .Y(_03473_),
    .B1(_03472_));
 sg13g2_nor2_1 _17754_ (.A(_02794_),
    .B(_02797_),
    .Y(_03474_));
 sg13g2_a21oi_1 _17755_ (.A1(\soc_inst.cpu_core.alu.b[19] ),
    .A2(\soc_inst.cpu_core.alu.a[19] ),
    .Y(_03475_),
    .B1(_03474_));
 sg13g2_o21ai_1 _17756_ (.B1(_03475_),
    .Y(_03476_),
    .A1(_03430_),
    .A2(_03471_));
 sg13g2_nor3_1 _17757_ (.A(_02792_),
    .B(_03473_),
    .C(_03476_),
    .Y(_03477_));
 sg13g2_o21ai_1 _17758_ (.B1(_02792_),
    .Y(_03478_),
    .A1(_03473_),
    .A2(_03476_));
 sg13g2_nand2_1 _17759_ (.Y(_03479_),
    .A(net4427),
    .B(_03478_));
 sg13g2_mux2_1 _17760_ (.A0(net4860),
    .A1(net4861),
    .S(net4840),
    .X(_03480_));
 sg13g2_mux2_1 _17761_ (.A0(_03480_),
    .A1(_03437_),
    .S(net4831),
    .X(_03481_));
 sg13g2_mux2_1 _17762_ (.A0(_03398_),
    .A1(_03481_),
    .S(net4722),
    .X(_03482_));
 sg13g2_a22oi_1 _17763_ (.Y(_03483_),
    .B1(_03482_),
    .B2(net4210),
    .A2(_03312_),
    .A1(net4209));
 sg13g2_a21oi_1 _17764_ (.A1(_03119_),
    .A2(_03483_),
    .Y(_03484_),
    .B1(net4802));
 sg13g2_nor2_1 _17765_ (.A(_03129_),
    .B(_03407_),
    .Y(_03485_));
 sg13g2_o21ai_1 _17766_ (.B1(net4437),
    .Y(_03486_),
    .A1(\soc_inst.cpu_core.alu.b[20] ),
    .A2(net4860));
 sg13g2_o21ai_1 _17767_ (.B1(_03486_),
    .Y(_03487_),
    .A1(_02793_),
    .A2(_03011_));
 sg13g2_o21ai_1 _17768_ (.B1(_03379_),
    .Y(_03488_),
    .A1(_02791_),
    .A2(net4432));
 sg13g2_nor4_1 _17769_ (.A(_03484_),
    .B(_03485_),
    .C(_03487_),
    .D(_03488_),
    .Y(_03489_));
 sg13g2_o21ai_1 _17770_ (.B1(_03489_),
    .Y(_03490_),
    .A1(_03477_),
    .A2(_03479_));
 sg13g2_a21oi_2 _17771_ (.B1(_03490_),
    .Y(_03491_),
    .A2(_03470_),
    .A1(_03468_));
 sg13g2_nand2_1 _17772_ (.Y(_03492_),
    .A(net4914),
    .B(net736));
 sg13g2_o21ai_1 _17773_ (.B1(_03492_),
    .Y(_01406_),
    .A1(net4111),
    .A2(_03491_));
 sg13g2_a21o_1 _17774_ (.A2(_03468_),
    .A1(_02806_),
    .B1(_02789_),
    .X(_03493_));
 sg13g2_nand3_1 _17775_ (.B(_02806_),
    .C(_03468_),
    .A(_02789_),
    .Y(_03494_));
 sg13g2_nand3_1 _17776_ (.B(_03493_),
    .C(_03494_),
    .A(net4447),
    .Y(_03495_));
 sg13g2_nand3_1 _17777_ (.B(_02791_),
    .C(_03478_),
    .A(_02790_),
    .Y(_03496_));
 sg13g2_a21o_1 _17778_ (.A2(_03478_),
    .A1(_02791_),
    .B1(_02790_),
    .X(_03497_));
 sg13g2_nand3_1 _17779_ (.B(_03496_),
    .C(_03497_),
    .A(net4425),
    .Y(_03498_));
 sg13g2_and2_1 _17780_ (.A(net4820),
    .B(_03420_),
    .X(_03499_));
 sg13g2_o21ai_1 _17781_ (.B1(_02958_),
    .Y(_03500_),
    .A1(_05798_),
    .A2(net4839));
 sg13g2_mux2_1 _17782_ (.A0(_03500_),
    .A1(_03455_),
    .S(net4827),
    .X(_03501_));
 sg13g2_a21oi_1 _17783_ (.A1(net4722),
    .A2(_03501_),
    .Y(_03502_),
    .B1(_03499_));
 sg13g2_a21o_1 _17784_ (.A2(_03501_),
    .A1(net4722),
    .B1(_03499_),
    .X(_03503_));
 sg13g2_a221oi_1 _17785_ (.B2(net4210),
    .C1(_03146_),
    .B1(_03503_),
    .A1(net4209),
    .Y(_03504_),
    .A2(_03335_));
 sg13g2_nand2b_1 _17786_ (.Y(_03505_),
    .B(net4436),
    .A_N(_02788_));
 sg13g2_o21ai_1 _17787_ (.B1(_03505_),
    .Y(_03506_),
    .A1(_02787_),
    .A2(_02936_));
 sg13g2_a221oi_1 _17788_ (.B2(net4804),
    .C1(_03506_),
    .B1(_03212_),
    .A1(_02789_),
    .Y(_03507_),
    .A2(net4428));
 sg13g2_o21ai_1 _17789_ (.B1(_03507_),
    .Y(_03508_),
    .A1(net4804),
    .A2(_03504_));
 sg13g2_a21oi_1 _17790_ (.A1(_03158_),
    .A2(net4208),
    .Y(_03509_),
    .B1(_03508_));
 sg13g2_nand3_1 _17791_ (.B(_03498_),
    .C(_03509_),
    .A(_03495_),
    .Y(_03510_));
 sg13g2_a22oi_1 _17792_ (.Y(_03511_),
    .B1(_02673_),
    .B2(_03510_),
    .A2(net2643),
    .A1(net4898));
 sg13g2_inv_1 _17793_ (.Y(_01407_),
    .A(_03511_));
 sg13g2_nand3_1 _17794_ (.B(_02805_),
    .C(_03493_),
    .A(_02785_),
    .Y(_03512_));
 sg13g2_a21oi_1 _17795_ (.A1(_02805_),
    .A2(_03493_),
    .Y(_03513_),
    .B1(_02785_));
 sg13g2_nor2_1 _17796_ (.A(net4444),
    .B(_03513_),
    .Y(_03514_));
 sg13g2_and2_1 _17797_ (.A(_02788_),
    .B(_03497_),
    .X(_03515_));
 sg13g2_nor2_1 _17798_ (.A(_02784_),
    .B(_03515_),
    .Y(_03516_));
 sg13g2_xnor2_1 _17799_ (.Y(_03517_),
    .A(_02785_),
    .B(_03515_));
 sg13g2_o21ai_1 _17800_ (.B1(_02869_),
    .Y(_03518_),
    .A1(_05796_),
    .A2(net4839));
 sg13g2_mux2_1 _17801_ (.A0(_03518_),
    .A1(_03480_),
    .S(net4828),
    .X(_03519_));
 sg13g2_mux2_1 _17802_ (.A0(_03438_),
    .A1(_03519_),
    .S(net4721),
    .X(_03520_));
 sg13g2_a22oi_1 _17803_ (.Y(_03521_),
    .B1(_03520_),
    .B2(net4210),
    .A2(_03352_),
    .A1(net4209));
 sg13g2_a21o_1 _17804_ (.A2(_03521_),
    .A1(_03174_),
    .B1(net4802),
    .X(_03522_));
 sg13g2_nand2_1 _17805_ (.Y(_03523_),
    .A(_03188_),
    .B(net4208));
 sg13g2_o21ai_1 _17806_ (.B1(net4437),
    .Y(_03524_),
    .A1(\soc_inst.cpu_core.alu.b[22] ),
    .A2(\soc_inst.cpu_core.alu.a[22] ));
 sg13g2_o21ai_1 _17807_ (.B1(_03524_),
    .Y(_03525_),
    .A1(_02783_),
    .A2(net4432));
 sg13g2_a21oi_1 _17808_ (.A1(_02785_),
    .A2(net4428),
    .Y(_03526_),
    .B1(_03525_));
 sg13g2_nand4_1 _17809_ (.B(_03522_),
    .C(_03523_),
    .A(net4067),
    .Y(_03527_),
    .D(_03526_));
 sg13g2_a221oi_1 _17810_ (.B2(net4425),
    .C1(_03527_),
    .B1(_03517_),
    .A1(_03512_),
    .Y(_03528_),
    .A2(_03514_));
 sg13g2_nand2_1 _17811_ (.Y(_03529_),
    .A(net4900),
    .B(net2213));
 sg13g2_o21ai_1 _17812_ (.B1(_03529_),
    .Y(_01408_),
    .A1(net4111),
    .A2(_03528_));
 sg13g2_nor2_1 _17813_ (.A(_02803_),
    .B(_03513_),
    .Y(_03530_));
 sg13g2_xnor2_1 _17814_ (.Y(_03531_),
    .A(_02782_),
    .B(_03530_));
 sg13g2_mux2_1 _17815_ (.A0(net4859),
    .A1(\soc_inst.cpu_core.alu.a[22] ),
    .S(net4841),
    .X(_03532_));
 sg13g2_mux2_1 _17816_ (.A0(_03532_),
    .A1(_03500_),
    .S(net4827),
    .X(_03533_));
 sg13g2_mux2_1 _17817_ (.A0(_03456_),
    .A1(_03533_),
    .S(net4721),
    .X(_03534_));
 sg13g2_a221oi_1 _17818_ (.B2(net4210),
    .C1(_03218_),
    .B1(_03534_),
    .A1(net4209),
    .Y(_03535_),
    .A2(_03375_));
 sg13g2_a21oi_1 _17819_ (.A1(_02780_),
    .A2(net4428),
    .Y(_03536_),
    .B1(net4437));
 sg13g2_nand2b_1 _17820_ (.Y(_03537_),
    .B(net4434),
    .A_N(_02780_));
 sg13g2_o21ai_1 _17821_ (.B1(_03537_),
    .Y(_03538_),
    .A1(_02779_),
    .A2(_03536_));
 sg13g2_a221oi_1 _17822_ (.B2(_03206_),
    .C1(_03538_),
    .B1(net4208),
    .A1(net4802),
    .Y(_03539_),
    .A2(_03212_));
 sg13g2_o21ai_1 _17823_ (.B1(_03539_),
    .Y(_03540_),
    .A1(net4802),
    .A2(_03535_));
 sg13g2_a21oi_1 _17824_ (.A1(\soc_inst.cpu_core.alu.b[22] ),
    .A2(\soc_inst.cpu_core.alu.a[22] ),
    .Y(_03541_),
    .B1(_03516_));
 sg13g2_xnor2_1 _17825_ (.Y(_03542_),
    .A(_02781_),
    .B(_03541_));
 sg13g2_a221oi_1 _17826_ (.B2(net4425),
    .C1(_03540_),
    .B1(_03542_),
    .A1(net4446),
    .Y(_03543_),
    .A2(_03531_));
 sg13g2_nand2_1 _17827_ (.Y(_03544_),
    .A(net4897),
    .B(net1974));
 sg13g2_o21ai_1 _17828_ (.B1(_03544_),
    .Y(_01409_),
    .A1(net4111),
    .A2(_03543_));
 sg13g2_nor2_1 _17829_ (.A(_02782_),
    .B(_02784_),
    .Y(_03545_));
 sg13g2_nand3_1 _17830_ (.B(_02792_),
    .C(_03545_),
    .A(_02789_),
    .Y(_03546_));
 sg13g2_inv_1 _17831_ (.Y(_03547_),
    .A(_03546_));
 sg13g2_o21ai_1 _17832_ (.B1(_03547_),
    .Y(_03548_),
    .A1(_03473_),
    .A2(_03476_));
 sg13g2_o21ai_1 _17833_ (.B1(_02780_),
    .Y(_03549_),
    .A1(_02779_),
    .A2(_02783_));
 sg13g2_o21ai_1 _17834_ (.B1(_02788_),
    .Y(_03550_),
    .A1(_02787_),
    .A2(_02791_));
 sg13g2_a21oi_2 _17835_ (.B1(_03549_),
    .Y(_03551_),
    .A2(_03550_),
    .A1(_03545_));
 sg13g2_nand3_1 _17836_ (.B(_03548_),
    .C(_03551_),
    .A(_02835_),
    .Y(_03552_));
 sg13g2_a21oi_2 _17837_ (.B1(_02835_),
    .Y(_03553_),
    .A2(_03551_),
    .A1(_03548_));
 sg13g2_nor2_1 _17838_ (.A(net4424),
    .B(_03553_),
    .Y(_03554_));
 sg13g2_o21ai_1 _17839_ (.B1(_02936_),
    .Y(_03555_),
    .A1(_02832_),
    .A2(_03011_));
 sg13g2_a221oi_1 _17840_ (.B2(_02833_),
    .C1(_03378_),
    .B1(_03555_),
    .A1(_02832_),
    .Y(_03556_),
    .A2(net4435));
 sg13g2_o21ai_1 _17841_ (.B1(_03556_),
    .Y(_03557_),
    .A1(_02911_),
    .A2(_03236_));
 sg13g2_nor2_1 _17842_ (.A(net4735),
    .B(_03232_),
    .Y(_03558_));
 sg13g2_a21o_1 _17843_ (.A2(net4841),
    .A1(net4859),
    .B1(_02887_),
    .X(_03559_));
 sg13g2_mux2_1 _17844_ (.A0(_03559_),
    .A1(_03518_),
    .S(net4827),
    .X(_03560_));
 sg13g2_nand2_1 _17845_ (.Y(_03561_),
    .A(net4820),
    .B(_03481_));
 sg13g2_a21oi_1 _17846_ (.A1(net4721),
    .A2(_03560_),
    .Y(_03562_),
    .B1(net4813));
 sg13g2_a221oi_1 _17847_ (.B2(_03562_),
    .C1(_02947_),
    .B1(_03561_),
    .A1(net4813),
    .Y(_03563_),
    .A2(_03400_));
 sg13g2_nor3_1 _17848_ (.A(_03557_),
    .B(_03558_),
    .C(_03563_),
    .Y(_03564_));
 sg13g2_nand2_1 _17849_ (.Y(_03565_),
    .A(_02819_),
    .B(_02835_));
 sg13g2_xnor2_1 _17850_ (.Y(_03566_),
    .A(_02819_),
    .B(_02835_));
 sg13g2_o21ai_1 _17851_ (.B1(_03564_),
    .Y(_03567_),
    .A1(net4444),
    .A2(_03566_));
 sg13g2_a21oi_2 _17852_ (.B1(_03567_),
    .Y(_03568_),
    .A2(_03554_),
    .A1(_03552_));
 sg13g2_nand2_1 _17853_ (.Y(_03569_),
    .A(net4905),
    .B(net2619));
 sg13g2_o21ai_1 _17854_ (.B1(_03569_),
    .Y(_01410_),
    .A1(net4111),
    .A2(_03568_));
 sg13g2_or3_1 _17855_ (.A(net4442),
    .B(_02832_),
    .C(_03553_),
    .X(_03570_));
 sg13g2_o21ai_1 _17856_ (.B1(net4442),
    .Y(_03571_),
    .A1(_02832_),
    .A2(_03553_));
 sg13g2_nand3_1 _17857_ (.B(_03570_),
    .C(_03571_),
    .A(net4426),
    .Y(_03572_));
 sg13g2_nor2_1 _17858_ (.A(net4442),
    .B(_03565_),
    .Y(_03573_));
 sg13g2_nand3_1 _17859_ (.B(_02837_),
    .C(_03565_),
    .A(_02830_),
    .Y(_03574_));
 sg13g2_nor3_1 _17860_ (.A(net4445),
    .B(_02838_),
    .C(_03573_),
    .Y(_03575_));
 sg13g2_mux2_1 _17861_ (.A0(net4858),
    .A1(\soc_inst.cpu_core.alu.a[24] ),
    .S(net4841),
    .X(_03576_));
 sg13g2_mux2_1 _17862_ (.A0(_03576_),
    .A1(_03532_),
    .S(net4824),
    .X(_03577_));
 sg13g2_nor2_1 _17863_ (.A(net4817),
    .B(_03577_),
    .Y(_03578_));
 sg13g2_o21ai_1 _17864_ (.B1(net4731),
    .Y(_03579_),
    .A1(net4720),
    .A2(_03501_));
 sg13g2_nor2_1 _17865_ (.A(_03578_),
    .B(_03579_),
    .Y(_03580_));
 sg13g2_and2_1 _17866_ (.A(net4815),
    .B(_03421_),
    .X(_03581_));
 sg13g2_o21ai_1 _17867_ (.B1(net4211),
    .Y(_03582_),
    .A1(_03580_),
    .A2(_03581_));
 sg13g2_nor2_1 _17868_ (.A(_02829_),
    .B(net4433),
    .Y(_03583_));
 sg13g2_a221oi_1 _17869_ (.B2(net4442),
    .C1(_03583_),
    .B1(net4429),
    .A1(_02828_),
    .Y(_03584_),
    .A2(net4439));
 sg13g2_a22oi_1 _17870_ (.Y(_03585_),
    .B1(_03406_),
    .B2(_03255_),
    .A2(_03262_),
    .A1(net4735));
 sg13g2_nand4_1 _17871_ (.B(_03582_),
    .C(_03584_),
    .A(net4067),
    .Y(_03586_),
    .D(_03585_));
 sg13g2_a21oi_1 _17872_ (.A1(_03574_),
    .A2(_03575_),
    .Y(_03587_),
    .B1(_03586_));
 sg13g2_a21oi_2 _17873_ (.B1(net4112),
    .Y(_03588_),
    .A2(_03587_),
    .A1(_03572_));
 sg13g2_a21o_1 _17874_ (.A2(net2919),
    .A1(net4891),
    .B1(_03588_),
    .X(_01411_));
 sg13g2_nand3_1 _17875_ (.B(_02829_),
    .C(_03571_),
    .A(_02821_),
    .Y(_03589_));
 sg13g2_a21oi_1 _17876_ (.A1(_02829_),
    .A2(_03571_),
    .Y(_03590_),
    .B1(_02821_));
 sg13g2_nor2_1 _17877_ (.A(net4424),
    .B(_03590_),
    .Y(_03591_));
 sg13g2_o21ai_1 _17878_ (.B1(_02839_),
    .Y(_03592_),
    .A1(net4442),
    .A2(_03565_));
 sg13g2_xnor2_1 _17879_ (.Y(_03593_),
    .A(_02820_),
    .B(_03592_));
 sg13g2_mux2_1 _17880_ (.A0(net4856),
    .A1(net4858),
    .S(net4841),
    .X(_03594_));
 sg13g2_mux2_1 _17881_ (.A0(_03594_),
    .A1(_03559_),
    .S(net4825),
    .X(_03595_));
 sg13g2_mux2_1 _17882_ (.A0(_03519_),
    .A1(_03595_),
    .S(net4719),
    .X(_03596_));
 sg13g2_nor2_1 _17883_ (.A(net4810),
    .B(_03596_),
    .Y(_03597_));
 sg13g2_o21ai_1 _17884_ (.B1(net4212),
    .Y(_03598_),
    .A1(net4731),
    .A2(_03439_));
 sg13g2_nand2_1 _17885_ (.Y(_03599_),
    .A(_02820_),
    .B(net4429));
 sg13g2_o21ai_1 _17886_ (.B1(net4439),
    .Y(_03600_),
    .A1(\soc_inst.cpu_core.alu.b[26] ),
    .A2(net4856));
 sg13g2_nand3_1 _17887_ (.B(net4856),
    .C(net4435),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .Y(_03601_));
 sg13g2_nand4_1 _17888_ (.B(_03599_),
    .C(_03600_),
    .A(net4067),
    .Y(_03602_),
    .D(_03601_));
 sg13g2_a221oi_1 _17889_ (.B2(_03278_),
    .C1(_03602_),
    .B1(_03406_),
    .A1(net4735),
    .Y(_03603_),
    .A2(_03282_));
 sg13g2_o21ai_1 _17890_ (.B1(_03603_),
    .Y(_03604_),
    .A1(_03597_),
    .A2(_03598_));
 sg13g2_a221oi_1 _17891_ (.B2(_02670_),
    .C1(_03604_),
    .B1(_03593_),
    .A1(_03589_),
    .Y(_03605_),
    .A2(_03591_));
 sg13g2_nand2_1 _17892_ (.Y(_03606_),
    .A(net4887),
    .B(net2648));
 sg13g2_o21ai_1 _17893_ (.B1(_03606_),
    .Y(_01412_),
    .A1(net4112),
    .A2(_03605_));
 sg13g2_a21oi_1 _17894_ (.A1(\soc_inst.cpu_core.alu.b[26] ),
    .A2(net4857),
    .Y(_03607_),
    .B1(_03590_));
 sg13g2_xnor2_1 _17895_ (.Y(_03608_),
    .A(_02825_),
    .B(_03607_));
 sg13g2_a21o_1 _17896_ (.A2(_03592_),
    .A1(_02821_),
    .B1(_02840_),
    .X(_03609_));
 sg13g2_nor2_1 _17897_ (.A(_02826_),
    .B(_03609_),
    .Y(_03610_));
 sg13g2_nand2_1 _17898_ (.Y(_03611_),
    .A(_02826_),
    .B(_03609_));
 sg13g2_nor2_1 _17899_ (.A(net4445),
    .B(_03610_),
    .Y(_03612_));
 sg13g2_a21oi_1 _17900_ (.A1(net4856),
    .A2(net4843),
    .Y(_03613_),
    .B1(_02963_));
 sg13g2_nand2_1 _17901_ (.Y(_03614_),
    .A(net4825),
    .B(_03576_));
 sg13g2_o21ai_1 _17902_ (.B1(_03614_),
    .Y(_03615_),
    .A1(net4829),
    .A2(_03613_));
 sg13g2_nand2b_1 _17903_ (.Y(_03616_),
    .B(net4819),
    .A_N(_03533_));
 sg13g2_o21ai_1 _17904_ (.B1(_03616_),
    .Y(_03617_),
    .A1(net4818),
    .A2(_03615_));
 sg13g2_nand2_1 _17905_ (.Y(_03618_),
    .A(net4810),
    .B(_03457_));
 sg13g2_o21ai_1 _17906_ (.B1(_03618_),
    .Y(_03619_),
    .A1(net4810),
    .A2(_03617_));
 sg13g2_nand2b_1 _17907_ (.Y(_03620_),
    .B(net4435),
    .A_N(_02824_));
 sg13g2_a22oi_1 _17908_ (.Y(_03621_),
    .B1(net4429),
    .B2(_02825_),
    .A2(net4439),
    .A1(_02823_));
 sg13g2_nand3_1 _17909_ (.B(_03620_),
    .C(_03621_),
    .A(net4067),
    .Y(_03622_));
 sg13g2_a221oi_1 _17910_ (.B2(net4211),
    .C1(_03622_),
    .B1(_03619_),
    .A1(_03298_),
    .Y(_03623_),
    .A2(_03406_));
 sg13g2_o21ai_1 _17911_ (.B1(_03623_),
    .Y(_03624_),
    .A1(net4806),
    .A2(_03291_));
 sg13g2_a221oi_1 _17912_ (.B2(_03612_),
    .C1(_03624_),
    .B1(_03611_),
    .A1(net4426),
    .Y(_03625_),
    .A2(_03608_));
 sg13g2_nand2_1 _17913_ (.Y(_03626_),
    .A(net4919),
    .B(net2476));
 sg13g2_o21ai_1 _17914_ (.B1(_03626_),
    .Y(_01413_),
    .A1(net4112),
    .A2(_03625_));
 sg13g2_nand4_1 _17915_ (.B(_02825_),
    .C(net4442),
    .A(_02820_),
    .Y(_03627_),
    .D(_02834_));
 sg13g2_a21oi_1 _17916_ (.A1(_03548_),
    .A2(_03551_),
    .Y(_03628_),
    .B1(_03627_));
 sg13g2_nand3_1 _17917_ (.B(net4857),
    .C(_02823_),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .Y(_03629_));
 sg13g2_o21ai_1 _17918_ (.B1(_02829_),
    .Y(_03630_),
    .A1(_02827_),
    .A2(_02831_));
 sg13g2_nand3_1 _17919_ (.B(_02825_),
    .C(_03630_),
    .A(_02820_),
    .Y(_03631_));
 sg13g2_nand3_1 _17920_ (.B(_03629_),
    .C(_03631_),
    .A(_02824_),
    .Y(_03632_));
 sg13g2_nor3_1 _17921_ (.A(_02848_),
    .B(_03628_),
    .C(_03632_),
    .Y(_03633_));
 sg13g2_o21ai_1 _17922_ (.B1(_02848_),
    .Y(_03634_),
    .A1(_03628_),
    .A2(_03632_));
 sg13g2_nand2_1 _17923_ (.Y(_03635_),
    .A(net4425),
    .B(_03634_));
 sg13g2_xnor2_1 _17924_ (.Y(_03636_),
    .A(_02844_),
    .B(_02849_));
 sg13g2_or2_1 _17925_ (.X(_03637_),
    .B(_03482_),
    .A(net4730));
 sg13g2_a21o_1 _17926_ (.A2(net4842),
    .A1(\soc_inst.cpu_core.alu.a[27] ),
    .B1(_02881_),
    .X(_03638_));
 sg13g2_a22oi_1 _17927_ (.Y(_03639_),
    .B1(_03638_),
    .B2(_02924_),
    .A2(_03594_),
    .A1(_02923_));
 sg13g2_a21oi_1 _17928_ (.A1(net4819),
    .A2(_03560_),
    .Y(_03640_),
    .B1(net4810));
 sg13g2_a21oi_1 _17929_ (.A1(_03639_),
    .A2(_03640_),
    .Y(_03641_),
    .B1(_02947_));
 sg13g2_o21ai_1 _17930_ (.B1(net4437),
    .Y(_03642_),
    .A1(\soc_inst.cpu_core.alu.b[28] ),
    .A2(\soc_inst.cpu_core.alu.a[28] ));
 sg13g2_nand2_1 _17931_ (.Y(_03643_),
    .A(_02848_),
    .B(net4428));
 sg13g2_nand2b_1 _17932_ (.Y(_03644_),
    .B(net4434),
    .A_N(_02847_));
 sg13g2_nand4_1 _17933_ (.B(_03642_),
    .C(_03643_),
    .A(net4067),
    .Y(_03645_),
    .D(_03644_));
 sg13g2_a21oi_1 _17934_ (.A1(_03637_),
    .A2(_03641_),
    .Y(_03646_),
    .B1(_03645_));
 sg13g2_o21ai_1 _17935_ (.B1(_03646_),
    .Y(_03647_),
    .A1(net4802),
    .A2(_03318_));
 sg13g2_a221oi_1 _17936_ (.B2(net4446),
    .C1(_03647_),
    .B1(_03636_),
    .A1(_03314_),
    .Y(_03648_),
    .A2(net4208));
 sg13g2_o21ai_1 _17937_ (.B1(_03648_),
    .Y(_03649_),
    .A1(_03633_),
    .A2(_03635_));
 sg13g2_a22oi_1 _17938_ (.Y(_03650_),
    .B1(_02673_),
    .B2(_03649_),
    .A2(net2793),
    .A1(net4901));
 sg13g2_inv_1 _17939_ (.Y(_01414_),
    .A(_03650_));
 sg13g2_nand3_1 _17940_ (.B(_02847_),
    .C(_03634_),
    .A(_02846_),
    .Y(_03651_));
 sg13g2_nor2_1 _17941_ (.A(_02846_),
    .B(_02849_),
    .Y(_03652_));
 sg13g2_o21ai_1 _17942_ (.B1(_03652_),
    .Y(_03653_),
    .A1(_03628_),
    .A2(_03632_));
 sg13g2_or2_1 _17943_ (.X(_03654_),
    .B(_02847_),
    .A(_02846_));
 sg13g2_nand4_1 _17944_ (.B(_03651_),
    .C(_03653_),
    .A(net4425),
    .Y(_03655_),
    .D(_03654_));
 sg13g2_nor2_1 _17945_ (.A(_02846_),
    .B(_02852_),
    .Y(_03656_));
 sg13g2_o21ai_1 _17946_ (.B1(_03656_),
    .Y(_03657_),
    .A1(_02844_),
    .A2(_02848_));
 sg13g2_nor3_1 _17947_ (.A(net4445),
    .B(_02851_),
    .C(_02853_),
    .Y(_03658_));
 sg13g2_and2_1 _17948_ (.A(_03657_),
    .B(_03658_),
    .X(_03659_));
 sg13g2_nor2_1 _17949_ (.A(net4720),
    .B(_03577_),
    .Y(_03660_));
 sg13g2_nor2_1 _17950_ (.A(_02964_),
    .B(_02968_),
    .Y(_03661_));
 sg13g2_a221oi_1 _17951_ (.B2(_02924_),
    .C1(_03660_),
    .B1(_03661_),
    .A1(_02923_),
    .Y(_03662_),
    .A2(_03613_));
 sg13g2_a21oi_1 _17952_ (.A1(net4810),
    .A2(_03502_),
    .Y(_03663_),
    .B1(_02947_));
 sg13g2_o21ai_1 _17953_ (.B1(_03663_),
    .Y(_03664_),
    .A1(net4810),
    .A2(_03662_));
 sg13g2_nor2_1 _17954_ (.A(_03337_),
    .B(_03407_),
    .Y(_03665_));
 sg13g2_o21ai_1 _17955_ (.B1(net4437),
    .Y(_03666_),
    .A1(\soc_inst.cpu_core.alu.b[29] ),
    .A2(\soc_inst.cpu_core.alu.a[29] ));
 sg13g2_o21ai_1 _17956_ (.B1(_03666_),
    .Y(_03667_),
    .A1(_02846_),
    .A2(_03011_));
 sg13g2_o21ai_1 _17957_ (.B1(net4067),
    .Y(_03668_),
    .A1(_02845_),
    .A2(net4433));
 sg13g2_nor2_1 _17958_ (.A(net4803),
    .B(_03339_),
    .Y(_03669_));
 sg13g2_nor4_1 _17959_ (.A(_03665_),
    .B(_03667_),
    .C(_03668_),
    .D(_03669_),
    .Y(_03670_));
 sg13g2_nand3_1 _17960_ (.B(_03664_),
    .C(_03670_),
    .A(_03655_),
    .Y(_03671_));
 sg13g2_o21ai_1 _17961_ (.B1(_02673_),
    .Y(_03672_),
    .A1(_03659_),
    .A2(_03671_));
 sg13g2_o21ai_1 _17962_ (.B1(_03672_),
    .Y(_01415_),
    .A1(net4751),
    .A2(_05779_));
 sg13g2_and2_1 _17963_ (.A(_02845_),
    .B(_03654_),
    .X(_03673_));
 sg13g2_a21oi_1 _17964_ (.A1(_03653_),
    .A2(_03673_),
    .Y(_03674_),
    .B1(_02857_));
 sg13g2_nand3_1 _17965_ (.B(_03653_),
    .C(_03673_),
    .A(_02857_),
    .Y(_03675_));
 sg13g2_nor2_1 _17966_ (.A(net4424),
    .B(_03674_),
    .Y(_03676_));
 sg13g2_o21ai_1 _17967_ (.B1(net4446),
    .Y(_03677_),
    .A1(_02855_),
    .A2(_02857_));
 sg13g2_or2_1 _17968_ (.X(_03678_),
    .B(_03520_),
    .A(net4730));
 sg13g2_a21oi_1 _17969_ (.A1(\soc_inst.cpu_core.alu.a[29] ),
    .A2(net4843),
    .Y(_03679_),
    .B1(_02883_));
 sg13g2_nor2_1 _17970_ (.A(net4659),
    .B(_03679_),
    .Y(_03680_));
 sg13g2_a221oi_1 _17971_ (.B2(_02923_),
    .C1(_03680_),
    .B1(_03638_),
    .A1(net4817),
    .Y(_03681_),
    .A2(_03595_));
 sg13g2_a21oi_1 _17972_ (.A1(net4730),
    .A2(_03681_),
    .Y(_03682_),
    .B1(_02947_));
 sg13g2_nand2_1 _17973_ (.Y(_03683_),
    .A(net4735),
    .B(_03356_));
 sg13g2_o21ai_1 _17974_ (.B1(_02936_),
    .Y(_03684_),
    .A1(_02856_),
    .A2(_03011_));
 sg13g2_o21ai_1 _17975_ (.B1(_03684_),
    .Y(_03685_),
    .A1(\soc_inst.cpu_core.alu.b[30] ),
    .A2(\soc_inst.cpu_core.alu.a[30] ));
 sg13g2_a21oi_1 _17976_ (.A1(_02856_),
    .A2(net4434),
    .Y(_03686_),
    .B1(_03378_));
 sg13g2_nand3_1 _17977_ (.B(_03685_),
    .C(_03686_),
    .A(_03683_),
    .Y(_03687_));
 sg13g2_a221oi_1 _17978_ (.B2(_03682_),
    .C1(_03687_),
    .B1(_03678_),
    .A1(_03354_),
    .Y(_03688_),
    .A2(net4208));
 sg13g2_o21ai_1 _17979_ (.B1(_03688_),
    .Y(_03689_),
    .A1(_02858_),
    .A2(_03677_));
 sg13g2_a21o_1 _17980_ (.A2(_03676_),
    .A1(_03675_),
    .B1(_03689_),
    .X(_03690_));
 sg13g2_and2_1 _17981_ (.A(net4901),
    .B(net2940),
    .X(_03691_));
 sg13g2_a21o_1 _17982_ (.A2(_03690_),
    .A1(_02673_),
    .B1(_03691_),
    .X(_01416_));
 sg13g2_nor2_1 _17983_ (.A(_02856_),
    .B(_03674_),
    .Y(_03692_));
 sg13g2_xnor2_1 _17984_ (.Y(_03693_),
    .A(_02676_),
    .B(_03692_));
 sg13g2_xor2_1 _17985_ (.B(_02860_),
    .A(_02676_),
    .X(_03694_));
 sg13g2_nand2_1 _17986_ (.Y(_03695_),
    .A(net4817),
    .B(_03615_));
 sg13g2_o21ai_1 _17987_ (.B1(_02923_),
    .Y(_03696_),
    .A1(_02964_),
    .A2(_02968_));
 sg13g2_nand3_1 _17988_ (.B(net4843),
    .C(_02924_),
    .A(\soc_inst.cpu_core.alu.a[30] ),
    .Y(_03697_));
 sg13g2_nand4_1 _17989_ (.B(_03695_),
    .C(_03696_),
    .A(_03215_),
    .Y(_03698_),
    .D(_03697_));
 sg13g2_a221oi_1 _17990_ (.B2(net4210),
    .C1(_03382_),
    .B1(_03698_),
    .A1(net4209),
    .Y(_03699_),
    .A2(_03534_));
 sg13g2_a21oi_1 _17991_ (.A1(_02676_),
    .A2(net4431),
    .Y(_03700_),
    .B1(_03212_));
 sg13g2_nand3_1 _17992_ (.B(net4854),
    .C(net4434),
    .A(\soc_inst.cpu_core.alu.b[31] ),
    .Y(_03701_));
 sg13g2_o21ai_1 _17993_ (.B1(net4437),
    .Y(_03702_),
    .A1(\soc_inst.cpu_core.alu.b[31] ),
    .A2(net4854));
 sg13g2_nand3_1 _17994_ (.B(_03701_),
    .C(_03702_),
    .A(_03700_),
    .Y(_03703_));
 sg13g2_a21oi_1 _17995_ (.A1(_03376_),
    .A2(net4208),
    .Y(_03704_),
    .B1(_03703_));
 sg13g2_o21ai_1 _17996_ (.B1(_03704_),
    .Y(_03705_),
    .A1(net4805),
    .A2(_03699_));
 sg13g2_a221oi_1 _17997_ (.B2(net4446),
    .C1(_03705_),
    .B1(_03694_),
    .A1(net4425),
    .Y(_03706_),
    .A2(_03693_));
 sg13g2_nand2_1 _17998_ (.Y(_03707_),
    .A(net4885),
    .B(net2291));
 sg13g2_o21ai_1 _17999_ (.B1(_03707_),
    .Y(_01417_),
    .A1(net4112),
    .A2(_03706_));
 sg13g2_nand2_1 _18000_ (.Y(_03708_),
    .A(net4971),
    .B(net350));
 sg13g2_o21ai_1 _18001_ (.B1(_03708_),
    .Y(_01418_),
    .A1(_09212_),
    .A2(_09217_));
 sg13g2_a21oi_1 _18002_ (.A1(net4973),
    .A2(_05720_),
    .Y(_01419_),
    .B1(net542));
 sg13g2_nand3b_1 _18003_ (.B(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .C(\soc_inst.cpu_core.mem_reg_we ),
    .Y(_03709_),
    .A_N(\soc_inst.cpu_core._unused_mem_rd_addr[0] ));
 sg13g2_nor2_1 _18004_ (.A(_07213_),
    .B(_03709_),
    .Y(_03710_));
 sg13g2_nor2_1 _18005_ (.A(net1164),
    .B(net4418),
    .Y(_03711_));
 sg13g2_a21oi_1 _18006_ (.A1(net3945),
    .A2(net4418),
    .Y(_01420_),
    .B1(_03711_));
 sg13g2_nor2_1 _18007_ (.A(net1080),
    .B(net4417),
    .Y(_03712_));
 sg13g2_a21oi_1 _18008_ (.A1(net3943),
    .A2(net4417),
    .Y(_01421_),
    .B1(_03712_));
 sg13g2_nor2_1 _18009_ (.A(net1289),
    .B(net4422),
    .Y(_03713_));
 sg13g2_a21oi_1 _18010_ (.A1(net3940),
    .A2(net4422),
    .Y(_01422_),
    .B1(_03713_));
 sg13g2_nor2_1 _18011_ (.A(net1442),
    .B(net4417),
    .Y(_03714_));
 sg13g2_a21oi_1 _18012_ (.A1(net3938),
    .A2(net4417),
    .Y(_01423_),
    .B1(_03714_));
 sg13g2_nor2_1 _18013_ (.A(net1489),
    .B(net4419),
    .Y(_03715_));
 sg13g2_a21oi_1 _18014_ (.A1(net3835),
    .A2(net4419),
    .Y(_01424_),
    .B1(_03715_));
 sg13g2_nor2_1 _18015_ (.A(net1292),
    .B(net4419),
    .Y(_03716_));
 sg13g2_a21oi_1 _18016_ (.A1(net3935),
    .A2(net4419),
    .Y(_01425_),
    .B1(_03716_));
 sg13g2_nor2_1 _18017_ (.A(net1652),
    .B(net4419),
    .Y(_03717_));
 sg13g2_a21oi_1 _18018_ (.A1(net3932),
    .A2(net4419),
    .Y(_01426_),
    .B1(_03717_));
 sg13g2_nor2_1 _18019_ (.A(net1498),
    .B(net4417),
    .Y(_03718_));
 sg13g2_a21oi_1 _18020_ (.A1(net3930),
    .A2(net4417),
    .Y(_01427_),
    .B1(_03718_));
 sg13g2_nor2_1 _18021_ (.A(net1624),
    .B(net4414),
    .Y(_03719_));
 sg13g2_a21oi_1 _18022_ (.A1(net3929),
    .A2(net4414),
    .Y(_01428_),
    .B1(_03719_));
 sg13g2_nor2_1 _18023_ (.A(net767),
    .B(net4421),
    .Y(_03720_));
 sg13g2_a21oi_1 _18024_ (.A1(net3927),
    .A2(net4421),
    .Y(_01429_),
    .B1(_03720_));
 sg13g2_nor2_1 _18025_ (.A(net1068),
    .B(net4418),
    .Y(_03721_));
 sg13g2_a21oi_1 _18026_ (.A1(net3925),
    .A2(net4418),
    .Y(_01430_),
    .B1(_03721_));
 sg13g2_nor2_1 _18027_ (.A(net1375),
    .B(net4417),
    .Y(_03722_));
 sg13g2_a21oi_1 _18028_ (.A1(net3922),
    .A2(net4417),
    .Y(_01431_),
    .B1(_03722_));
 sg13g2_nor2_1 _18029_ (.A(net685),
    .B(net4420),
    .Y(_03723_));
 sg13g2_a21oi_1 _18030_ (.A1(net3833),
    .A2(net4420),
    .Y(_01432_),
    .B1(_03723_));
 sg13g2_nor2_1 _18031_ (.A(net1342),
    .B(net4414),
    .Y(_03724_));
 sg13g2_a21oi_1 _18032_ (.A1(net3919),
    .A2(net4414),
    .Y(_01433_),
    .B1(_03724_));
 sg13g2_nor2_1 _18033_ (.A(net1045),
    .B(net4420),
    .Y(_03725_));
 sg13g2_a21oi_1 _18034_ (.A1(net3917),
    .A2(net4420),
    .Y(_01434_),
    .B1(_03725_));
 sg13g2_nor2_1 _18035_ (.A(net1577),
    .B(net4416),
    .Y(_03726_));
 sg13g2_a21oi_1 _18036_ (.A1(net3916),
    .A2(net4416),
    .Y(_01435_),
    .B1(_03726_));
 sg13g2_nor2_1 _18037_ (.A(net729),
    .B(net4414),
    .Y(_03727_));
 sg13g2_a21oi_1 _18038_ (.A1(net3911),
    .A2(net4414),
    .Y(_01436_),
    .B1(_03727_));
 sg13g2_nor2_1 _18039_ (.A(net1796),
    .B(net4415),
    .Y(_03728_));
 sg13g2_a21oi_1 _18040_ (.A1(net3831),
    .A2(net4415),
    .Y(_01437_),
    .B1(_03728_));
 sg13g2_nor2_1 _18041_ (.A(net1793),
    .B(net4413),
    .Y(_03729_));
 sg13g2_a21oi_1 _18042_ (.A1(net3910),
    .A2(net4413),
    .Y(_01438_),
    .B1(_03729_));
 sg13g2_nor2_1 _18043_ (.A(net1403),
    .B(net4415),
    .Y(_03730_));
 sg13g2_a21oi_1 _18044_ (.A1(net3906),
    .A2(net4415),
    .Y(_01439_),
    .B1(_03730_));
 sg13g2_nor2_1 _18045_ (.A(net976),
    .B(net4413),
    .Y(_03731_));
 sg13g2_a21oi_1 _18046_ (.A1(net3905),
    .A2(net4413),
    .Y(_01440_),
    .B1(_03731_));
 sg13g2_nor2_1 _18047_ (.A(net813),
    .B(net4416),
    .Y(_03732_));
 sg13g2_a21oi_1 _18048_ (.A1(net3902),
    .A2(net4416),
    .Y(_01441_),
    .B1(_03732_));
 sg13g2_nor2_1 _18049_ (.A(net1340),
    .B(net4415),
    .Y(_03733_));
 sg13g2_a21oi_1 _18050_ (.A1(net3900),
    .A2(net4415),
    .Y(_01442_),
    .B1(_03733_));
 sg13g2_nor2_1 _18051_ (.A(net1194),
    .B(net4413),
    .Y(_03734_));
 sg13g2_a21oi_1 _18052_ (.A1(net3899),
    .A2(net4413),
    .Y(_01443_),
    .B1(_03734_));
 sg13g2_nor2_1 _18053_ (.A(net963),
    .B(net4421),
    .Y(_03735_));
 sg13g2_a21oi_1 _18054_ (.A1(net3830),
    .A2(net4421),
    .Y(_01444_),
    .B1(_03735_));
 sg13g2_nor2_1 _18055_ (.A(net1732),
    .B(net4421),
    .Y(_03736_));
 sg13g2_a21oi_1 _18056_ (.A1(net3828),
    .A2(net4421),
    .Y(_01445_),
    .B1(_03736_));
 sg13g2_nor2_1 _18057_ (.A(net1586),
    .B(net4418),
    .Y(_03737_));
 sg13g2_a21oi_1 _18058_ (.A1(net3825),
    .A2(net4418),
    .Y(_01446_),
    .B1(_03737_));
 sg13g2_nor2_1 _18059_ (.A(net1410),
    .B(net4416),
    .Y(_03738_));
 sg13g2_a21oi_1 _18060_ (.A1(net3896),
    .A2(net4416),
    .Y(_01447_),
    .B1(_03738_));
 sg13g2_nor2_1 _18061_ (.A(net1535),
    .B(net4413),
    .Y(_03739_));
 sg13g2_a21oi_1 _18062_ (.A1(net3823),
    .A2(net4413),
    .Y(_01448_),
    .B1(_03739_));
 sg13g2_nor2_1 _18063_ (.A(net1873),
    .B(net4415),
    .Y(_03740_));
 sg13g2_a21oi_1 _18064_ (.A1(net3819),
    .A2(net4415),
    .Y(_01449_),
    .B1(_03740_));
 sg13g2_nor2_1 _18065_ (.A(net798),
    .B(net4419),
    .Y(_03741_));
 sg13g2_a21oi_1 _18066_ (.A1(net3893),
    .A2(net4419),
    .Y(_01450_),
    .B1(_03741_));
 sg13g2_nor2_1 _18067_ (.A(net1617),
    .B(net4418),
    .Y(_03742_));
 sg13g2_a21oi_1 _18068_ (.A1(net3817),
    .A2(net4418),
    .Y(_01451_),
    .B1(_03742_));
 sg13g2_nand3b_1 _18069_ (.B(\soc_inst.cpu_core.mem_reg_we ),
    .C(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .Y(_03743_),
    .A_N(\soc_inst.cpu_core._unused_mem_rd_addr[1] ));
 sg13g2_nor2_2 _18070_ (.A(_07213_),
    .B(_03743_),
    .Y(_03744_));
 sg13g2_nor2_1 _18071_ (.A(net1101),
    .B(net4409),
    .Y(_03745_));
 sg13g2_a21oi_1 _18072_ (.A1(net3944),
    .A2(net4409),
    .Y(_01452_),
    .B1(_03745_));
 sg13g2_nor2_1 _18073_ (.A(net782),
    .B(net4409),
    .Y(_03746_));
 sg13g2_a21oi_1 _18074_ (.A1(net3943),
    .A2(net4408),
    .Y(_01453_),
    .B1(_03746_));
 sg13g2_nor2_1 _18075_ (.A(net772),
    .B(net4408),
    .Y(_03747_));
 sg13g2_a21oi_1 _18076_ (.A1(net3940),
    .A2(net4408),
    .Y(_01454_),
    .B1(_03747_));
 sg13g2_nor2_1 _18077_ (.A(net1269),
    .B(net4408),
    .Y(_03748_));
 sg13g2_a21oi_1 _18078_ (.A1(net3938),
    .A2(net4408),
    .Y(_01455_),
    .B1(_03748_));
 sg13g2_nor2_1 _18079_ (.A(net2044),
    .B(net4410),
    .Y(_03749_));
 sg13g2_a21oi_1 _18080_ (.A1(net3835),
    .A2(net4410),
    .Y(_01456_),
    .B1(_03749_));
 sg13g2_nor2_1 _18081_ (.A(net1368),
    .B(net4410),
    .Y(_03750_));
 sg13g2_a21oi_1 _18082_ (.A1(net3935),
    .A2(net4410),
    .Y(_01457_),
    .B1(_03750_));
 sg13g2_nor2_1 _18083_ (.A(net791),
    .B(net4410),
    .Y(_03751_));
 sg13g2_a21oi_1 _18084_ (.A1(net3934),
    .A2(net4410),
    .Y(_01458_),
    .B1(_03751_));
 sg13g2_nor2_1 _18085_ (.A(net1447),
    .B(net4412),
    .Y(_03752_));
 sg13g2_a21oi_1 _18086_ (.A1(net3931),
    .A2(net4408),
    .Y(_01459_),
    .B1(_03752_));
 sg13g2_nor2_1 _18087_ (.A(net1891),
    .B(net4404),
    .Y(_03753_));
 sg13g2_a21oi_1 _18088_ (.A1(net3928),
    .A2(net4404),
    .Y(_01460_),
    .B1(_03753_));
 sg13g2_nor2_1 _18089_ (.A(net1231),
    .B(net4411),
    .Y(_03754_));
 sg13g2_a21oi_1 _18090_ (.A1(net3926),
    .A2(net4411),
    .Y(_01461_),
    .B1(_03754_));
 sg13g2_nor2_1 _18091_ (.A(net1610),
    .B(net4409),
    .Y(_03755_));
 sg13g2_a21oi_1 _18092_ (.A1(net3924),
    .A2(net4409),
    .Y(_01462_),
    .B1(_03755_));
 sg13g2_nor2_1 _18093_ (.A(net1011),
    .B(net4408),
    .Y(_03756_));
 sg13g2_a21oi_1 _18094_ (.A1(net3923),
    .A2(net4408),
    .Y(_01463_),
    .B1(_03756_));
 sg13g2_nor2_1 _18095_ (.A(net984),
    .B(net4412),
    .Y(_03757_));
 sg13g2_a21oi_1 _18096_ (.A1(net3833),
    .A2(net4411),
    .Y(_01464_),
    .B1(_03757_));
 sg13g2_nor2_1 _18097_ (.A(net1082),
    .B(net4404),
    .Y(_03758_));
 sg13g2_a21oi_1 _18098_ (.A1(net3920),
    .A2(net4404),
    .Y(_01465_),
    .B1(_03758_));
 sg13g2_nor2_1 _18099_ (.A(net1224),
    .B(net4410),
    .Y(_03759_));
 sg13g2_a21oi_1 _18100_ (.A1(net3917),
    .A2(net4410),
    .Y(_01466_),
    .B1(_03759_));
 sg13g2_nor2_1 _18101_ (.A(net1275),
    .B(net4406),
    .Y(_03760_));
 sg13g2_a21oi_1 _18102_ (.A1(net3914),
    .A2(net4406),
    .Y(_01467_),
    .B1(_03760_));
 sg13g2_nor2_1 _18103_ (.A(net1223),
    .B(net4404),
    .Y(_03761_));
 sg13g2_a21oi_1 _18104_ (.A1(net3911),
    .A2(net4404),
    .Y(_01468_),
    .B1(_03761_));
 sg13g2_nor2_1 _18105_ (.A(net1237),
    .B(net4405),
    .Y(_03762_));
 sg13g2_a21oi_1 _18106_ (.A1(net3831),
    .A2(net4405),
    .Y(_01469_),
    .B1(_03762_));
 sg13g2_nor2_1 _18107_ (.A(net893),
    .B(net4403),
    .Y(_03763_));
 sg13g2_a21oi_1 _18108_ (.A1(net3909),
    .A2(net4403),
    .Y(_01470_),
    .B1(_03763_));
 sg13g2_nor2_1 _18109_ (.A(net1413),
    .B(net4405),
    .Y(_03764_));
 sg13g2_a21oi_1 _18110_ (.A1(net3906),
    .A2(net4405),
    .Y(_01471_),
    .B1(_03764_));
 sg13g2_nor2_1 _18111_ (.A(net924),
    .B(net4403),
    .Y(_03765_));
 sg13g2_a21oi_1 _18112_ (.A1(net3904),
    .A2(net4403),
    .Y(_01472_),
    .B1(_03765_));
 sg13g2_nor2_1 _18113_ (.A(net982),
    .B(net4405),
    .Y(_03766_));
 sg13g2_a21oi_1 _18114_ (.A1(net3902),
    .A2(net4405),
    .Y(_01473_),
    .B1(_03766_));
 sg13g2_nor2_1 _18115_ (.A(net969),
    .B(net4405),
    .Y(_03767_));
 sg13g2_a21oi_1 _18116_ (.A1(net3901),
    .A2(net4405),
    .Y(_01474_),
    .B1(_03767_));
 sg13g2_nor2_1 _18117_ (.A(net1704),
    .B(net4403),
    .Y(_03768_));
 sg13g2_a21oi_1 _18118_ (.A1(net3897),
    .A2(net4403),
    .Y(_01475_),
    .B1(_03768_));
 sg13g2_nor2_1 _18119_ (.A(net1284),
    .B(net4406),
    .Y(_03769_));
 sg13g2_a21oi_1 _18120_ (.A1(net3830),
    .A2(net4406),
    .Y(_01476_),
    .B1(_03769_));
 sg13g2_nor2_1 _18121_ (.A(net1595),
    .B(net4411),
    .Y(_03770_));
 sg13g2_a21oi_1 _18122_ (.A1(net3827),
    .A2(net4411),
    .Y(_01477_),
    .B1(_03770_));
 sg13g2_nor2_1 _18123_ (.A(net1697),
    .B(net4409),
    .Y(_03771_));
 sg13g2_a21oi_1 _18124_ (.A1(net3824),
    .A2(net4409),
    .Y(_01478_),
    .B1(_03771_));
 sg13g2_nor2_1 _18125_ (.A(net992),
    .B(net4406),
    .Y(_03772_));
 sg13g2_a21oi_1 _18126_ (.A1(net3895),
    .A2(net4407),
    .Y(_01479_),
    .B1(_03772_));
 sg13g2_nor2_1 _18127_ (.A(net1566),
    .B(net4403),
    .Y(_03773_));
 sg13g2_a21oi_1 _18128_ (.A1(net3821),
    .A2(net4403),
    .Y(_01480_),
    .B1(_03773_));
 sg13g2_nor2_1 _18129_ (.A(net846),
    .B(net4406),
    .Y(_03774_));
 sg13g2_a21oi_1 _18130_ (.A1(net3819),
    .A2(net4406),
    .Y(_01481_),
    .B1(_03774_));
 sg13g2_nor2_1 _18131_ (.A(net1640),
    .B(net4411),
    .Y(_03775_));
 sg13g2_a21oi_1 _18132_ (.A1(net3893),
    .A2(net4411),
    .Y(_01482_),
    .B1(_03775_));
 sg13g2_nor2_1 _18133_ (.A(net1616),
    .B(net4404),
    .Y(_03776_));
 sg13g2_a21oi_1 _18134_ (.A1(net3817),
    .A2(net4404),
    .Y(_01483_),
    .B1(_03776_));
 sg13g2_nor4_2 _18135_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .C(_05481_),
    .Y(_03777_),
    .D(_07213_));
 sg13g2_nor2_1 _18136_ (.A(net687),
    .B(net4399),
    .Y(_03778_));
 sg13g2_a21oi_1 _18137_ (.A1(net3945),
    .A2(net4399),
    .Y(_01484_),
    .B1(_03778_));
 sg13g2_nor2_1 _18138_ (.A(net1110),
    .B(net4398),
    .Y(_03779_));
 sg13g2_a21oi_1 _18139_ (.A1(net3942),
    .A2(net4398),
    .Y(_01485_),
    .B1(_03779_));
 sg13g2_nor2_1 _18140_ (.A(net1098),
    .B(net4398),
    .Y(_03780_));
 sg13g2_a21oi_1 _18141_ (.A1(net3940),
    .A2(net4399),
    .Y(_01486_),
    .B1(_03780_));
 sg13g2_nor2_1 _18142_ (.A(net1219),
    .B(net4398),
    .Y(_03781_));
 sg13g2_a21oi_1 _18143_ (.A1(net3938),
    .A2(net4398),
    .Y(_01487_),
    .B1(_03781_));
 sg13g2_nor2_1 _18144_ (.A(net1680),
    .B(net4401),
    .Y(_03782_));
 sg13g2_a21oi_1 _18145_ (.A1(net3836),
    .A2(net4401),
    .Y(_01488_),
    .B1(_03782_));
 sg13g2_nor2_1 _18146_ (.A(net1349),
    .B(net4401),
    .Y(_03783_));
 sg13g2_a21oi_1 _18147_ (.A1(net3935),
    .A2(net4401),
    .Y(_01489_),
    .B1(_03783_));
 sg13g2_nor2_1 _18148_ (.A(net995),
    .B(net4401),
    .Y(_03784_));
 sg13g2_a21oi_1 _18149_ (.A1(net3932),
    .A2(net4401),
    .Y(_01490_),
    .B1(_03784_));
 sg13g2_nor2_1 _18150_ (.A(net1352),
    .B(net4402),
    .Y(_03785_));
 sg13g2_a21oi_1 _18151_ (.A1(net3931),
    .A2(net4398),
    .Y(_01491_),
    .B1(_03785_));
 sg13g2_nor2_1 _18152_ (.A(net904),
    .B(net4394),
    .Y(_03786_));
 sg13g2_a21oi_1 _18153_ (.A1(net3928),
    .A2(net4394),
    .Y(_01492_),
    .B1(_03786_));
 sg13g2_nor2_1 _18154_ (.A(net1230),
    .B(net4400),
    .Y(_03787_));
 sg13g2_a21oi_1 _18155_ (.A1(net3926),
    .A2(net4400),
    .Y(_01493_),
    .B1(_03787_));
 sg13g2_nor2_1 _18156_ (.A(net1178),
    .B(net4399),
    .Y(_03788_));
 sg13g2_a21oi_1 _18157_ (.A1(net3924),
    .A2(net4399),
    .Y(_01494_),
    .B1(_03788_));
 sg13g2_nor2_1 _18158_ (.A(net1100),
    .B(net4398),
    .Y(_03789_));
 sg13g2_a21oi_1 _18159_ (.A1(net3922),
    .A2(net4398),
    .Y(_01495_),
    .B1(_03789_));
 sg13g2_nor2_1 _18160_ (.A(net1551),
    .B(net4400),
    .Y(_03790_));
 sg13g2_a21oi_1 _18161_ (.A1(net3833),
    .A2(net4400),
    .Y(_01496_),
    .B1(_03790_));
 sg13g2_nor2_1 _18162_ (.A(net1316),
    .B(net4394),
    .Y(_03791_));
 sg13g2_a21oi_1 _18163_ (.A1(net3921),
    .A2(net4394),
    .Y(_01497_),
    .B1(_03791_));
 sg13g2_nor2_1 _18164_ (.A(net1337),
    .B(net4400),
    .Y(_03792_));
 sg13g2_a21oi_1 _18165_ (.A1(net3917),
    .A2(net4400),
    .Y(_01498_),
    .B1(_03792_));
 sg13g2_nor2_1 _18166_ (.A(net1864),
    .B(net4396),
    .Y(_03793_));
 sg13g2_a21oi_1 _18167_ (.A1(net3914),
    .A2(net4396),
    .Y(_01499_),
    .B1(_03793_));
 sg13g2_nor2_1 _18168_ (.A(net1583),
    .B(net4393),
    .Y(_03794_));
 sg13g2_a21oi_1 _18169_ (.A1(net3911),
    .A2(net4393),
    .Y(_01500_),
    .B1(_03794_));
 sg13g2_nor2_1 _18170_ (.A(net1338),
    .B(net4395),
    .Y(_03795_));
 sg13g2_a21oi_1 _18171_ (.A1(net3831),
    .A2(net4396),
    .Y(_01501_),
    .B1(_03795_));
 sg13g2_nor2_1 _18172_ (.A(net1233),
    .B(net4393),
    .Y(_03796_));
 sg13g2_a21oi_1 _18173_ (.A1(net3909),
    .A2(net4393),
    .Y(_01502_),
    .B1(_03796_));
 sg13g2_nor2_1 _18174_ (.A(net894),
    .B(net4395),
    .Y(_03797_));
 sg13g2_a21oi_1 _18175_ (.A1(net3908),
    .A2(net4395),
    .Y(_01503_),
    .B1(_03797_));
 sg13g2_nor2_1 _18176_ (.A(net1788),
    .B(net4393),
    .Y(_03798_));
 sg13g2_a21oi_1 _18177_ (.A1(net3904),
    .A2(net4393),
    .Y(_01504_),
    .B1(_03798_));
 sg13g2_nor2_1 _18178_ (.A(net1142),
    .B(net4395),
    .Y(_03799_));
 sg13g2_a21oi_1 _18179_ (.A1(net3902),
    .A2(net4396),
    .Y(_01505_),
    .B1(_03799_));
 sg13g2_nor2_1 _18180_ (.A(net891),
    .B(net4395),
    .Y(_03800_));
 sg13g2_a21oi_1 _18181_ (.A1(net3901),
    .A2(net4395),
    .Y(_01506_),
    .B1(_03800_));
 sg13g2_nor2_1 _18182_ (.A(net1402),
    .B(net4393),
    .Y(_03801_));
 sg13g2_a21oi_1 _18183_ (.A1(net3897),
    .A2(net4393),
    .Y(_01507_),
    .B1(_03801_));
 sg13g2_nor2_1 _18184_ (.A(net1165),
    .B(net4396),
    .Y(_03802_));
 sg13g2_a21oi_1 _18185_ (.A1(net3829),
    .A2(net4396),
    .Y(_01508_),
    .B1(_03802_));
 sg13g2_nor2_1 _18186_ (.A(net1735),
    .B(net4400),
    .Y(_03803_));
 sg13g2_a21oi_1 _18187_ (.A1(net3826),
    .A2(net4400),
    .Y(_01509_),
    .B1(_03803_));
 sg13g2_nor2_1 _18188_ (.A(net1058),
    .B(net4399),
    .Y(_03804_));
 sg13g2_a21oi_1 _18189_ (.A1(net3824),
    .A2(net4399),
    .Y(_01510_),
    .B1(_03804_));
 sg13g2_nor2_1 _18190_ (.A(net1370),
    .B(net4396),
    .Y(_03805_));
 sg13g2_a21oi_1 _18191_ (.A1(net3895),
    .A2(net4397),
    .Y(_01511_),
    .B1(_03805_));
 sg13g2_nor2_1 _18192_ (.A(net792),
    .B(net4394),
    .Y(_03806_));
 sg13g2_a21oi_1 _18193_ (.A1(net3822),
    .A2(net4394),
    .Y(_01512_),
    .B1(_03806_));
 sg13g2_nor2_1 _18194_ (.A(net1139),
    .B(net4395),
    .Y(_03807_));
 sg13g2_a21oi_1 _18195_ (.A1(net3819),
    .A2(net4395),
    .Y(_01513_),
    .B1(_03807_));
 sg13g2_nor2_1 _18196_ (.A(net920),
    .B(net4401),
    .Y(_03808_));
 sg13g2_a21oi_1 _18197_ (.A1(net3893),
    .A2(net4401),
    .Y(_01514_),
    .B1(_03808_));
 sg13g2_nor2_1 _18198_ (.A(net2440),
    .B(net4397),
    .Y(_03809_));
 sg13g2_a21oi_1 _18199_ (.A1(net3818),
    .A2(net4394),
    .Y(_01515_),
    .B1(_03809_));
 sg13g2_nand2b_2 _18200_ (.Y(_03810_),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .A_N(\soc_inst.cpu_core._unused_mem_rd_addr[2] ));
 sg13g2_nor2_1 _18201_ (.A(_07212_),
    .B(_03810_),
    .Y(_03811_));
 sg13g2_nor2_1 _18202_ (.A(net1759),
    .B(net4388),
    .Y(_03812_));
 sg13g2_a21oi_1 _18203_ (.A1(net3944),
    .A2(net4388),
    .Y(_01516_),
    .B1(_03812_));
 sg13g2_nor2_1 _18204_ (.A(net1181),
    .B(net4387),
    .Y(_03813_));
 sg13g2_a21oi_1 _18205_ (.A1(net3942),
    .A2(net4388),
    .Y(_01517_),
    .B1(_03813_));
 sg13g2_nor2_1 _18206_ (.A(net839),
    .B(net4387),
    .Y(_03814_));
 sg13g2_a21oi_1 _18207_ (.A1(net3941),
    .A2(net4391),
    .Y(_01518_),
    .B1(_03814_));
 sg13g2_nor2_1 _18208_ (.A(net1367),
    .B(net4387),
    .Y(_03815_));
 sg13g2_a21oi_1 _18209_ (.A1(net3939),
    .A2(net4387),
    .Y(_01519_),
    .B1(_03815_));
 sg13g2_nor2_1 _18210_ (.A(net892),
    .B(net4390),
    .Y(_03816_));
 sg13g2_a21oi_1 _18211_ (.A1(net3836),
    .A2(net4391),
    .Y(_01520_),
    .B1(_03816_));
 sg13g2_nor2_1 _18212_ (.A(net1703),
    .B(net4390),
    .Y(_03817_));
 sg13g2_a21oi_1 _18213_ (.A1(net3936),
    .A2(net4390),
    .Y(_01521_),
    .B1(_03817_));
 sg13g2_nor2_1 _18214_ (.A(net1755),
    .B(net4390),
    .Y(_03818_));
 sg13g2_a21oi_1 _18215_ (.A1(net3932),
    .A2(net4390),
    .Y(_01522_),
    .B1(_03818_));
 sg13g2_nor2_1 _18216_ (.A(net1348),
    .B(net4387),
    .Y(_03819_));
 sg13g2_a21oi_1 _18217_ (.A1(net3931),
    .A2(net4387),
    .Y(_01523_),
    .B1(_03819_));
 sg13g2_nor2_1 _18218_ (.A(net1910),
    .B(net4384),
    .Y(_03820_));
 sg13g2_a21oi_1 _18219_ (.A1(net3928),
    .A2(net4384),
    .Y(_01524_),
    .B1(_03820_));
 sg13g2_nor2_1 _18220_ (.A(net1227),
    .B(net4389),
    .Y(_03821_));
 sg13g2_a21oi_1 _18221_ (.A1(net3926),
    .A2(net4389),
    .Y(_01525_),
    .B1(_03821_));
 sg13g2_nor2_1 _18222_ (.A(net1655),
    .B(net4388),
    .Y(_03822_));
 sg13g2_a21oi_1 _18223_ (.A1(net3925),
    .A2(net4388),
    .Y(_01526_),
    .B1(_03822_));
 sg13g2_nor2_1 _18224_ (.A(net1111),
    .B(net4387),
    .Y(_03823_));
 sg13g2_a21oi_1 _18225_ (.A1(net3922),
    .A2(net4387),
    .Y(_01527_),
    .B1(_03823_));
 sg13g2_nor2_1 _18226_ (.A(net1240),
    .B(net4391),
    .Y(_03824_));
 sg13g2_a21oi_1 _18227_ (.A1(net3833),
    .A2(net4391),
    .Y(_01528_),
    .B1(_03824_));
 sg13g2_nor2_1 _18228_ (.A(net744),
    .B(net4384),
    .Y(_03825_));
 sg13g2_a21oi_1 _18229_ (.A1(net3919),
    .A2(net4384),
    .Y(_01529_),
    .B1(_03825_));
 sg13g2_nor2_1 _18230_ (.A(net1108),
    .B(net4390),
    .Y(_03826_));
 sg13g2_a21oi_1 _18231_ (.A1(net3918),
    .A2(net4390),
    .Y(_01530_),
    .B1(_03826_));
 sg13g2_nor2_1 _18232_ (.A(net900),
    .B(net4386),
    .Y(_03827_));
 sg13g2_a21oi_1 _18233_ (.A1(net3914),
    .A2(net4386),
    .Y(_01531_),
    .B1(_03827_));
 sg13g2_nor2_1 _18234_ (.A(net1326),
    .B(net4384),
    .Y(_03828_));
 sg13g2_a21oi_1 _18235_ (.A1(net3911),
    .A2(net4384),
    .Y(_01532_),
    .B1(_03828_));
 sg13g2_nor2_1 _18236_ (.A(net1303),
    .B(net4385),
    .Y(_03829_));
 sg13g2_a21oi_1 _18237_ (.A1(net3832),
    .A2(net4385),
    .Y(_01533_),
    .B1(_03829_));
 sg13g2_nor2_1 _18238_ (.A(net1290),
    .B(net4383),
    .Y(_03830_));
 sg13g2_a21oi_1 _18239_ (.A1(net3909),
    .A2(net4383),
    .Y(_01534_),
    .B1(_03830_));
 sg13g2_nor2_1 _18240_ (.A(net1781),
    .B(net4385),
    .Y(_03831_));
 sg13g2_a21oi_1 _18241_ (.A1(net3906),
    .A2(net4385),
    .Y(_01535_),
    .B1(_03831_));
 sg13g2_nor2_1 _18242_ (.A(net1835),
    .B(net4383),
    .Y(_03832_));
 sg13g2_a21oi_1 _18243_ (.A1(net3904),
    .A2(net4383),
    .Y(_01536_),
    .B1(_03832_));
 sg13g2_nor2_1 _18244_ (.A(net771),
    .B(net4386),
    .Y(_03833_));
 sg13g2_a21oi_1 _18245_ (.A1(net3902),
    .A2(net4386),
    .Y(_01537_),
    .B1(_03833_));
 sg13g2_nor2_1 _18246_ (.A(net1134),
    .B(net4385),
    .Y(_03834_));
 sg13g2_a21oi_1 _18247_ (.A1(net3901),
    .A2(net4385),
    .Y(_01538_),
    .B1(_03834_));
 sg13g2_nor2_1 _18248_ (.A(net1210),
    .B(net4383),
    .Y(_03835_));
 sg13g2_a21oi_1 _18249_ (.A1(net3897),
    .A2(net4383),
    .Y(_01539_),
    .B1(_03835_));
 sg13g2_nor2_1 _18250_ (.A(net1542),
    .B(net4389),
    .Y(_03836_));
 sg13g2_a21oi_1 _18251_ (.A1(net3829),
    .A2(net4389),
    .Y(_01540_),
    .B1(_03836_));
 sg13g2_nor2_1 _18252_ (.A(net702),
    .B(net4389),
    .Y(_03837_));
 sg13g2_a21oi_1 _18253_ (.A1(net3826),
    .A2(net4389),
    .Y(_01541_),
    .B1(_03837_));
 sg13g2_nor2_1 _18254_ (.A(net624),
    .B(net4388),
    .Y(_03838_));
 sg13g2_a21oi_1 _18255_ (.A1(net3824),
    .A2(net4388),
    .Y(_01542_),
    .B1(_03838_));
 sg13g2_nor2_1 _18256_ (.A(net728),
    .B(net4386),
    .Y(_03839_));
 sg13g2_a21oi_1 _18257_ (.A1(net3895),
    .A2(net4386),
    .Y(_01543_),
    .B1(_03839_));
 sg13g2_nor2_1 _18258_ (.A(net1401),
    .B(net4383),
    .Y(_03840_));
 sg13g2_a21oi_1 _18259_ (.A1(net3822),
    .A2(net4383),
    .Y(_01544_),
    .B1(_03840_));
 sg13g2_nor2_1 _18260_ (.A(net1009),
    .B(net4385),
    .Y(_03841_));
 sg13g2_a21oi_1 _18261_ (.A1(net3819),
    .A2(net4385),
    .Y(_01545_),
    .B1(_03841_));
 sg13g2_nor2_1 _18262_ (.A(net1216),
    .B(net4389),
    .Y(_03842_));
 sg13g2_a21oi_1 _18263_ (.A1(net3894),
    .A2(net4389),
    .Y(_01546_),
    .B1(_03842_));
 sg13g2_nor2_1 _18264_ (.A(net1205),
    .B(net4384),
    .Y(_03843_));
 sg13g2_a21oi_1 _18265_ (.A1(net3817),
    .A2(net4384),
    .Y(_01547_),
    .B1(_03843_));
 sg13g2_nor2_2 _18266_ (.A(_03709_),
    .B(_03810_),
    .Y(_03844_));
 sg13g2_nor2_1 _18267_ (.A(net1060),
    .B(net4378),
    .Y(_03845_));
 sg13g2_a21oi_1 _18268_ (.A1(net3944),
    .A2(net4378),
    .Y(_01548_),
    .B1(_03845_));
 sg13g2_nor2_1 _18269_ (.A(net1843),
    .B(net4379),
    .Y(_03846_));
 sg13g2_a21oi_1 _18270_ (.A1(net3942),
    .A2(net4379),
    .Y(_01549_),
    .B1(_03846_));
 sg13g2_nor2_1 _18271_ (.A(net1127),
    .B(net4378),
    .Y(_03847_));
 sg13g2_a21oi_1 _18272_ (.A1(net3940),
    .A2(net4378),
    .Y(_01550_),
    .B1(_03847_));
 sg13g2_nor2_1 _18273_ (.A(net1783),
    .B(net4379),
    .Y(_03848_));
 sg13g2_a21oi_1 _18274_ (.A1(net3939),
    .A2(net4379),
    .Y(_01551_),
    .B1(_03848_));
 sg13g2_nor2_1 _18275_ (.A(net1081),
    .B(net4381),
    .Y(_03849_));
 sg13g2_a21oi_1 _18276_ (.A1(net3836),
    .A2(net4381),
    .Y(_01552_),
    .B1(_03849_));
 sg13g2_nor2_1 _18277_ (.A(net2217),
    .B(net4381),
    .Y(_03850_));
 sg13g2_a21oi_1 _18278_ (.A1(net3936),
    .A2(net4381),
    .Y(_01553_),
    .B1(_03850_));
 sg13g2_nor2_1 _18279_ (.A(net1580),
    .B(net4381),
    .Y(_03851_));
 sg13g2_a21oi_1 _18280_ (.A1(net3932),
    .A2(net4381),
    .Y(_01554_),
    .B1(_03851_));
 sg13g2_nor2_1 _18281_ (.A(net1357),
    .B(net4379),
    .Y(_03852_));
 sg13g2_a21oi_1 _18282_ (.A1(net3931),
    .A2(net4379),
    .Y(_01555_),
    .B1(_03852_));
 sg13g2_nor2_1 _18283_ (.A(net1053),
    .B(net4374),
    .Y(_03853_));
 sg13g2_a21oi_1 _18284_ (.A1(net3928),
    .A2(net4374),
    .Y(_01556_),
    .B1(_03853_));
 sg13g2_nor2_1 _18285_ (.A(net1428),
    .B(net4375),
    .Y(_03854_));
 sg13g2_a21oi_1 _18286_ (.A1(net3926),
    .A2(net4375),
    .Y(_01557_),
    .B1(_03854_));
 sg13g2_nor2_1 _18287_ (.A(net1014),
    .B(net4378),
    .Y(_03855_));
 sg13g2_a21oi_1 _18288_ (.A1(net3924),
    .A2(net4378),
    .Y(_01558_),
    .B1(_03855_));
 sg13g2_nor2_1 _18289_ (.A(net1291),
    .B(net4379),
    .Y(_03856_));
 sg13g2_a21oi_1 _18290_ (.A1(net3923),
    .A2(net4379),
    .Y(_01559_),
    .B1(_03856_));
 sg13g2_nor2_1 _18291_ (.A(net980),
    .B(net4380),
    .Y(_03857_));
 sg13g2_a21oi_1 _18292_ (.A1(net3833),
    .A2(net4380),
    .Y(_01560_),
    .B1(_03857_));
 sg13g2_nor2_1 _18293_ (.A(net727),
    .B(net4374),
    .Y(_03858_));
 sg13g2_a21oi_1 _18294_ (.A1(net3920),
    .A2(net4374),
    .Y(_01561_),
    .B1(_03858_));
 sg13g2_nor2_1 _18295_ (.A(net786),
    .B(net4380),
    .Y(_03859_));
 sg13g2_a21oi_1 _18296_ (.A1(net3917),
    .A2(net4380),
    .Y(_01562_),
    .B1(_03859_));
 sg13g2_nor2_1 _18297_ (.A(net1176),
    .B(net4375),
    .Y(_03860_));
 sg13g2_a21oi_1 _18298_ (.A1(net3914),
    .A2(net4375),
    .Y(_01563_),
    .B1(_03860_));
 sg13g2_nor2_1 _18299_ (.A(net1140),
    .B(net4374),
    .Y(_03861_));
 sg13g2_a21oi_1 _18300_ (.A1(net3912),
    .A2(net4374),
    .Y(_01564_),
    .B1(_03861_));
 sg13g2_nor2_1 _18301_ (.A(net1626),
    .B(net4376),
    .Y(_03862_));
 sg13g2_a21oi_1 _18302_ (.A1(net3832),
    .A2(net4376),
    .Y(_01565_),
    .B1(_03862_));
 sg13g2_nor2_1 _18303_ (.A(net1149),
    .B(net4373),
    .Y(_03863_));
 sg13g2_a21oi_1 _18304_ (.A1(net3909),
    .A2(net4373),
    .Y(_01566_),
    .B1(_03863_));
 sg13g2_nor2_1 _18305_ (.A(net1356),
    .B(net4376),
    .Y(_03864_));
 sg13g2_a21oi_1 _18306_ (.A1(net3907),
    .A2(net4376),
    .Y(_01567_),
    .B1(_03864_));
 sg13g2_nor2_1 _18307_ (.A(net773),
    .B(net4373),
    .Y(_03865_));
 sg13g2_a21oi_1 _18308_ (.A1(net3904),
    .A2(net4373),
    .Y(_01568_),
    .B1(_03865_));
 sg13g2_nor2_1 _18309_ (.A(net1548),
    .B(net4376),
    .Y(_03866_));
 sg13g2_a21oi_1 _18310_ (.A1(net3903),
    .A2(net4376),
    .Y(_01569_),
    .B1(_03866_));
 sg13g2_nor2_1 _18311_ (.A(net814),
    .B(net4376),
    .Y(_03867_));
 sg13g2_a21oi_1 _18312_ (.A1(net3901),
    .A2(net4376),
    .Y(_01570_),
    .B1(_03867_));
 sg13g2_nor2_1 _18313_ (.A(net886),
    .B(net4373),
    .Y(_03868_));
 sg13g2_a21oi_1 _18314_ (.A1(net3897),
    .A2(net4373),
    .Y(_01571_),
    .B1(_03868_));
 sg13g2_nor2_1 _18315_ (.A(net1502),
    .B(net4375),
    .Y(_03869_));
 sg13g2_a21oi_1 _18316_ (.A1(net3829),
    .A2(net4375),
    .Y(_01572_),
    .B1(_03869_));
 sg13g2_nor2_1 _18317_ (.A(net1274),
    .B(net4380),
    .Y(_03870_));
 sg13g2_a21oi_1 _18318_ (.A1(net3826),
    .A2(net4380),
    .Y(_01573_),
    .B1(_03870_));
 sg13g2_nor2_1 _18319_ (.A(net972),
    .B(net4378),
    .Y(_03871_));
 sg13g2_a21oi_1 _18320_ (.A1(net3824),
    .A2(net4378),
    .Y(_01574_),
    .B1(_03871_));
 sg13g2_nor2_1 _18321_ (.A(net805),
    .B(net4377),
    .Y(_03872_));
 sg13g2_a21oi_1 _18322_ (.A1(net3896),
    .A2(net4375),
    .Y(_01575_),
    .B1(_03872_));
 sg13g2_nor2_1 _18323_ (.A(net1372),
    .B(net4373),
    .Y(_03873_));
 sg13g2_a21oi_1 _18324_ (.A1(net3821),
    .A2(net4373),
    .Y(_01576_),
    .B1(_03873_));
 sg13g2_nor2_1 _18325_ (.A(net803),
    .B(net4377),
    .Y(_03874_));
 sg13g2_a21oi_1 _18326_ (.A1(net3820),
    .A2(net4375),
    .Y(_01577_),
    .B1(_03874_));
 sg13g2_nor2_1 _18327_ (.A(net1163),
    .B(net4380),
    .Y(_03875_));
 sg13g2_a21oi_1 _18328_ (.A1(net3893),
    .A2(net4380),
    .Y(_01578_),
    .B1(_03875_));
 sg13g2_nor2_1 _18329_ (.A(net1281),
    .B(net4374),
    .Y(_03876_));
 sg13g2_a21oi_1 _18330_ (.A1(net3818),
    .A2(net4374),
    .Y(_01579_),
    .B1(_03876_));
 sg13g2_nor2_1 _18331_ (.A(_03743_),
    .B(_03810_),
    .Y(_03877_));
 sg13g2_nor2_1 _18332_ (.A(net758),
    .B(net4369),
    .Y(_03878_));
 sg13g2_a21oi_1 _18333_ (.A1(net3945),
    .A2(net4369),
    .Y(_01580_),
    .B1(_03878_));
 sg13g2_nor2_1 _18334_ (.A(net1637),
    .B(net4367),
    .Y(_03879_));
 sg13g2_a21oi_1 _18335_ (.A1(net3942),
    .A2(net4368),
    .Y(_01581_),
    .B1(_03879_));
 sg13g2_nor2_1 _18336_ (.A(net1043),
    .B(net4368),
    .Y(_03880_));
 sg13g2_a21oi_1 _18337_ (.A1(net3941),
    .A2(net4368),
    .Y(_01582_),
    .B1(_03880_));
 sg13g2_nor2_1 _18338_ (.A(net799),
    .B(net4367),
    .Y(_03881_));
 sg13g2_a21oi_1 _18339_ (.A1(net3938),
    .A2(net4367),
    .Y(_01583_),
    .B1(_03881_));
 sg13g2_nor2_1 _18340_ (.A(net785),
    .B(net4371),
    .Y(_03882_));
 sg13g2_a21oi_1 _18341_ (.A1(net3835),
    .A2(net4371),
    .Y(_01584_),
    .B1(_03882_));
 sg13g2_nor2_1 _18342_ (.A(net800),
    .B(net4367),
    .Y(_03883_));
 sg13g2_a21oi_1 _18343_ (.A1(net3935),
    .A2(net4368),
    .Y(_01585_),
    .B1(_03883_));
 sg13g2_nor2_1 _18344_ (.A(net1238),
    .B(net4371),
    .Y(_03884_));
 sg13g2_a21oi_1 _18345_ (.A1(net3932),
    .A2(net4371),
    .Y(_01586_),
    .B1(_03884_));
 sg13g2_nor2_1 _18346_ (.A(net1119),
    .B(net4367),
    .Y(_03885_));
 sg13g2_a21oi_1 _18347_ (.A1(net3930),
    .A2(net4367),
    .Y(_01587_),
    .B1(_03885_));
 sg13g2_nor2_1 _18348_ (.A(net868),
    .B(net4363),
    .Y(_03886_));
 sg13g2_a21oi_1 _18349_ (.A1(net3929),
    .A2(net4363),
    .Y(_01588_),
    .B1(_03886_));
 sg13g2_nor2_1 _18350_ (.A(net1360),
    .B(net4370),
    .Y(_03887_));
 sg13g2_a21oi_1 _18351_ (.A1(net3927),
    .A2(net4370),
    .Y(_01589_),
    .B1(_03887_));
 sg13g2_nor2_1 _18352_ (.A(net977),
    .B(net4369),
    .Y(_03888_));
 sg13g2_a21oi_1 _18353_ (.A1(net3925),
    .A2(net4369),
    .Y(_01590_),
    .B1(_03888_));
 sg13g2_nor2_1 _18354_ (.A(net1310),
    .B(net4367),
    .Y(_03889_));
 sg13g2_a21oi_1 _18355_ (.A1(net3923),
    .A2(net4367),
    .Y(_01591_),
    .B1(_03889_));
 sg13g2_nor2_1 _18356_ (.A(net958),
    .B(net4371),
    .Y(_03890_));
 sg13g2_a21oi_1 _18357_ (.A1(net3834),
    .A2(net4371),
    .Y(_01592_),
    .B1(_03890_));
 sg13g2_nor2_1 _18358_ (.A(net1191),
    .B(net4363),
    .Y(_03891_));
 sg13g2_a21oi_1 _18359_ (.A1(net3920),
    .A2(net4363),
    .Y(_01593_),
    .B1(_03891_));
 sg13g2_nor2_1 _18360_ (.A(net1539),
    .B(net4370),
    .Y(_03892_));
 sg13g2_a21oi_1 _18361_ (.A1(net3918),
    .A2(net4370),
    .Y(_01594_),
    .B1(_03892_));
 sg13g2_nor2_1 _18362_ (.A(net1212),
    .B(net4365),
    .Y(_03893_));
 sg13g2_a21oi_1 _18363_ (.A1(net3914),
    .A2(net4365),
    .Y(_01595_),
    .B1(_03893_));
 sg13g2_nor2_1 _18364_ (.A(net1056),
    .B(net4362),
    .Y(_03894_));
 sg13g2_a21oi_1 _18365_ (.A1(net3913),
    .A2(net4362),
    .Y(_01596_),
    .B1(_03894_));
 sg13g2_nor2_1 _18366_ (.A(net1117),
    .B(net4364),
    .Y(_03895_));
 sg13g2_a21oi_1 _18367_ (.A1(net3832),
    .A2(net4365),
    .Y(_01597_),
    .B1(_03895_));
 sg13g2_nor2_1 _18368_ (.A(net1453),
    .B(net4362),
    .Y(_03896_));
 sg13g2_a21oi_1 _18369_ (.A1(net3910),
    .A2(net4362),
    .Y(_01598_),
    .B1(_03896_));
 sg13g2_nor2_1 _18370_ (.A(net973),
    .B(net4364),
    .Y(_03897_));
 sg13g2_a21oi_1 _18371_ (.A1(net3907),
    .A2(net4364),
    .Y(_01599_),
    .B1(_03897_));
 sg13g2_nor2_1 _18372_ (.A(net1418),
    .B(net4362),
    .Y(_03898_));
 sg13g2_a21oi_1 _18373_ (.A1(net3905),
    .A2(net4362),
    .Y(_01600_),
    .B1(_03898_));
 sg13g2_nor2_1 _18374_ (.A(net913),
    .B(net4364),
    .Y(_03899_));
 sg13g2_a21oi_1 _18375_ (.A1(net3903),
    .A2(net4365),
    .Y(_01601_),
    .B1(_03899_));
 sg13g2_nor2_1 _18376_ (.A(net828),
    .B(net4364),
    .Y(_03900_));
 sg13g2_a21oi_1 _18377_ (.A1(net3900),
    .A2(net4364),
    .Y(_01602_),
    .B1(_03900_));
 sg13g2_nor2_1 _18378_ (.A(net1478),
    .B(net4362),
    .Y(_03901_));
 sg13g2_a21oi_1 _18379_ (.A1(net3897),
    .A2(net4362),
    .Y(_01603_),
    .B1(_03901_));
 sg13g2_nor2_1 _18380_ (.A(net1190),
    .B(net4365),
    .Y(_03902_));
 sg13g2_a21oi_1 _18381_ (.A1(net3829),
    .A2(net4365),
    .Y(_01604_),
    .B1(_03902_));
 sg13g2_nor2_1 _18382_ (.A(net1998),
    .B(net4370),
    .Y(_03903_));
 sg13g2_a21oi_1 _18383_ (.A1(net3826),
    .A2(net4370),
    .Y(_01605_),
    .B1(_03903_));
 sg13g2_nor2_1 _18384_ (.A(net834),
    .B(net4369),
    .Y(_03904_));
 sg13g2_a21oi_1 _18385_ (.A1(net3824),
    .A2(net4369),
    .Y(_01606_),
    .B1(_03904_));
 sg13g2_nor2_1 _18386_ (.A(net722),
    .B(net4365),
    .Y(_03905_));
 sg13g2_a21oi_1 _18387_ (.A1(net3896),
    .A2(net4366),
    .Y(_01607_),
    .B1(_03905_));
 sg13g2_nor2_1 _18388_ (.A(net964),
    .B(net4363),
    .Y(_03906_));
 sg13g2_a21oi_1 _18389_ (.A1(net3821),
    .A2(net4363),
    .Y(_01608_),
    .B1(_03906_));
 sg13g2_nor2_1 _18390_ (.A(net880),
    .B(net4364),
    .Y(_03907_));
 sg13g2_a21oi_1 _18391_ (.A1(net3819),
    .A2(net4364),
    .Y(_01609_),
    .B1(_03907_));
 sg13g2_nor2_1 _18392_ (.A(net1700),
    .B(net4370),
    .Y(_03908_));
 sg13g2_a21oi_1 _18393_ (.A1(net3893),
    .A2(net4370),
    .Y(_01610_),
    .B1(_03908_));
 sg13g2_nor2_1 _18394_ (.A(net1601),
    .B(net4363),
    .Y(_03909_));
 sg13g2_a21oi_1 _18395_ (.A1(net3818),
    .A2(net4366),
    .Y(_01611_),
    .B1(_03909_));
 sg13g2_nor4_2 _18396_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .C(_05481_),
    .Y(_03910_),
    .D(_03810_));
 sg13g2_nor2_1 _18397_ (.A(net1151),
    .B(net4357),
    .Y(_03911_));
 sg13g2_a21oi_1 _18398_ (.A1(net3944),
    .A2(net4357),
    .Y(_01612_),
    .B1(_03911_));
 sg13g2_nor2_1 _18399_ (.A(net2069),
    .B(net4358),
    .Y(_03912_));
 sg13g2_a21oi_1 _18400_ (.A1(net3943),
    .A2(net4358),
    .Y(_01613_),
    .B1(_03912_));
 sg13g2_nor2_1 _18401_ (.A(net766),
    .B(net4357),
    .Y(_03913_));
 sg13g2_a21oi_1 _18402_ (.A1(net3941),
    .A2(net4357),
    .Y(_01614_),
    .B1(_03913_));
 sg13g2_nor2_1 _18403_ (.A(net1997),
    .B(net4358),
    .Y(_03914_));
 sg13g2_a21oi_1 _18404_ (.A1(net3939),
    .A2(net4358),
    .Y(_01615_),
    .B1(_03914_));
 sg13g2_nor2_1 _18405_ (.A(net929),
    .B(net4360),
    .Y(_03915_));
 sg13g2_a21oi_1 _18406_ (.A1(net3836),
    .A2(net4360),
    .Y(_01616_),
    .B1(_03915_));
 sg13g2_nor2_1 _18407_ (.A(net1615),
    .B(net4360),
    .Y(_03916_));
 sg13g2_a21oi_1 _18408_ (.A1(net3936),
    .A2(net4360),
    .Y(_01617_),
    .B1(_03916_));
 sg13g2_nor2_1 _18409_ (.A(net1473),
    .B(net4360),
    .Y(_03917_));
 sg13g2_a21oi_1 _18410_ (.A1(net3933),
    .A2(net4360),
    .Y(_01618_),
    .B1(_03917_));
 sg13g2_nor2_1 _18411_ (.A(net1155),
    .B(net4358),
    .Y(_03918_));
 sg13g2_a21oi_1 _18412_ (.A1(net3930),
    .A2(net4358),
    .Y(_01619_),
    .B1(_03918_));
 sg13g2_nor2_1 _18413_ (.A(net1837),
    .B(net4353),
    .Y(_03919_));
 sg13g2_a21oi_1 _18414_ (.A1(net3929),
    .A2(net4353),
    .Y(_01620_),
    .B1(_03919_));
 sg13g2_nor2_1 _18415_ (.A(net1638),
    .B(net4359),
    .Y(_03920_));
 sg13g2_a21oi_1 _18416_ (.A1(net3926),
    .A2(net4359),
    .Y(_01621_),
    .B1(_03920_));
 sg13g2_nor2_1 _18417_ (.A(net1625),
    .B(net4357),
    .Y(_03921_));
 sg13g2_a21oi_1 _18418_ (.A1(net3925),
    .A2(net4357),
    .Y(_01622_),
    .B1(_03921_));
 sg13g2_nor2_1 _18419_ (.A(net851),
    .B(net4358),
    .Y(_03922_));
 sg13g2_a21oi_1 _18420_ (.A1(net3923),
    .A2(net4358),
    .Y(_01623_),
    .B1(_03922_));
 sg13g2_nor2_1 _18421_ (.A(net895),
    .B(net4360),
    .Y(_03923_));
 sg13g2_a21oi_1 _18422_ (.A1(net3834),
    .A2(net4360),
    .Y(_01624_),
    .B1(_03923_));
 sg13g2_nor2_1 _18423_ (.A(net1585),
    .B(net4353),
    .Y(_03924_));
 sg13g2_a21oi_1 _18424_ (.A1(net3919),
    .A2(net4353),
    .Y(_01625_),
    .B1(_03924_));
 sg13g2_nor2_1 _18425_ (.A(net1226),
    .B(net4359),
    .Y(_03925_));
 sg13g2_a21oi_1 _18426_ (.A1(net3917),
    .A2(net4359),
    .Y(_01626_),
    .B1(_03925_));
 sg13g2_nor2_1 _18427_ (.A(net816),
    .B(net4355),
    .Y(_03926_));
 sg13g2_a21oi_1 _18428_ (.A1(net3914),
    .A2(net4355),
    .Y(_01627_),
    .B1(_03926_));
 sg13g2_nor2_1 _18429_ (.A(net1346),
    .B(net4353),
    .Y(_03927_));
 sg13g2_a21oi_1 _18430_ (.A1(net3912),
    .A2(net4353),
    .Y(_01628_),
    .B1(_03927_));
 sg13g2_nor2_1 _18431_ (.A(net1325),
    .B(net4354),
    .Y(_03928_));
 sg13g2_a21oi_1 _18432_ (.A1(net3832),
    .A2(net4354),
    .Y(_01629_),
    .B1(_03928_));
 sg13g2_nor2_1 _18433_ (.A(net830),
    .B(net4352),
    .Y(_03929_));
 sg13g2_a21oi_1 _18434_ (.A1(net3909),
    .A2(net4352),
    .Y(_01630_),
    .B1(_03929_));
 sg13g2_nor2_1 _18435_ (.A(net996),
    .B(net4354),
    .Y(_03930_));
 sg13g2_a21oi_1 _18436_ (.A1(net3906),
    .A2(net4354),
    .Y(_01631_),
    .B1(_03930_));
 sg13g2_nor2_1 _18437_ (.A(net747),
    .B(net4352),
    .Y(_03931_));
 sg13g2_a21oi_1 _18438_ (.A1(net3905),
    .A2(net4352),
    .Y(_01632_),
    .B1(_03931_));
 sg13g2_nor2_1 _18439_ (.A(net1691),
    .B(net4355),
    .Y(_03932_));
 sg13g2_a21oi_1 _18440_ (.A1(net3902),
    .A2(net4355),
    .Y(_01633_),
    .B1(_03932_));
 sg13g2_nor2_1 _18441_ (.A(net1508),
    .B(net4354),
    .Y(_03933_));
 sg13g2_a21oi_1 _18442_ (.A1(net3901),
    .A2(net4354),
    .Y(_01634_),
    .B1(_03933_));
 sg13g2_nor2_1 _18443_ (.A(net985),
    .B(net4352),
    .Y(_03934_));
 sg13g2_a21oi_1 _18444_ (.A1(net3898),
    .A2(net4352),
    .Y(_01635_),
    .B1(_03934_));
 sg13g2_nor2_1 _18445_ (.A(net1630),
    .B(net4355),
    .Y(_03935_));
 sg13g2_a21oi_1 _18446_ (.A1(net3829),
    .A2(net4355),
    .Y(_01636_),
    .B1(_03935_));
 sg13g2_nor2_1 _18447_ (.A(net1029),
    .B(net4359),
    .Y(_03936_));
 sg13g2_a21oi_1 _18448_ (.A1(net3827),
    .A2(net4359),
    .Y(_01637_),
    .B1(_03936_));
 sg13g2_nor2_1 _18449_ (.A(net1129),
    .B(net4357),
    .Y(_03937_));
 sg13g2_a21oi_1 _18450_ (.A1(net3824),
    .A2(net4357),
    .Y(_01638_),
    .B1(_03937_));
 sg13g2_nor2_1 _18451_ (.A(net1124),
    .B(net4355),
    .Y(_03938_));
 sg13g2_a21oi_1 _18452_ (.A1(net3896),
    .A2(net4356),
    .Y(_01639_),
    .B1(_03938_));
 sg13g2_nor2_1 _18453_ (.A(net677),
    .B(net4352),
    .Y(_03939_));
 sg13g2_a21oi_1 _18454_ (.A1(net3822),
    .A2(net4352),
    .Y(_01640_),
    .B1(_03939_));
 sg13g2_nor2_1 _18455_ (.A(net1768),
    .B(net4354),
    .Y(_03940_));
 sg13g2_a21oi_1 _18456_ (.A1(net3819),
    .A2(net4354),
    .Y(_01641_),
    .B1(_03940_));
 sg13g2_nor2_1 _18457_ (.A(net757),
    .B(net4359),
    .Y(_03941_));
 sg13g2_a21oi_1 _18458_ (.A1(net3894),
    .A2(net4359),
    .Y(_01642_),
    .B1(_03941_));
 sg13g2_nor2_1 _18459_ (.A(net1328),
    .B(net4353),
    .Y(_03942_));
 sg13g2_a21oi_1 _18460_ (.A1(net3817),
    .A2(net4353),
    .Y(_01643_),
    .B1(_03942_));
 sg13g2_nand2b_2 _18461_ (.Y(_03943_),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .A_N(\soc_inst.cpu_core._unused_mem_rd_addr[3] ));
 sg13g2_nor2_2 _18462_ (.A(_07212_),
    .B(_03943_),
    .Y(_03944_));
 sg13g2_nor2_1 _18463_ (.A(net1089),
    .B(net4348),
    .Y(_03945_));
 sg13g2_a21oi_1 _18464_ (.A1(net3944),
    .A2(net4348),
    .Y(_01644_),
    .B1(_03945_));
 sg13g2_nor2_1 _18465_ (.A(net1550),
    .B(net4347),
    .Y(_03946_));
 sg13g2_a21oi_1 _18466_ (.A1(net3942),
    .A2(net4347),
    .Y(_01645_),
    .B1(_03946_));
 sg13g2_nor2_1 _18467_ (.A(net1565),
    .B(net4348),
    .Y(_03947_));
 sg13g2_a21oi_1 _18468_ (.A1(net3940),
    .A2(net4348),
    .Y(_01646_),
    .B1(_03947_));
 sg13g2_nor2_1 _18469_ (.A(net2004),
    .B(net4347),
    .Y(_03948_));
 sg13g2_a21oi_1 _18470_ (.A1(net3938),
    .A2(net4347),
    .Y(_01647_),
    .B1(_03948_));
 sg13g2_nor2_1 _18471_ (.A(net2123),
    .B(net4349),
    .Y(_03949_));
 sg13g2_a21oi_1 _18472_ (.A1(net3835),
    .A2(net4349),
    .Y(_01648_),
    .B1(_03949_));
 sg13g2_nor2_1 _18473_ (.A(net1287),
    .B(net4349),
    .Y(_03950_));
 sg13g2_a21oi_1 _18474_ (.A1(net3935),
    .A2(net4351),
    .Y(_01649_),
    .B1(_03950_));
 sg13g2_nor2_1 _18475_ (.A(net1273),
    .B(net4349),
    .Y(_03951_));
 sg13g2_a21oi_1 _18476_ (.A1(net3933),
    .A2(net4349),
    .Y(_01650_),
    .B1(_03951_));
 sg13g2_nor2_1 _18477_ (.A(net1537),
    .B(net4347),
    .Y(_03952_));
 sg13g2_a21oi_1 _18478_ (.A1(net3930),
    .A2(net4347),
    .Y(_01651_),
    .B1(_03952_));
 sg13g2_nor2_1 _18479_ (.A(net1394),
    .B(net4343),
    .Y(_03953_));
 sg13g2_a21oi_1 _18480_ (.A1(net3928),
    .A2(net4343),
    .Y(_01652_),
    .B1(_03953_));
 sg13g2_nor2_1 _18481_ (.A(net1690),
    .B(net4350),
    .Y(_03954_));
 sg13g2_a21oi_1 _18482_ (.A1(net3927),
    .A2(net4350),
    .Y(_01653_),
    .B1(_03954_));
 sg13g2_nor2_1 _18483_ (.A(net988),
    .B(net4348),
    .Y(_03955_));
 sg13g2_a21oi_1 _18484_ (.A1(net3924),
    .A2(net4348),
    .Y(_01654_),
    .B1(_03955_));
 sg13g2_nor2_1 _18485_ (.A(net1505),
    .B(net4347),
    .Y(_03956_));
 sg13g2_a21oi_1 _18486_ (.A1(net3922),
    .A2(net4347),
    .Y(_01655_),
    .B1(_03956_));
 sg13g2_nor2_1 _18487_ (.A(net1106),
    .B(net4350),
    .Y(_03957_));
 sg13g2_a21oi_1 _18488_ (.A1(net3834),
    .A2(net4349),
    .Y(_01656_),
    .B1(_03957_));
 sg13g2_nor2_1 _18489_ (.A(net1818),
    .B(net4343),
    .Y(_03958_));
 sg13g2_a21oi_1 _18490_ (.A1(net3919),
    .A2(net4343),
    .Y(_01657_),
    .B1(_03958_));
 sg13g2_nor2_1 _18491_ (.A(net1076),
    .B(net4350),
    .Y(_03959_));
 sg13g2_a21oi_1 _18492_ (.A1(net3917),
    .A2(net4350),
    .Y(_01658_),
    .B1(_03959_));
 sg13g2_nor2_1 _18493_ (.A(net1776),
    .B(net4345),
    .Y(_03960_));
 sg13g2_a21oi_1 _18494_ (.A1(net3915),
    .A2(net4345),
    .Y(_01659_),
    .B1(_03960_));
 sg13g2_nor2_1 _18495_ (.A(net1681),
    .B(net4343),
    .Y(_03961_));
 sg13g2_a21oi_1 _18496_ (.A1(net3912),
    .A2(net4343),
    .Y(_01660_),
    .B1(_03961_));
 sg13g2_nor2_1 _18497_ (.A(net1192),
    .B(net4344),
    .Y(_03962_));
 sg13g2_a21oi_1 _18498_ (.A1(net3832),
    .A2(net4344),
    .Y(_01661_),
    .B1(_03962_));
 sg13g2_nor2_1 _18499_ (.A(net1329),
    .B(net4342),
    .Y(_03963_));
 sg13g2_a21oi_1 _18500_ (.A1(net3910),
    .A2(net4342),
    .Y(_01662_),
    .B1(_03963_));
 sg13g2_nor2_1 _18501_ (.A(net1319),
    .B(net4344),
    .Y(_03964_));
 sg13g2_a21oi_1 _18502_ (.A1(net3907),
    .A2(net4344),
    .Y(_01663_),
    .B1(_03964_));
 sg13g2_nor2_1 _18503_ (.A(net1112),
    .B(net4342),
    .Y(_03965_));
 sg13g2_a21oi_1 _18504_ (.A1(net3904),
    .A2(net4342),
    .Y(_01664_),
    .B1(_03965_));
 sg13g2_nor2_1 _18505_ (.A(net1885),
    .B(net4345),
    .Y(_03966_));
 sg13g2_a21oi_1 _18506_ (.A1(net3903),
    .A2(net4345),
    .Y(_01665_),
    .B1(_03966_));
 sg13g2_nor2_1 _18507_ (.A(net1309),
    .B(net4344),
    .Y(_03967_));
 sg13g2_a21oi_1 _18508_ (.A1(net3900),
    .A2(net4344),
    .Y(_01666_),
    .B1(_03967_));
 sg13g2_nor2_1 _18509_ (.A(net1474),
    .B(net4342),
    .Y(_03968_));
 sg13g2_a21oi_1 _18510_ (.A1(net3898),
    .A2(net4342),
    .Y(_01667_),
    .B1(_03968_));
 sg13g2_nor2_1 _18511_ (.A(net1040),
    .B(net4345),
    .Y(_03969_));
 sg13g2_a21oi_1 _18512_ (.A1(net3829),
    .A2(net4345),
    .Y(_01668_),
    .B1(_03969_));
 sg13g2_nor2_1 _18513_ (.A(net1002),
    .B(net4350),
    .Y(_03970_));
 sg13g2_a21oi_1 _18514_ (.A1(net3826),
    .A2(net4350),
    .Y(_01669_),
    .B1(_03970_));
 sg13g2_nor2_1 _18515_ (.A(net1819),
    .B(net4348),
    .Y(_03971_));
 sg13g2_a21oi_1 _18516_ (.A1(net3824),
    .A2(net4348),
    .Y(_01670_),
    .B1(_03971_));
 sg13g2_nor2_1 _18517_ (.A(net1545),
    .B(net4345),
    .Y(_03972_));
 sg13g2_a21oi_1 _18518_ (.A1(net3895),
    .A2(net4346),
    .Y(_01671_),
    .B1(_03972_));
 sg13g2_nor2_1 _18519_ (.A(net1295),
    .B(net4342),
    .Y(_03973_));
 sg13g2_a21oi_1 _18520_ (.A1(net3822),
    .A2(net4342),
    .Y(_01672_),
    .B1(_03973_));
 sg13g2_nor2_1 _18521_ (.A(net1513),
    .B(net4344),
    .Y(_03974_));
 sg13g2_a21oi_1 _18522_ (.A1(net3819),
    .A2(net4344),
    .Y(_01673_),
    .B1(_03974_));
 sg13g2_nor2_1 _18523_ (.A(net1761),
    .B(net4349),
    .Y(_03975_));
 sg13g2_a21oi_1 _18524_ (.A1(net3894),
    .A2(net4349),
    .Y(_01674_),
    .B1(_03975_));
 sg13g2_nor2_1 _18525_ (.A(net1760),
    .B(net4343),
    .Y(_03976_));
 sg13g2_a21oi_1 _18526_ (.A1(net3817),
    .A2(net4343),
    .Y(_01675_),
    .B1(_03976_));
 sg13g2_nor2_2 _18527_ (.A(_03709_),
    .B(_03943_),
    .Y(_03977_));
 sg13g2_nor2_1 _18528_ (.A(net688),
    .B(net4337),
    .Y(_03978_));
 sg13g2_a21oi_1 _18529_ (.A1(net3945),
    .A2(net4337),
    .Y(_01676_),
    .B1(_03978_));
 sg13g2_nor2_1 _18530_ (.A(net1118),
    .B(net4338),
    .Y(_03979_));
 sg13g2_a21oi_1 _18531_ (.A1(net3942),
    .A2(net4338),
    .Y(_01677_),
    .B1(_03979_));
 sg13g2_nor2_1 _18532_ (.A(net831),
    .B(net4337),
    .Y(_03980_));
 sg13g2_a21oi_1 _18533_ (.A1(net3940),
    .A2(net4337),
    .Y(_01678_),
    .B1(_03980_));
 sg13g2_nor2_1 _18534_ (.A(net1452),
    .B(net4338),
    .Y(_03981_));
 sg13g2_a21oi_1 _18535_ (.A1(net3939),
    .A2(net4338),
    .Y(_01679_),
    .B1(_03981_));
 sg13g2_nor2_1 _18536_ (.A(net1456),
    .B(net4340),
    .Y(_03982_));
 sg13g2_a21oi_1 _18537_ (.A1(net3836),
    .A2(net4340),
    .Y(_01680_),
    .B1(_03982_));
 sg13g2_nor2_1 _18538_ (.A(net1041),
    .B(net4340),
    .Y(_03983_));
 sg13g2_a21oi_1 _18539_ (.A1(net3935),
    .A2(net4340),
    .Y(_01681_),
    .B1(_03983_));
 sg13g2_nor2_1 _18540_ (.A(net1747),
    .B(net4340),
    .Y(_03984_));
 sg13g2_a21oi_1 _18541_ (.A1(net3933),
    .A2(net4340),
    .Y(_01682_),
    .B1(_03984_));
 sg13g2_nor2_1 _18542_ (.A(net751),
    .B(net4338),
    .Y(_03985_));
 sg13g2_a21oi_1 _18543_ (.A1(net3930),
    .A2(net4338),
    .Y(_01683_),
    .B1(_03985_));
 sg13g2_nor2_1 _18544_ (.A(net1666),
    .B(net4333),
    .Y(_03986_));
 sg13g2_a21oi_1 _18545_ (.A1(_07305_),
    .A2(net4336),
    .Y(_01684_),
    .B1(_03986_));
 sg13g2_nor2_1 _18546_ (.A(net1336),
    .B(net4339),
    .Y(_03987_));
 sg13g2_a21oi_1 _18547_ (.A1(net3927),
    .A2(net4339),
    .Y(_01685_),
    .B1(_03987_));
 sg13g2_nor2_1 _18548_ (.A(net1186),
    .B(net4337),
    .Y(_03988_));
 sg13g2_a21oi_1 _18549_ (.A1(net3924),
    .A2(net4337),
    .Y(_01686_),
    .B1(_03988_));
 sg13g2_nor2_1 _18550_ (.A(net1125),
    .B(net4338),
    .Y(_03989_));
 sg13g2_a21oi_1 _18551_ (.A1(net3923),
    .A2(net4338),
    .Y(_01687_),
    .B1(_03989_));
 sg13g2_nor2_1 _18552_ (.A(net1150),
    .B(net4340),
    .Y(_03990_));
 sg13g2_a21oi_1 _18553_ (.A1(net3834),
    .A2(net4340),
    .Y(_01688_),
    .B1(_03990_));
 sg13g2_nor2_1 _18554_ (.A(net1088),
    .B(net4333),
    .Y(_03991_));
 sg13g2_a21oi_1 _18555_ (.A1(net3919),
    .A2(net4333),
    .Y(_01689_),
    .B1(_03991_));
 sg13g2_nor2_1 _18556_ (.A(net1039),
    .B(net4339),
    .Y(_03992_));
 sg13g2_a21oi_1 _18557_ (.A1(net3918),
    .A2(net4339),
    .Y(_01690_),
    .B1(_03992_));
 sg13g2_nor2_1 _18558_ (.A(net1943),
    .B(net4335),
    .Y(_03993_));
 sg13g2_a21oi_1 _18559_ (.A1(net3916),
    .A2(net4335),
    .Y(_01691_),
    .B1(_03993_));
 sg13g2_nor2_1 _18560_ (.A(net1797),
    .B(net4332),
    .Y(_03994_));
 sg13g2_a21oi_1 _18561_ (.A1(net3911),
    .A2(net4332),
    .Y(_01692_),
    .B1(_03994_));
 sg13g2_nor2_1 _18562_ (.A(net1811),
    .B(net4334),
    .Y(_03995_));
 sg13g2_a21oi_1 _18563_ (.A1(net3831),
    .A2(net4334),
    .Y(_01693_),
    .B1(_03995_));
 sg13g2_nor2_1 _18564_ (.A(net1414),
    .B(net4332),
    .Y(_03996_));
 sg13g2_a21oi_1 _18565_ (.A1(net3909),
    .A2(net4332),
    .Y(_01694_),
    .B1(_03996_));
 sg13g2_nor2_1 _18566_ (.A(net1965),
    .B(net4334),
    .Y(_03997_));
 sg13g2_a21oi_1 _18567_ (.A1(net3906),
    .A2(net4334),
    .Y(_01695_),
    .B1(_03997_));
 sg13g2_nor2_1 _18568_ (.A(net1643),
    .B(net4333),
    .Y(_03998_));
 sg13g2_a21oi_1 _18569_ (.A1(net3904),
    .A2(net4333),
    .Y(_01696_),
    .B1(_03998_));
 sg13g2_nor2_1 _18570_ (.A(net1673),
    .B(net4334),
    .Y(_03999_));
 sg13g2_a21oi_1 _18571_ (.A1(net3903),
    .A2(net4334),
    .Y(_01697_),
    .B1(_03999_));
 sg13g2_nor2_1 _18572_ (.A(net1006),
    .B(net4334),
    .Y(_04000_));
 sg13g2_a21oi_1 _18573_ (.A1(net3900),
    .A2(net4334),
    .Y(_01698_),
    .B1(_04000_));
 sg13g2_nor2_1 _18574_ (.A(net1463),
    .B(net4332),
    .Y(_04001_));
 sg13g2_a21oi_1 _18575_ (.A1(net3897),
    .A2(net4332),
    .Y(_01699_),
    .B1(_04001_));
 sg13g2_nor2_1 _18576_ (.A(net1087),
    .B(net4335),
    .Y(_04002_));
 sg13g2_a21oi_1 _18577_ (.A1(net3829),
    .A2(net4335),
    .Y(_01700_),
    .B1(_04002_));
 sg13g2_nor2_1 _18578_ (.A(net1844),
    .B(net4339),
    .Y(_04003_));
 sg13g2_a21oi_1 _18579_ (.A1(net3826),
    .A2(net4339),
    .Y(_01701_),
    .B1(_04003_));
 sg13g2_nor2_1 _18580_ (.A(net2053),
    .B(net4337),
    .Y(_04004_));
 sg13g2_a21oi_1 _18581_ (.A1(net3825),
    .A2(net4337),
    .Y(_01702_),
    .B1(_04004_));
 sg13g2_nor2_1 _18582_ (.A(net1956),
    .B(net4335),
    .Y(_04005_));
 sg13g2_a21oi_1 _18583_ (.A1(net3895),
    .A2(net4335),
    .Y(_01703_),
    .B1(_04005_));
 sg13g2_nor2_1 _18584_ (.A(net765),
    .B(net4332),
    .Y(_04006_));
 sg13g2_a21oi_1 _18585_ (.A1(net3821),
    .A2(net4332),
    .Y(_01704_),
    .B1(_04006_));
 sg13g2_nor2_1 _18586_ (.A(net1092),
    .B(net4335),
    .Y(_04007_));
 sg13g2_a21oi_1 _18587_ (.A1(net3820),
    .A2(net4335),
    .Y(_01705_),
    .B1(_04007_));
 sg13g2_nor2_1 _18588_ (.A(net1010),
    .B(net4339),
    .Y(_04008_));
 sg13g2_a21oi_1 _18589_ (.A1(net3894),
    .A2(net4339),
    .Y(_01706_),
    .B1(_04008_));
 sg13g2_nor2_1 _18590_ (.A(net1430),
    .B(net4333),
    .Y(_04009_));
 sg13g2_a21oi_1 _18591_ (.A1(net3817),
    .A2(net4333),
    .Y(_01707_),
    .B1(_04009_));
 sg13g2_nor2_1 _18592_ (.A(_03743_),
    .B(_03943_),
    .Y(_04010_));
 sg13g2_nor2_1 _18593_ (.A(net1800),
    .B(net4328),
    .Y(_04011_));
 sg13g2_a21oi_1 _18594_ (.A1(net3944),
    .A2(net4328),
    .Y(_01708_),
    .B1(_04011_));
 sg13g2_nor2_1 _18595_ (.A(net829),
    .B(net4326),
    .Y(_04012_));
 sg13g2_a21oi_1 _18596_ (.A1(net3943),
    .A2(net4326),
    .Y(_01709_),
    .B1(_04012_));
 sg13g2_nor2_1 _18597_ (.A(net845),
    .B(net4327),
    .Y(_04013_));
 sg13g2_a21oi_1 _18598_ (.A1(net3940),
    .A2(net4327),
    .Y(_01710_),
    .B1(_04013_));
 sg13g2_nor2_1 _18599_ (.A(net1593),
    .B(net4326),
    .Y(_04014_));
 sg13g2_a21oi_1 _18600_ (.A1(net3938),
    .A2(net4326),
    .Y(_01711_),
    .B1(_04014_));
 sg13g2_nor2_1 _18601_ (.A(net1055),
    .B(net4330),
    .Y(_04015_));
 sg13g2_a21oi_1 _18602_ (.A1(net3835),
    .A2(net4330),
    .Y(_01712_),
    .B1(_04015_));
 sg13g2_nor2_1 _18603_ (.A(net726),
    .B(net4327),
    .Y(_04016_));
 sg13g2_a21oi_1 _18604_ (.A1(net3937),
    .A2(net4327),
    .Y(_01713_),
    .B1(_04016_));
 sg13g2_nor2_1 _18605_ (.A(net991),
    .B(net4330),
    .Y(_04017_));
 sg13g2_a21oi_1 _18606_ (.A1(net3934),
    .A2(net4330),
    .Y(_01714_),
    .B1(_04017_));
 sg13g2_nor2_1 _18607_ (.A(net1001),
    .B(net4326),
    .Y(_04018_));
 sg13g2_a21oi_1 _18608_ (.A1(net3930),
    .A2(net4326),
    .Y(_01715_),
    .B1(_04018_));
 sg13g2_nor2_1 _18609_ (.A(net1050),
    .B(net4323),
    .Y(_04019_));
 sg13g2_a21oi_1 _18610_ (.A1(net3929),
    .A2(net4331),
    .Y(_01716_),
    .B1(_04019_));
 sg13g2_nor2_1 _18611_ (.A(net1385),
    .B(net4329),
    .Y(_04020_));
 sg13g2_a21oi_1 _18612_ (.A1(net3927),
    .A2(net4329),
    .Y(_01717_),
    .B1(_04020_));
 sg13g2_nor2_1 _18613_ (.A(net1633),
    .B(net4328),
    .Y(_04021_));
 sg13g2_a21oi_1 _18614_ (.A1(net3924),
    .A2(net4328),
    .Y(_01718_),
    .B1(_04021_));
 sg13g2_nor2_1 _18615_ (.A(net1536),
    .B(net4326),
    .Y(_04022_));
 sg13g2_a21oi_1 _18616_ (.A1(net3922),
    .A2(net4326),
    .Y(_01719_),
    .B1(_04022_));
 sg13g2_nor2_1 _18617_ (.A(net1135),
    .B(net4331),
    .Y(_04023_));
 sg13g2_a21oi_1 _18618_ (.A1(net3833),
    .A2(net4330),
    .Y(_01720_),
    .B1(_04023_));
 sg13g2_nor2_1 _18619_ (.A(net1429),
    .B(net4323),
    .Y(_04024_));
 sg13g2_a21oi_1 _18620_ (.A1(net3919),
    .A2(net4323),
    .Y(_01721_),
    .B1(_04024_));
 sg13g2_nor2_1 _18621_ (.A(net923),
    .B(net4330),
    .Y(_04025_));
 sg13g2_a21oi_1 _18622_ (.A1(net3918),
    .A2(net4330),
    .Y(_01722_),
    .B1(_04025_));
 sg13g2_nor2_1 _18623_ (.A(net1015),
    .B(net4325),
    .Y(_04026_));
 sg13g2_a21oi_1 _18624_ (.A1(net3914),
    .A2(net4325),
    .Y(_01723_),
    .B1(_04026_));
 sg13g2_nor2_1 _18625_ (.A(net1363),
    .B(net4322),
    .Y(_04027_));
 sg13g2_a21oi_1 _18626_ (.A1(net3911),
    .A2(net4322),
    .Y(_01724_),
    .B1(_04027_));
 sg13g2_nor2_1 _18627_ (.A(net1627),
    .B(net4324),
    .Y(_04028_));
 sg13g2_a21oi_1 _18628_ (.A1(net3832),
    .A2(net4324),
    .Y(_01725_),
    .B1(_04028_));
 sg13g2_nor2_1 _18629_ (.A(net1318),
    .B(net4322),
    .Y(_04029_));
 sg13g2_a21oi_1 _18630_ (.A1(net3910),
    .A2(net4322),
    .Y(_01726_),
    .B1(_04029_));
 sg13g2_nor2_1 _18631_ (.A(net1931),
    .B(net4324),
    .Y(_04030_));
 sg13g2_a21oi_1 _18632_ (.A1(net3906),
    .A2(net4324),
    .Y(_01727_),
    .B1(_04030_));
 sg13g2_nor2_1 _18633_ (.A(net1083),
    .B(net4322),
    .Y(_04031_));
 sg13g2_a21oi_1 _18634_ (.A1(net3905),
    .A2(net4323),
    .Y(_01728_),
    .B1(_04031_));
 sg13g2_nor2_1 _18635_ (.A(net1044),
    .B(net4325),
    .Y(_04032_));
 sg13g2_a21oi_1 _18636_ (.A1(net3903),
    .A2(net4324),
    .Y(_01729_),
    .B1(_04032_));
 sg13g2_nor2_1 _18637_ (.A(net698),
    .B(net4324),
    .Y(_04033_));
 sg13g2_a21oi_1 _18638_ (.A1(net3900),
    .A2(net4324),
    .Y(_01730_),
    .B1(_04033_));
 sg13g2_nor2_1 _18639_ (.A(net686),
    .B(net4322),
    .Y(_04034_));
 sg13g2_a21oi_1 _18640_ (.A1(net3898),
    .A2(net4322),
    .Y(_01731_),
    .B1(_04034_));
 sg13g2_nor2_1 _18641_ (.A(net997),
    .B(net4329),
    .Y(_04035_));
 sg13g2_a21oi_1 _18642_ (.A1(net3830),
    .A2(net4329),
    .Y(_01732_),
    .B1(_04035_));
 sg13g2_nor2_1 _18643_ (.A(net804),
    .B(net4329),
    .Y(_04036_));
 sg13g2_a21oi_1 _18644_ (.A1(net3826),
    .A2(net4329),
    .Y(_01733_),
    .B1(_04036_));
 sg13g2_nor2_1 _18645_ (.A(net1084),
    .B(net4328),
    .Y(_04037_));
 sg13g2_a21oi_1 _18646_ (.A1(net3825),
    .A2(net4328),
    .Y(_01734_),
    .B1(_04037_));
 sg13g2_nor2_1 _18647_ (.A(net716),
    .B(net4325),
    .Y(_04038_));
 sg13g2_a21oi_1 _18648_ (.A1(net3896),
    .A2(net4325),
    .Y(_01735_),
    .B1(_04038_));
 sg13g2_nor2_1 _18649_ (.A(net840),
    .B(net4322),
    .Y(_04039_));
 sg13g2_a21oi_1 _18650_ (.A1(net3821),
    .A2(net4323),
    .Y(_01736_),
    .B1(_04039_));
 sg13g2_nor2_1 _18651_ (.A(net1371),
    .B(net4325),
    .Y(_04040_));
 sg13g2_a21oi_1 _18652_ (.A1(net3819),
    .A2(net4324),
    .Y(_01737_),
    .B1(_04040_));
 sg13g2_nor2_1 _18653_ (.A(net1008),
    .B(net4329),
    .Y(_04041_));
 sg13g2_a21oi_1 _18654_ (.A1(net3893),
    .A2(net4329),
    .Y(_01738_),
    .B1(_04041_));
 sg13g2_nor2_1 _18655_ (.A(net1177),
    .B(net4323),
    .Y(_04042_));
 sg13g2_a21oi_1 _18656_ (.A1(net3817),
    .A2(net4323),
    .Y(_01739_),
    .B1(_04042_));
 sg13g2_nor4_1 _18657_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .C(_05481_),
    .D(_03943_),
    .Y(_04043_));
 sg13g2_nor2_1 _18658_ (.A(net907),
    .B(net4318),
    .Y(_04044_));
 sg13g2_a21oi_1 _18659_ (.A1(net3945),
    .A2(net4318),
    .Y(_01740_),
    .B1(_04044_));
 sg13g2_nor2_1 _18660_ (.A(net1538),
    .B(net4316),
    .Y(_04045_));
 sg13g2_a21oi_1 _18661_ (.A1(net3942),
    .A2(net4316),
    .Y(_01741_),
    .B1(_04045_));
 sg13g2_nor2_1 _18662_ (.A(net1153),
    .B(net4317),
    .Y(_04046_));
 sg13g2_a21oi_1 _18663_ (.A1(net3941),
    .A2(net4317),
    .Y(_01742_),
    .B1(_04046_));
 sg13g2_nor2_1 _18664_ (.A(net1824),
    .B(net4316),
    .Y(_04047_));
 sg13g2_a21oi_1 _18665_ (.A1(net3939),
    .A2(net4316),
    .Y(_01743_),
    .B1(_04047_));
 sg13g2_nor2_1 _18666_ (.A(net1543),
    .B(net4320),
    .Y(_04048_));
 sg13g2_a21oi_1 _18667_ (.A1(net3836),
    .A2(net4320),
    .Y(_01744_),
    .B1(_04048_));
 sg13g2_nor2_1 _18668_ (.A(net1028),
    .B(net4317),
    .Y(_04049_));
 sg13g2_a21oi_1 _18669_ (.A1(net3936),
    .A2(net4317),
    .Y(_01745_),
    .B1(_04049_));
 sg13g2_nor2_1 _18670_ (.A(net1507),
    .B(net4320),
    .Y(_04050_));
 sg13g2_a21oi_1 _18671_ (.A1(net3933),
    .A2(net4320),
    .Y(_01746_),
    .B1(_04050_));
 sg13g2_nor2_1 _18672_ (.A(net1481),
    .B(net4316),
    .Y(_04051_));
 sg13g2_a21oi_1 _18673_ (.A1(net3930),
    .A2(net4316),
    .Y(_01747_),
    .B1(_04051_));
 sg13g2_nor2_1 _18674_ (.A(net1221),
    .B(net4312),
    .Y(_04052_));
 sg13g2_a21oi_1 _18675_ (.A1(net3928),
    .A2(net4312),
    .Y(_01748_),
    .B1(_04052_));
 sg13g2_nor2_1 _18676_ (.A(net908),
    .B(net4319),
    .Y(_04053_));
 sg13g2_a21oi_1 _18677_ (.A1(net3926),
    .A2(net4319),
    .Y(_01749_),
    .B1(_04053_));
 sg13g2_nor2_1 _18678_ (.A(net1764),
    .B(net4318),
    .Y(_04054_));
 sg13g2_a21oi_1 _18679_ (.A1(net3924),
    .A2(net4318),
    .Y(_01750_),
    .B1(_04054_));
 sg13g2_nor2_1 _18680_ (.A(net1327),
    .B(net4316),
    .Y(_04055_));
 sg13g2_a21oi_1 _18681_ (.A1(net3923),
    .A2(net4316),
    .Y(_01751_),
    .B1(_04055_));
 sg13g2_nor2_1 _18682_ (.A(net1152),
    .B(net4319),
    .Y(_04056_));
 sg13g2_a21oi_1 _18683_ (.A1(net3833),
    .A2(net4319),
    .Y(_01752_),
    .B1(_04056_));
 sg13g2_nor2_1 _18684_ (.A(net1059),
    .B(net4312),
    .Y(_04057_));
 sg13g2_a21oi_1 _18685_ (.A1(net3920),
    .A2(net4312),
    .Y(_01753_),
    .B1(_04057_));
 sg13g2_nor2_1 _18686_ (.A(net1443),
    .B(net4319),
    .Y(_04058_));
 sg13g2_a21oi_1 _18687_ (.A1(net3917),
    .A2(net4319),
    .Y(_01754_),
    .B1(_04058_));
 sg13g2_nor2_1 _18688_ (.A(net1863),
    .B(net4314),
    .Y(_04059_));
 sg13g2_a21oi_1 _18689_ (.A1(net3915),
    .A2(net4314),
    .Y(_01755_),
    .B1(_04059_));
 sg13g2_nor2_1 _18690_ (.A(net1782),
    .B(net4312),
    .Y(_04060_));
 sg13g2_a21oi_1 _18691_ (.A1(net3912),
    .A2(net4312),
    .Y(_01756_),
    .B1(_04060_));
 sg13g2_nor2_1 _18692_ (.A(net2010),
    .B(net4313),
    .Y(_04061_));
 sg13g2_a21oi_1 _18693_ (.A1(net3831),
    .A2(net4313),
    .Y(_01757_),
    .B1(_04061_));
 sg13g2_nor2_1 _18694_ (.A(net1862),
    .B(net4311),
    .Y(_04062_));
 sg13g2_a21oi_1 _18695_ (.A1(net3910),
    .A2(net4311),
    .Y(_01758_),
    .B1(_04062_));
 sg13g2_nor2_1 _18696_ (.A(net1472),
    .B(net4313),
    .Y(_04063_));
 sg13g2_a21oi_1 _18697_ (.A1(net3906),
    .A2(net4313),
    .Y(_01759_),
    .B1(_04063_));
 sg13g2_nor2_1 _18698_ (.A(net2191),
    .B(net4311),
    .Y(_04064_));
 sg13g2_a21oi_1 _18699_ (.A1(net3905),
    .A2(net4311),
    .Y(_01760_),
    .B1(_04064_));
 sg13g2_nor2_1 _18700_ (.A(net1220),
    .B(net4313),
    .Y(_04065_));
 sg13g2_a21oi_1 _18701_ (.A1(net3902),
    .A2(net4313),
    .Y(_01761_),
    .B1(_04065_));
 sg13g2_nor2_1 _18702_ (.A(net1522),
    .B(net4313),
    .Y(_04066_));
 sg13g2_a21oi_1 _18703_ (.A1(net3900),
    .A2(net4313),
    .Y(_01762_),
    .B1(_04066_));
 sg13g2_nor2_1 _18704_ (.A(net820),
    .B(net4311),
    .Y(_04067_));
 sg13g2_a21oi_1 _18705_ (.A1(net3899),
    .A2(net4311),
    .Y(_01763_),
    .B1(_04067_));
 sg13g2_nor2_1 _18706_ (.A(net951),
    .B(net4314),
    .Y(_04068_));
 sg13g2_a21oi_1 _18707_ (.A1(net3830),
    .A2(net4314),
    .Y(_01764_),
    .B1(_04068_));
 sg13g2_nor2_1 _18708_ (.A(net1479),
    .B(net4319),
    .Y(_04069_));
 sg13g2_a21oi_1 _18709_ (.A1(net3827),
    .A2(net4319),
    .Y(_01765_),
    .B1(_04069_));
 sg13g2_nor2_1 _18710_ (.A(net1675),
    .B(net4318),
    .Y(_04070_));
 sg13g2_a21oi_1 _18711_ (.A1(net3825),
    .A2(net4318),
    .Y(_01766_),
    .B1(_04070_));
 sg13g2_nor2_1 _18712_ (.A(net1717),
    .B(net4314),
    .Y(_04071_));
 sg13g2_a21oi_1 _18713_ (.A1(net3896),
    .A2(net4314),
    .Y(_01767_),
    .B1(_04071_));
 sg13g2_nor2_1 _18714_ (.A(net1708),
    .B(net4311),
    .Y(_04072_));
 sg13g2_a21oi_1 _18715_ (.A1(net3823),
    .A2(net4311),
    .Y(_01768_),
    .B1(_04072_));
 sg13g2_nor2_1 _18716_ (.A(net787),
    .B(net4314),
    .Y(_04073_));
 sg13g2_a21oi_1 _18717_ (.A1(net3820),
    .A2(net4314),
    .Y(_01769_),
    .B1(_04073_));
 sg13g2_nor2_1 _18718_ (.A(net1121),
    .B(net4320),
    .Y(_04074_));
 sg13g2_a21oi_1 _18719_ (.A1(net3894),
    .A2(net4320),
    .Y(_01770_),
    .B1(_04074_));
 sg13g2_nor2_1 _18720_ (.A(net1051),
    .B(net4312),
    .Y(_04075_));
 sg13g2_a21oi_1 _18721_ (.A1(net3818),
    .A2(net4312),
    .Y(_01771_),
    .B1(_04075_));
 sg13g2_nor3_2 _18722_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .C(_07212_),
    .Y(_04076_));
 sg13g2_nor2_1 _18723_ (.A(net1444),
    .B(net4307),
    .Y(_04077_));
 sg13g2_a21oi_1 _18724_ (.A1(net3944),
    .A2(net4307),
    .Y(_01772_),
    .B1(_04077_));
 sg13g2_nor2_1 _18725_ (.A(net1549),
    .B(net4306),
    .Y(_04078_));
 sg13g2_a21oi_1 _18726_ (.A1(net3943),
    .A2(net4306),
    .Y(_01773_),
    .B1(_04078_));
 sg13g2_nor2_1 _18727_ (.A(net1727),
    .B(net4306),
    .Y(_04079_));
 sg13g2_a21oi_1 _18728_ (.A1(net3941),
    .A2(net4307),
    .Y(_01774_),
    .B1(_04079_));
 sg13g2_nor2_1 _18729_ (.A(net1795),
    .B(net4306),
    .Y(_04080_));
 sg13g2_a21oi_1 _18730_ (.A1(net3938),
    .A2(net4306),
    .Y(_01775_),
    .B1(_04080_));
 sg13g2_nor2_1 _18731_ (.A(net922),
    .B(net4308),
    .Y(_04081_));
 sg13g2_a21oi_1 _18732_ (.A1(net3835),
    .A2(net4308),
    .Y(_01776_),
    .B1(_04081_));
 sg13g2_nor2_1 _18733_ (.A(net1353),
    .B(net4308),
    .Y(_04082_));
 sg13g2_a21oi_1 _18734_ (.A1(net3936),
    .A2(net4310),
    .Y(_01777_),
    .B1(_04082_));
 sg13g2_nor2_1 _18735_ (.A(net699),
    .B(net4308),
    .Y(_04083_));
 sg13g2_a21oi_1 _18736_ (.A1(net3932),
    .A2(net4308),
    .Y(_01778_),
    .B1(_04083_));
 sg13g2_nor2_1 _18737_ (.A(net987),
    .B(net4310),
    .Y(_04084_));
 sg13g2_a21oi_1 _18738_ (.A1(net3931),
    .A2(net4306),
    .Y(_01779_),
    .B1(_04084_));
 sg13g2_nor2_1 _18739_ (.A(net1298),
    .B(net4302),
    .Y(_04085_));
 sg13g2_a21oi_1 _18740_ (.A1(net3928),
    .A2(net4302),
    .Y(_01780_),
    .B1(_04085_));
 sg13g2_nor2_1 _18741_ (.A(net1484),
    .B(net4309),
    .Y(_04086_));
 sg13g2_a21oi_1 _18742_ (.A1(net3927),
    .A2(net4309),
    .Y(_01781_),
    .B1(_04086_));
 sg13g2_nor2_1 _18743_ (.A(net1264),
    .B(net4307),
    .Y(_04087_));
 sg13g2_a21oi_1 _18744_ (.A1(net3924),
    .A2(net4307),
    .Y(_01782_),
    .B1(_04087_));
 sg13g2_nor2_1 _18745_ (.A(net2021),
    .B(net4306),
    .Y(_04088_));
 sg13g2_a21oi_1 _18746_ (.A1(net3922),
    .A2(net4306),
    .Y(_01783_),
    .B1(_04088_));
 sg13g2_nor2_1 _18747_ (.A(net1007),
    .B(net4308),
    .Y(_04089_));
 sg13g2_a21oi_1 _18748_ (.A1(net3834),
    .A2(net4309),
    .Y(_01784_),
    .B1(_04089_));
 sg13g2_nor2_1 _18749_ (.A(net1042),
    .B(net4302),
    .Y(_04090_));
 sg13g2_a21oi_1 _18750_ (.A1(net3919),
    .A2(net4302),
    .Y(_01785_),
    .B1(_04090_));
 sg13g2_nor2_1 _18751_ (.A(net1662),
    .B(net4309),
    .Y(_04091_));
 sg13g2_a21oi_1 _18752_ (.A1(net3918),
    .A2(net4309),
    .Y(_01786_),
    .B1(_04091_));
 sg13g2_nor2_1 _18753_ (.A(net966),
    .B(net4304),
    .Y(_04092_));
 sg13g2_a21oi_1 _18754_ (.A1(net3914),
    .A2(net4304),
    .Y(_01787_),
    .B1(_04092_));
 sg13g2_nor2_1 _18755_ (.A(net1519),
    .B(net4302),
    .Y(_04093_));
 sg13g2_a21oi_1 _18756_ (.A1(net3912),
    .A2(net4302),
    .Y(_01788_),
    .B1(_04093_));
 sg13g2_nor2_1 _18757_ (.A(net1143),
    .B(net4303),
    .Y(_04094_));
 sg13g2_a21oi_1 _18758_ (.A1(net3831),
    .A2(net4303),
    .Y(_01789_),
    .B1(_04094_));
 sg13g2_nor2_1 _18759_ (.A(net1682),
    .B(net4301),
    .Y(_04095_));
 sg13g2_a21oi_1 _18760_ (.A1(net3909),
    .A2(net4301),
    .Y(_01790_),
    .B1(_04095_));
 sg13g2_nor2_1 _18761_ (.A(net823),
    .B(net4303),
    .Y(_04096_));
 sg13g2_a21oi_1 _18762_ (.A1(net3908),
    .A2(net4303),
    .Y(_01791_),
    .B1(_04096_));
 sg13g2_nor2_1 _18763_ (.A(net1077),
    .B(net4301),
    .Y(_04097_));
 sg13g2_a21oi_1 _18764_ (.A1(net3905),
    .A2(net4301),
    .Y(_01792_),
    .B1(_04097_));
 sg13g2_nor2_1 _18765_ (.A(net796),
    .B(net4303),
    .Y(_04098_));
 sg13g2_a21oi_1 _18766_ (.A1(net3902),
    .A2(net4303),
    .Y(_01793_),
    .B1(_04098_));
 sg13g2_nor2_1 _18767_ (.A(net965),
    .B(net4303),
    .Y(_04099_));
 sg13g2_a21oi_1 _18768_ (.A1(net3901),
    .A2(net4303),
    .Y(_01794_),
    .B1(_04099_));
 sg13g2_nor2_1 _18769_ (.A(net1945),
    .B(net4301),
    .Y(_04100_));
 sg13g2_a21oi_1 _18770_ (.A1(net3897),
    .A2(net4301),
    .Y(_01795_),
    .B1(_04100_));
 sg13g2_nor2_1 _18771_ (.A(net1471),
    .B(net4304),
    .Y(_04101_));
 sg13g2_a21oi_1 _18772_ (.A1(_07468_),
    .A2(net4304),
    .Y(_01796_),
    .B1(_04101_));
 sg13g2_nor2_1 _18773_ (.A(net1771),
    .B(net4309),
    .Y(_04102_));
 sg13g2_a21oi_1 _18774_ (.A1(net3826),
    .A2(net4309),
    .Y(_01797_),
    .B1(_04102_));
 sg13g2_nor2_1 _18775_ (.A(net1823),
    .B(net4307),
    .Y(_04103_));
 sg13g2_a21oi_1 _18776_ (.A1(net3825),
    .A2(net4307),
    .Y(_01798_),
    .B1(_04103_));
 sg13g2_nor2_1 _18777_ (.A(net1254),
    .B(net4304),
    .Y(_04104_));
 sg13g2_a21oi_1 _18778_ (.A1(net3895),
    .A2(net4304),
    .Y(_01799_),
    .B1(_04104_));
 sg13g2_nor2_1 _18779_ (.A(net1270),
    .B(net4301),
    .Y(_04105_));
 sg13g2_a21oi_1 _18780_ (.A1(net3821),
    .A2(net4301),
    .Y(_01800_),
    .B1(_04105_));
 sg13g2_nor2_1 _18781_ (.A(net625),
    .B(net4304),
    .Y(_04106_));
 sg13g2_a21oi_1 _18782_ (.A1(net3820),
    .A2(net4304),
    .Y(_01801_),
    .B1(_04106_));
 sg13g2_nor2_1 _18783_ (.A(net1424),
    .B(net4308),
    .Y(_04107_));
 sg13g2_a21oi_1 _18784_ (.A1(net3894),
    .A2(net4308),
    .Y(_01802_),
    .B1(_04107_));
 sg13g2_nor2_1 _18785_ (.A(net1324),
    .B(net4302),
    .Y(_04108_));
 sg13g2_a21oi_1 _18786_ (.A1(net3817),
    .A2(net4302),
    .Y(_01803_),
    .B1(_04108_));
 sg13g2_nor3_2 _18787_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .C(_03709_),
    .Y(_04109_));
 sg13g2_nor2_1 _18788_ (.A(net865),
    .B(net4297),
    .Y(_04110_));
 sg13g2_a21oi_1 _18789_ (.A1(net3945),
    .A2(net4297),
    .Y(_01804_),
    .B1(_04110_));
 sg13g2_nor2_1 _18790_ (.A(net1562),
    .B(net4300),
    .Y(_04111_));
 sg13g2_a21oi_1 _18791_ (.A1(net3942),
    .A2(net4296),
    .Y(_01805_),
    .B1(_04111_));
 sg13g2_nor2_1 _18792_ (.A(net815),
    .B(net4297),
    .Y(_04112_));
 sg13g2_a21oi_1 _18793_ (.A1(net3941),
    .A2(net4297),
    .Y(_01806_),
    .B1(_04112_));
 sg13g2_nor2_1 _18794_ (.A(net1651),
    .B(net4296),
    .Y(_04113_));
 sg13g2_a21oi_1 _18795_ (.A1(net3939),
    .A2(net4296),
    .Y(_01807_),
    .B1(_04113_));
 sg13g2_nor2_1 _18796_ (.A(net1215),
    .B(net4298),
    .Y(_04114_));
 sg13g2_a21oi_1 _18797_ (.A1(net3836),
    .A2(net4298),
    .Y(_01808_),
    .B1(_04114_));
 sg13g2_nor2_1 _18798_ (.A(net1736),
    .B(net4298),
    .Y(_04115_));
 sg13g2_a21oi_1 _18799_ (.A1(net3935),
    .A2(net4296),
    .Y(_01809_),
    .B1(_04115_));
 sg13g2_nor2_1 _18800_ (.A(net1358),
    .B(net4298),
    .Y(_04116_));
 sg13g2_a21oi_1 _18801_ (.A1(net3932),
    .A2(net4298),
    .Y(_01810_),
    .B1(_04116_));
 sg13g2_nor2_1 _18802_ (.A(net1141),
    .B(net4296),
    .Y(_04117_));
 sg13g2_a21oi_1 _18803_ (.A1(net3930),
    .A2(net4296),
    .Y(_01811_),
    .B1(_04117_));
 sg13g2_nor2_1 _18804_ (.A(net1079),
    .B(net4292),
    .Y(_04118_));
 sg13g2_a21oi_1 _18805_ (.A1(net3929),
    .A2(net4292),
    .Y(_01812_),
    .B1(_04118_));
 sg13g2_nor2_1 _18806_ (.A(net983),
    .B(net4299),
    .Y(_04119_));
 sg13g2_a21oi_1 _18807_ (.A1(net3926),
    .A2(net4299),
    .Y(_01813_),
    .B1(_04119_));
 sg13g2_nor2_1 _18808_ (.A(net844),
    .B(net4297),
    .Y(_04120_));
 sg13g2_a21oi_1 _18809_ (.A1(net3925),
    .A2(net4297),
    .Y(_01814_),
    .B1(_04120_));
 sg13g2_nor2_1 _18810_ (.A(net1354),
    .B(net4296),
    .Y(_04121_));
 sg13g2_a21oi_1 _18811_ (.A1(net3922),
    .A2(net4296),
    .Y(_01815_),
    .B1(_04121_));
 sg13g2_nor2_1 _18812_ (.A(net899),
    .B(net4298),
    .Y(_04122_));
 sg13g2_a21oi_1 _18813_ (.A1(net3834),
    .A2(net4299),
    .Y(_01816_),
    .B1(_04122_));
 sg13g2_nor2_1 _18814_ (.A(net1423),
    .B(net4292),
    .Y(_04123_));
 sg13g2_a21oi_1 _18815_ (.A1(net3921),
    .A2(net4292),
    .Y(_01817_),
    .B1(_04123_));
 sg13g2_nor2_1 _18816_ (.A(net1018),
    .B(net4299),
    .Y(_04124_));
 sg13g2_a21oi_1 _18817_ (.A1(net3918),
    .A2(net4299),
    .Y(_01818_),
    .B1(_04124_));
 sg13g2_nor2_1 _18818_ (.A(net1229),
    .B(net4294),
    .Y(_04125_));
 sg13g2_a21oi_1 _18819_ (.A1(net3915),
    .A2(net4294),
    .Y(_01819_),
    .B1(_04125_));
 sg13g2_nor2_1 _18820_ (.A(net735),
    .B(net4291),
    .Y(_04126_));
 sg13g2_a21oi_1 _18821_ (.A1(net3911),
    .A2(net4291),
    .Y(_01820_),
    .B1(_04126_));
 sg13g2_nor2_1 _18822_ (.A(net1794),
    .B(net4293),
    .Y(_04127_));
 sg13g2_a21oi_1 _18823_ (.A1(net3832),
    .A2(net4293),
    .Y(_01821_),
    .B1(_04127_));
 sg13g2_nor2_1 _18824_ (.A(net1374),
    .B(net4291),
    .Y(_04128_));
 sg13g2_a21oi_1 _18825_ (.A1(net3910),
    .A2(net4291),
    .Y(_01822_),
    .B1(_04128_));
 sg13g2_nor2_1 _18826_ (.A(net1546),
    .B(net4293),
    .Y(_04129_));
 sg13g2_a21oi_1 _18827_ (.A1(net3907),
    .A2(net4293),
    .Y(_01823_),
    .B1(_04129_));
 sg13g2_nor2_1 _18828_ (.A(net1451),
    .B(net4291),
    .Y(_04130_));
 sg13g2_a21oi_1 _18829_ (.A1(net3905),
    .A2(net4291),
    .Y(_01824_),
    .B1(_04130_));
 sg13g2_nor2_1 _18830_ (.A(net1260),
    .B(net4293),
    .Y(_04131_));
 sg13g2_a21oi_1 _18831_ (.A1(net3903),
    .A2(net4293),
    .Y(_01825_),
    .B1(_04131_));
 sg13g2_nor2_1 _18832_ (.A(net1378),
    .B(net4293),
    .Y(_04132_));
 sg13g2_a21oi_1 _18833_ (.A1(net3900),
    .A2(net4293),
    .Y(_01826_),
    .B1(_04132_));
 sg13g2_nor2_1 _18834_ (.A(net2111),
    .B(net4291),
    .Y(_04133_));
 sg13g2_a21oi_1 _18835_ (.A1(net3898),
    .A2(net4291),
    .Y(_01827_),
    .B1(_04133_));
 sg13g2_nor2_1 _18836_ (.A(net1241),
    .B(net4294),
    .Y(_04134_));
 sg13g2_a21oi_1 _18837_ (.A1(net3829),
    .A2(net4294),
    .Y(_01828_),
    .B1(_04134_));
 sg13g2_nor2_1 _18838_ (.A(net1052),
    .B(net4299),
    .Y(_04135_));
 sg13g2_a21oi_1 _18839_ (.A1(net3827),
    .A2(net4299),
    .Y(_01829_),
    .B1(_04135_));
 sg13g2_nor2_1 _18840_ (.A(net909),
    .B(net4297),
    .Y(_04136_));
 sg13g2_a21oi_1 _18841_ (.A1(net3825),
    .A2(net4297),
    .Y(_01830_),
    .B1(_04136_));
 sg13g2_nor2_1 _18842_ (.A(net1255),
    .B(net4294),
    .Y(_04137_));
 sg13g2_a21oi_1 _18843_ (.A1(net3896),
    .A2(net4294),
    .Y(_01831_),
    .B1(_04137_));
 sg13g2_nor2_1 _18844_ (.A(net684),
    .B(net4292),
    .Y(_04138_));
 sg13g2_a21oi_1 _18845_ (.A1(net3821),
    .A2(net4292),
    .Y(_01832_),
    .B1(_04138_));
 sg13g2_nor2_1 _18846_ (.A(net927),
    .B(net4294),
    .Y(_04139_));
 sg13g2_a21oi_1 _18847_ (.A1(net3820),
    .A2(net4294),
    .Y(_01833_),
    .B1(_04139_));
 sg13g2_nor2_1 _18848_ (.A(net2340),
    .B(net4298),
    .Y(_04140_));
 sg13g2_a21oi_1 _18849_ (.A1(net3894),
    .A2(net4298),
    .Y(_01834_),
    .B1(_04140_));
 sg13g2_nor2_1 _18850_ (.A(net2056),
    .B(net4295),
    .Y(_04141_));
 sg13g2_a21oi_1 _18851_ (.A1(net3818),
    .A2(net4292),
    .Y(_01835_),
    .B1(_04141_));
 sg13g2_nor3_2 _18852_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .C(_03743_),
    .Y(_04142_));
 sg13g2_nor2_1 _18853_ (.A(net872),
    .B(net4285),
    .Y(_04143_));
 sg13g2_a21oi_1 _18854_ (.A1(_07227_),
    .A2(net4285),
    .Y(_01836_),
    .B1(_04143_));
 sg13g2_nor2_1 _18855_ (.A(net986),
    .B(net4285),
    .Y(_04144_));
 sg13g2_a21oi_1 _18856_ (.A1(net3943),
    .A2(net4285),
    .Y(_01837_),
    .B1(_04144_));
 sg13g2_nor2_1 _18857_ (.A(net673),
    .B(net4285),
    .Y(_04145_));
 sg13g2_a21oi_1 _18858_ (.A1(net3941),
    .A2(net4285),
    .Y(_01838_),
    .B1(_04145_));
 sg13g2_nor2_1 _18859_ (.A(net732),
    .B(net4286),
    .Y(_04146_));
 sg13g2_a21oi_1 _18860_ (.A1(_07255_),
    .A2(net4286),
    .Y(_01839_),
    .B1(_04146_));
 sg13g2_nor2_1 _18861_ (.A(net512),
    .B(net4289),
    .Y(_04147_));
 sg13g2_a21oi_1 _18862_ (.A1(net3835),
    .A2(net4290),
    .Y(_01840_),
    .B1(_04147_));
 sg13g2_nor2_1 _18863_ (.A(net879),
    .B(net4289),
    .Y(_04148_));
 sg13g2_a21oi_1 _18864_ (.A1(net3937),
    .A2(net4289),
    .Y(_01841_),
    .B1(_04148_));
 sg13g2_nor2_1 _18865_ (.A(net1267),
    .B(net4289),
    .Y(_04149_));
 sg13g2_a21oi_1 _18866_ (.A1(_07282_),
    .A2(net4289),
    .Y(_01842_),
    .B1(_04149_));
 sg13g2_nor2_1 _18867_ (.A(net2016),
    .B(net4285),
    .Y(_04150_));
 sg13g2_a21oi_1 _18868_ (.A1(net3931),
    .A2(net4285),
    .Y(_01843_),
    .B1(_04150_));
 sg13g2_nor2_1 _18869_ (.A(net1594),
    .B(net4287),
    .Y(_04151_));
 sg13g2_a21oi_1 _18870_ (.A1(_07305_),
    .A2(net4282),
    .Y(_01844_),
    .B1(_04151_));
 sg13g2_nor2_1 _18871_ (.A(net548),
    .B(net4288),
    .Y(_04152_));
 sg13g2_a21oi_1 _18872_ (.A1(net3927),
    .A2(net4288),
    .Y(_01845_),
    .B1(_04152_));
 sg13g2_nor2_1 _18873_ (.A(net1171),
    .B(net4287),
    .Y(_04153_));
 sg13g2_a21oi_1 _18874_ (.A1(_07327_),
    .A2(net4287),
    .Y(_01846_),
    .B1(_04153_));
 sg13g2_nor2_1 _18875_ (.A(net1845),
    .B(net4286),
    .Y(_04154_));
 sg13g2_a21oi_1 _18876_ (.A1(_07339_),
    .A2(net4286),
    .Y(_01847_),
    .B1(_04154_));
 sg13g2_nor2_1 _18877_ (.A(net1335),
    .B(net4290),
    .Y(_04155_));
 sg13g2_a21oi_1 _18878_ (.A1(_07350_),
    .A2(net4289),
    .Y(_01848_),
    .B1(_04155_));
 sg13g2_nor2_1 _18879_ (.A(net715),
    .B(net4282),
    .Y(_04156_));
 sg13g2_a21oi_1 _18880_ (.A1(net3921),
    .A2(net4282),
    .Y(_01849_),
    .B1(_04156_));
 sg13g2_nor2_1 _18881_ (.A(net487),
    .B(net4289),
    .Y(_04157_));
 sg13g2_a21oi_1 _18882_ (.A1(net3918),
    .A2(net4289),
    .Y(_01850_),
    .B1(_04157_));
 sg13g2_nor2_1 _18883_ (.A(net555),
    .B(net4288),
    .Y(_04158_));
 sg13g2_a21oi_1 _18884_ (.A1(net3916),
    .A2(net4290),
    .Y(_01851_),
    .B1(_04158_));
 sg13g2_nor2_1 _18885_ (.A(net1027),
    .B(net4282),
    .Y(_04159_));
 sg13g2_a21oi_1 _18886_ (.A1(net3913),
    .A2(net4282),
    .Y(_01852_),
    .B1(_04159_));
 sg13g2_nor2_1 _18887_ (.A(net626),
    .B(net4283),
    .Y(_04160_));
 sg13g2_a21oi_1 _18888_ (.A1(net3831),
    .A2(net4283),
    .Y(_01853_),
    .B1(_04160_));
 sg13g2_nor2_1 _18889_ (.A(net723),
    .B(net4281),
    .Y(_04161_));
 sg13g2_a21oi_1 _18890_ (.A1(_07415_),
    .A2(net4281),
    .Y(_01854_),
    .B1(_04161_));
 sg13g2_nor2_1 _18891_ (.A(net768),
    .B(net4283),
    .Y(_04162_));
 sg13g2_a21oi_1 _18892_ (.A1(_07424_),
    .A2(net4283),
    .Y(_01855_),
    .B1(_04162_));
 sg13g2_nor2_1 _18893_ (.A(net1278),
    .B(net4281),
    .Y(_04163_));
 sg13g2_a21oi_1 _18894_ (.A1(net3904),
    .A2(net4281),
    .Y(_01856_),
    .B1(_04163_));
 sg13g2_nor2_1 _18895_ (.A(net561),
    .B(net4283),
    .Y(_04164_));
 sg13g2_a21oi_1 _18896_ (.A1(_07442_),
    .A2(net4283),
    .Y(_01857_),
    .B1(_04164_));
 sg13g2_nor2_1 _18897_ (.A(net769),
    .B(net4283),
    .Y(_04165_));
 sg13g2_a21oi_1 _18898_ (.A1(_07451_),
    .A2(net4283),
    .Y(_01858_),
    .B1(_04165_));
 sg13g2_nor2_1 _18899_ (.A(net739),
    .B(net4281),
    .Y(_04166_));
 sg13g2_a21oi_1 _18900_ (.A1(net3899),
    .A2(net4281),
    .Y(_01859_),
    .B1(_04166_));
 sg13g2_nor2_1 _18901_ (.A(net683),
    .B(net4288),
    .Y(_04167_));
 sg13g2_a21oi_1 _18902_ (.A1(_07468_),
    .A2(net4288),
    .Y(_01860_),
    .B1(_04167_));
 sg13g2_nor2_1 _18903_ (.A(net1268),
    .B(net4288),
    .Y(_04168_));
 sg13g2_a21oi_1 _18904_ (.A1(net3828),
    .A2(net4288),
    .Y(_01861_),
    .B1(_04168_));
 sg13g2_nor2_1 _18905_ (.A(net719),
    .B(net4287),
    .Y(_04169_));
 sg13g2_a21oi_1 _18906_ (.A1(net3825),
    .A2(net4287),
    .Y(_01862_),
    .B1(_04169_));
 sg13g2_nor2_1 _18907_ (.A(net1834),
    .B(net4282),
    .Y(_04170_));
 sg13g2_a21oi_1 _18908_ (.A1(net3895),
    .A2(net4282),
    .Y(_01863_),
    .B1(_04170_));
 sg13g2_nor2_1 _18909_ (.A(net654),
    .B(net4281),
    .Y(_04171_));
 sg13g2_a21oi_1 _18910_ (.A1(net3823),
    .A2(net4281),
    .Y(_01864_),
    .B1(_04171_));
 sg13g2_nor2_1 _18911_ (.A(net454),
    .B(net4284),
    .Y(_04172_));
 sg13g2_a21oi_1 _18912_ (.A1(net3820),
    .A2(net4284),
    .Y(_01865_),
    .B1(_04172_));
 sg13g2_nor2_1 _18913_ (.A(net2385),
    .B(net4286),
    .Y(_04173_));
 sg13g2_a21oi_1 _18914_ (.A1(net3893),
    .A2(net4286),
    .Y(_01866_),
    .B1(_04173_));
 sg13g2_nor2_1 _18915_ (.A(net1193),
    .B(net4288),
    .Y(_04174_));
 sg13g2_a21oi_1 _18916_ (.A1(_07524_),
    .A2(net4290),
    .Y(_01867_),
    .B1(_04174_));
 sg13g2_nand3_1 _18917_ (.B(_06695_),
    .C(_07606_),
    .A(net4248),
    .Y(_04175_));
 sg13g2_o21ai_1 _18918_ (.B1(net678),
    .Y(_04176_),
    .A1(_08476_),
    .A2(_04175_));
 sg13g2_or2_1 _18919_ (.X(_04177_),
    .B(_04175_),
    .A(_06738_));
 sg13g2_o21ai_1 _18920_ (.B1(_04176_),
    .Y(_01868_),
    .A1(_08474_),
    .A2(_04177_));
 sg13g2_o21ai_1 _18921_ (.B1(net643),
    .Y(_04178_),
    .A1(_08487_),
    .A2(_04175_));
 sg13g2_o21ai_1 _18922_ (.B1(_04178_),
    .Y(_01869_),
    .A1(_08485_),
    .A2(_04177_));
 sg13g2_nand2b_1 _18923_ (.Y(_04179_),
    .B(\soc_inst.cpu_core.id_rs1_data[24] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[24] ));
 sg13g2_nand2b_1 _18924_ (.Y(_04180_),
    .B(\soc_inst.cpu_core.id_rs1_data[25] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[25] ));
 sg13g2_nor2b_1 _18925_ (.A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .B_N(\soc_inst.cpu_core.id_rs2_data[25] ),
    .Y(_04181_));
 sg13g2_a21oi_1 _18926_ (.A1(_05666_),
    .A2(\soc_inst.cpu_core.id_rs2_data[26] ),
    .Y(_04182_),
    .B1(_04181_));
 sg13g2_and3_1 _18927_ (.X(_04183_),
    .A(_04179_),
    .B(_04180_),
    .C(_04182_));
 sg13g2_nor2b_1 _18928_ (.A(\soc_inst.cpu_core.id_rs1_data[31] ),
    .B_N(\soc_inst.cpu_core.id_rs2_data[31] ),
    .Y(_04184_));
 sg13g2_a21oi_1 _18929_ (.A1(_05663_),
    .A2(\soc_inst.cpu_core.id_rs2_data[30] ),
    .Y(_04185_),
    .B1(_04184_));
 sg13g2_a22oi_1 _18930_ (.Y(_04186_),
    .B1(\soc_inst.cpu_core.id_rs1_data[27] ),
    .B2(_05665_),
    .A2(_05664_),
    .A1(\soc_inst.cpu_core.id_rs1_data[28] ));
 sg13g2_nand2b_2 _18931_ (.Y(_04187_),
    .B(\soc_inst.cpu_core.id_rs1_data[31] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[31] ));
 sg13g2_nor2_1 _18932_ (.A(_05666_),
    .B(\soc_inst.cpu_core.id_rs2_data[26] ),
    .Y(_04188_));
 sg13g2_o21ai_1 _18933_ (.B1(_04187_),
    .Y(_04189_),
    .A1(_05666_),
    .A2(\soc_inst.cpu_core.id_rs2_data[26] ));
 sg13g2_nand2b_1 _18934_ (.Y(_04190_),
    .B(\soc_inst.cpu_core.id_rs2_data[27] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[27] ));
 sg13g2_o21ai_1 _18935_ (.B1(_04190_),
    .Y(_04191_),
    .A1(\soc_inst.cpu_core.id_rs1_data[24] ),
    .A2(_05667_));
 sg13g2_nand2b_1 _18936_ (.Y(_04192_),
    .B(\soc_inst.cpu_core.id_rs1_data[29] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[29] ));
 sg13g2_o21ai_1 _18937_ (.B1(_04192_),
    .Y(_04193_),
    .A1(_05663_),
    .A2(\soc_inst.cpu_core.id_rs2_data[30] ));
 sg13g2_nand2b_1 _18938_ (.Y(_04194_),
    .B(\soc_inst.cpu_core.id_rs2_data[29] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[29] ));
 sg13g2_o21ai_1 _18939_ (.B1(_04194_),
    .Y(_04195_),
    .A1(\soc_inst.cpu_core.id_rs1_data[28] ),
    .A2(_05664_));
 sg13g2_nor4_1 _18940_ (.A(_04189_),
    .B(_04191_),
    .C(_04193_),
    .D(_04195_),
    .Y(_04196_));
 sg13g2_nand4_1 _18941_ (.B(_04185_),
    .C(_04186_),
    .A(_04183_),
    .Y(_04197_),
    .D(_04196_));
 sg13g2_a22oi_1 _18942_ (.Y(_04198_),
    .B1(_05672_),
    .B2(\soc_inst.cpu_core.id_rs2_data[21] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[22] ),
    .A1(_05670_));
 sg13g2_a22oi_1 _18943_ (.Y(_04199_),
    .B1(_05676_),
    .B2(\soc_inst.cpu_core.id_rs2_data[18] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[19] ),
    .A1(_05674_));
 sg13g2_a22oi_1 _18944_ (.Y(_04200_),
    .B1(\soc_inst.cpu_core.id_rs1_data[22] ),
    .B2(_05671_),
    .A2(_05669_),
    .A1(\soc_inst.cpu_core.id_rs1_data[23] ));
 sg13g2_a22oi_1 _18945_ (.Y(_04201_),
    .B1(\soc_inst.cpu_core.id_rs1_data[19] ),
    .B2(_05675_),
    .A2(_05673_),
    .A1(\soc_inst.cpu_core.id_rs1_data[20] ));
 sg13g2_nand4_1 _18946_ (.B(_04199_),
    .C(_04200_),
    .A(_04198_),
    .Y(_04202_),
    .D(_04201_));
 sg13g2_nor2b_1 _18947_ (.A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .B_N(\soc_inst.cpu_core.id_rs2_data[17] ),
    .Y(_04203_));
 sg13g2_nor2b_1 _18948_ (.A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .B_N(\soc_inst.cpu_core.id_rs2_data[16] ),
    .Y(_04204_));
 sg13g2_nor2_1 _18949_ (.A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .B(_05673_),
    .Y(_04205_));
 sg13g2_nor2_1 _18950_ (.A(_05672_),
    .B(\soc_inst.cpu_core.id_rs2_data[21] ),
    .Y(_04206_));
 sg13g2_nor4_1 _18951_ (.A(_04203_),
    .B(_04204_),
    .C(_04205_),
    .D(_04206_),
    .Y(_04207_));
 sg13g2_nand2b_1 _18952_ (.Y(_04208_),
    .B(\soc_inst.cpu_core.id_rs1_data[16] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[16] ));
 sg13g2_nand2b_1 _18953_ (.Y(_04209_),
    .B(\soc_inst.cpu_core.id_rs1_data[17] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[17] ));
 sg13g2_nor2_1 _18954_ (.A(_05676_),
    .B(\soc_inst.cpu_core.id_rs2_data[18] ),
    .Y(_04210_));
 sg13g2_a21oi_1 _18955_ (.A1(_05668_),
    .A2(\soc_inst.cpu_core.id_rs2_data[23] ),
    .Y(_04211_),
    .B1(_04210_));
 sg13g2_nand4_1 _18956_ (.B(_04208_),
    .C(_04209_),
    .A(_04207_),
    .Y(_04212_),
    .D(_04211_));
 sg13g2_nor3_2 _18957_ (.A(_04197_),
    .B(_04202_),
    .C(_04212_),
    .Y(_04213_));
 sg13g2_a22oi_1 _18958_ (.Y(_04214_),
    .B1(_05660_),
    .B2(\soc_inst.cpu_core.id_rs2_data[14] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[15] ),
    .A1(_05658_));
 sg13g2_nand2b_1 _18959_ (.Y(_04215_),
    .B(\soc_inst.cpu_core.id_rs2_data[12] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[12] ));
 sg13g2_nand2b_1 _18960_ (.Y(_04216_),
    .B(\soc_inst.cpu_core.id_rs2_data[13] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[13] ));
 sg13g2_nand3_1 _18961_ (.B(_04215_),
    .C(_04216_),
    .A(_04214_),
    .Y(_04217_));
 sg13g2_nor2b_1 _18962_ (.A(\soc_inst.cpu_core.id_rs2_data[11] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[11] ),
    .Y(_04218_));
 sg13g2_a21o_1 _18963_ (.A2(_05661_),
    .A1(\soc_inst.cpu_core.id_rs1_data[10] ),
    .B1(_04218_),
    .X(_04219_));
 sg13g2_nand2b_1 _18964_ (.Y(_04220_),
    .B(\soc_inst.cpu_core.id_rs2_data[11] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[11] ));
 sg13g2_o21ai_1 _18965_ (.B1(_04220_),
    .Y(_04221_),
    .A1(\soc_inst.cpu_core.id_rs1_data[10] ),
    .A2(_05661_));
 sg13g2_nor2_1 _18966_ (.A(_04219_),
    .B(_04221_),
    .Y(_04222_));
 sg13g2_nor2b_1 _18967_ (.A(\soc_inst.cpu_core.id_rs2_data[9] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[9] ),
    .Y(_04223_));
 sg13g2_a21o_1 _18968_ (.A2(_05662_),
    .A1(\soc_inst.cpu_core.id_rs1_data[8] ),
    .B1(_04223_),
    .X(_04224_));
 sg13g2_nand2b_1 _18969_ (.Y(_04225_),
    .B(\soc_inst.cpu_core.id_rs1_data[13] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[13] ));
 sg13g2_o21ai_1 _18970_ (.B1(_04225_),
    .Y(_04226_),
    .A1(_05660_),
    .A2(\soc_inst.cpu_core.id_rs2_data[14] ));
 sg13g2_nand2b_1 _18971_ (.Y(_04227_),
    .B(\soc_inst.cpu_core.id_rs2_data[9] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[9] ));
 sg13g2_o21ai_1 _18972_ (.B1(_04227_),
    .Y(_04228_),
    .A1(\soc_inst.cpu_core.id_rs1_data[8] ),
    .A2(_05662_));
 sg13g2_nor3_1 _18973_ (.A(_04224_),
    .B(_04226_),
    .C(_04228_),
    .Y(_04229_));
 sg13g2_a22oi_1 _18974_ (.Y(_04230_),
    .B1(_05653_),
    .B2(\soc_inst.cpu_core.id_rs2_data[6] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[7] ),
    .A1(_05652_));
 sg13g2_nand2_1 _18975_ (.Y(_04231_),
    .A(_04229_),
    .B(_04230_));
 sg13g2_nor2_1 _18976_ (.A(_05653_),
    .B(\soc_inst.cpu_core.id_rs2_data[6] ),
    .Y(_04232_));
 sg13g2_a21oi_1 _18977_ (.A1(\soc_inst.cpu_core.id_rs1_data[5] ),
    .A2(_05655_),
    .Y(_04233_),
    .B1(_04232_));
 sg13g2_a22oi_1 _18978_ (.Y(_04234_),
    .B1(_05656_),
    .B2(\soc_inst.cpu_core.id_rs2_data[4] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[5] ),
    .A1(_05654_));
 sg13g2_nand2b_1 _18979_ (.Y(_04235_),
    .B(\soc_inst.cpu_core.id_rs2_data[2] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[2] ));
 sg13g2_nor2b_1 _18980_ (.A(\soc_inst.cpu_core.id_rs2_data[2] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[2] ),
    .Y(_04236_));
 sg13g2_nand2b_1 _18981_ (.Y(_04237_),
    .B(\soc_inst.cpu_core.id_rs1_data[2] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[2] ));
 sg13g2_nand2b_1 _18982_ (.Y(_04238_),
    .B(\soc_inst.cpu_core.id_rs2_data[3] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[3] ));
 sg13g2_nand3_1 _18983_ (.B(_04237_),
    .C(_04238_),
    .A(_04235_),
    .Y(_04239_));
 sg13g2_nand2b_1 _18984_ (.Y(_04240_),
    .B(\soc_inst.cpu_core.id_rs2_data[1] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[1] ));
 sg13g2_nand2b_1 _18985_ (.Y(_04241_),
    .B(\soc_inst.cpu_core.id_rs2_data[0] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[0] ));
 sg13g2_nor2b_1 _18986_ (.A(\soc_inst.cpu_core.id_rs2_data[1] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[1] ),
    .Y(_04242_));
 sg13g2_a21oi_1 _18987_ (.A1(_04240_),
    .A2(_04241_),
    .Y(_04243_),
    .B1(_04242_));
 sg13g2_nor2_1 _18988_ (.A(_05656_),
    .B(\soc_inst.cpu_core.id_rs2_data[4] ),
    .Y(_04244_));
 sg13g2_nor2b_1 _18989_ (.A(\soc_inst.cpu_core.id_rs2_data[3] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[3] ),
    .Y(_04245_));
 sg13g2_a221oi_1 _18990_ (.B2(_04238_),
    .C1(_04245_),
    .B1(_04236_),
    .A1(\soc_inst.cpu_core.id_rs1_data[4] ),
    .Y(_04246_),
    .A2(_05657_));
 sg13g2_o21ai_1 _18991_ (.B1(_04246_),
    .Y(_04247_),
    .A1(_04239_),
    .A2(_04243_));
 sg13g2_a221oi_1 _18992_ (.B2(_04247_),
    .C1(_04232_),
    .B1(_04234_),
    .A1(\soc_inst.cpu_core.id_rs1_data[5] ),
    .Y(_04248_),
    .A2(_05655_));
 sg13g2_nor2_1 _18993_ (.A(_05652_),
    .B(\soc_inst.cpu_core.id_rs2_data[7] ),
    .Y(_04249_));
 sg13g2_a22oi_1 _18994_ (.Y(_04250_),
    .B1(_04229_),
    .B2(_04249_),
    .A2(_04227_),
    .A1(_04224_));
 sg13g2_o21ai_1 _18995_ (.B1(_04250_),
    .Y(_04251_),
    .A1(_04231_),
    .A2(_04248_));
 sg13g2_nor2b_1 _18996_ (.A(\soc_inst.cpu_core.id_rs2_data[12] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[12] ),
    .Y(_04252_));
 sg13g2_a221oi_1 _18997_ (.B2(_04251_),
    .C1(_04252_),
    .B1(_04222_),
    .A1(_04219_),
    .Y(_04253_),
    .A2(_04220_));
 sg13g2_a22oi_1 _18998_ (.Y(_04254_),
    .B1(_04214_),
    .B2(_04226_),
    .A2(_05659_),
    .A1(\soc_inst.cpu_core.id_rs1_data[15] ));
 sg13g2_o21ai_1 _18999_ (.B1(_04254_),
    .Y(_04255_),
    .A1(_04217_),
    .A2(_04253_));
 sg13g2_a221oi_1 _19000_ (.B2(_04180_),
    .C1(_04181_),
    .B1(_04179_),
    .A1(_05666_),
    .Y(_04256_),
    .A2(\soc_inst.cpu_core.id_rs2_data[26] ));
 sg13g2_o21ai_1 _19001_ (.B1(_04190_),
    .Y(_04257_),
    .A1(_04188_),
    .A2(_04256_));
 sg13g2_a21oi_1 _19002_ (.A1(_04186_),
    .A2(_04257_),
    .Y(_04258_),
    .B1(_04195_));
 sg13g2_o21ai_1 _19003_ (.B1(_04185_),
    .Y(_04259_),
    .A1(_04193_),
    .A2(_04258_));
 sg13g2_nand2_1 _19004_ (.Y(_04260_),
    .A(_04187_),
    .B(_04259_));
 sg13g2_a21oi_1 _19005_ (.A1(_04208_),
    .A2(_04209_),
    .Y(_04261_),
    .B1(_04203_));
 sg13g2_o21ai_1 _19006_ (.B1(_04199_),
    .Y(_04262_),
    .A1(_04210_),
    .A2(_04261_));
 sg13g2_a21oi_1 _19007_ (.A1(_04201_),
    .A2(_04262_),
    .Y(_04263_),
    .B1(_04205_));
 sg13g2_o21ai_1 _19008_ (.B1(_04198_),
    .Y(_04264_),
    .A1(_04206_),
    .A2(_04263_));
 sg13g2_a221oi_1 _19009_ (.B2(_04264_),
    .C1(_04197_),
    .B1(_04200_),
    .A1(_05668_),
    .Y(_04265_),
    .A2(\soc_inst.cpu_core.id_rs2_data[23] ));
 sg13g2_or2_1 _19010_ (.X(_04266_),
    .B(_04265_),
    .A(_04260_));
 sg13g2_a21o_1 _19011_ (.A2(_04255_),
    .A1(_04213_),
    .B1(_04266_),
    .X(_04267_));
 sg13g2_nand2_1 _19012_ (.Y(_04268_),
    .A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[0] ));
 sg13g2_nor2b_1 _19013_ (.A(\soc_inst.cpu_core.id_funct3[0] ),
    .B_N(\soc_inst.cpu_core.id_funct3[2] ),
    .Y(_04269_));
 sg13g2_o21ai_1 _19014_ (.B1(\soc_inst.cpu_core.id_funct3[1] ),
    .Y(_04270_),
    .A1(_04267_),
    .A2(_04269_));
 sg13g2_a21oi_1 _19015_ (.A1(_04267_),
    .A2(_04268_),
    .Y(_04271_),
    .B1(_04270_));
 sg13g2_a21oi_1 _19016_ (.A1(_04187_),
    .A2(_04267_),
    .Y(_04272_),
    .B1(_04184_));
 sg13g2_nor2b_1 _19017_ (.A(\soc_inst.cpu_core.id_funct3[1] ),
    .B_N(_04269_),
    .Y(_04273_));
 sg13g2_nor3_1 _19018_ (.A(\soc_inst.cpu_core.id_funct3[1] ),
    .B(_04268_),
    .C(_04272_),
    .Y(_04274_));
 sg13g2_or2_1 _19019_ (.X(_04275_),
    .B(_04274_),
    .A(_04271_));
 sg13g2_a21o_2 _19020_ (.A2(_04273_),
    .A1(_04272_),
    .B1(_04275_),
    .X(_04276_));
 sg13g2_nand2_1 _19021_ (.Y(_04277_),
    .A(\soc_inst.cpu_core.id_funct3[0] ),
    .B(_09223_));
 sg13g2_nand2_1 _19022_ (.Y(_04278_),
    .A(\soc_inst.cpu_core.id_imm[0] ),
    .B(\soc_inst.cpu_core.id_pc[0] ));
 sg13g2_xor2_1 _19023_ (.B(\soc_inst.cpu_core.id_pc[0] ),
    .A(\soc_inst.cpu_core.id_imm[0] ),
    .X(_04279_));
 sg13g2_nand2_1 _19024_ (.Y(_04280_),
    .A(_04276_),
    .B(_04279_));
 sg13g2_o21ai_1 _19025_ (.B1(_04280_),
    .Y(_04281_),
    .A1(_05677_),
    .A2(_04276_));
 sg13g2_nor4_1 _19026_ (.A(_04217_),
    .B(_04219_),
    .C(_04221_),
    .D(_04239_),
    .Y(_04282_));
 sg13g2_nand4_1 _19027_ (.B(_04234_),
    .C(_04240_),
    .A(_04233_),
    .Y(_04283_),
    .D(_04241_));
 sg13g2_a221oi_1 _19028_ (.B2(_05659_),
    .C1(_04242_),
    .B1(\soc_inst.cpu_core.id_rs1_data[15] ),
    .A1(\soc_inst.cpu_core.id_rs1_data[0] ),
    .Y(_04284_),
    .A2(_05651_));
 sg13g2_nor2_1 _19029_ (.A(_04249_),
    .B(_04252_),
    .Y(_04285_));
 sg13g2_nand3_1 _19030_ (.B(_04284_),
    .C(_04285_),
    .A(_04230_),
    .Y(_04286_));
 sg13g2_nor4_1 _19031_ (.A(_04244_),
    .B(_04245_),
    .C(_04283_),
    .D(_04286_),
    .Y(_04287_));
 sg13g2_nand4_1 _19032_ (.B(_04229_),
    .C(_04282_),
    .A(_04213_),
    .Y(_04288_),
    .D(_04287_));
 sg13g2_nand2b_1 _19033_ (.Y(_04289_),
    .B(_04288_),
    .A_N(_04277_));
 sg13g2_and4_1 _19034_ (.A(\soc_inst.cpu_core.id_funct3[0] ),
    .B(_09223_),
    .C(_04279_),
    .D(_04288_),
    .X(_04290_));
 sg13g2_nor2_1 _19035_ (.A(_04277_),
    .B(_04288_),
    .Y(_04291_));
 sg13g2_inv_1 _19036_ (.Y(_04292_),
    .A(_04291_));
 sg13g2_a221oi_1 _19037_ (.B2(\soc_inst.cpu_core.id_pc[0] ),
    .C1(_04290_),
    .B1(_04291_),
    .A1(_04277_),
    .Y(_04293_),
    .A2(_04281_));
 sg13g2_or2_1 _19038_ (.X(_04294_),
    .B(_04293_),
    .A(_09224_));
 sg13g2_nand2_2 _19039_ (.Y(_04295_),
    .A(_09224_),
    .B(_04288_));
 sg13g2_inv_1 _19040_ (.Y(_04296_),
    .A(_04295_));
 sg13g2_and3_2 _19041_ (.X(_04297_),
    .A(\soc_inst.cpu_core.id_instr[5] ),
    .B(net4878),
    .C(_09215_));
 sg13g2_nand3_1 _19042_ (.B(\soc_inst.cpu_core.id_instr[6] ),
    .C(_09215_),
    .A(\soc_inst.cpu_core.id_instr[5] ),
    .Y(_04298_));
 sg13g2_or4_1 _19043_ (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[0] ),
    .C(\soc_inst.cpu_core.id_funct3[1] ),
    .D(_04288_),
    .X(_04299_));
 sg13g2_inv_1 _19044_ (.Y(_04300_),
    .A(_04299_));
 sg13g2_a221oi_1 _19045_ (.B2(_04279_),
    .C1(net4107),
    .B1(_04300_),
    .A1(\soc_inst.cpu_core.id_pc[0] ),
    .Y(_04301_),
    .A2(_04296_));
 sg13g2_nand2_1 _19046_ (.Y(_04302_),
    .A(net4119),
    .B(_04279_));
 sg13g2_a221oi_1 _19047_ (.B2(net4107),
    .C1(net4920),
    .B1(_04302_),
    .A1(_04294_),
    .Y(_04303_),
    .A2(_04301_));
 sg13g2_a21o_1 _19048_ (.A2(net4924),
    .A1(net1805),
    .B1(_04303_),
    .X(_01870_));
 sg13g2_nand2_1 _19049_ (.Y(_04304_),
    .A(\soc_inst.cpu_core.id_pc[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xnor2_1 _19050_ (.Y(_04305_),
    .A(\soc_inst.cpu_core.id_pc[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xnor2_1 _19051_ (.Y(_04306_),
    .A(_04278_),
    .B(_04305_));
 sg13g2_inv_1 _19052_ (.Y(_04307_),
    .A(_04306_));
 sg13g2_nand2_1 _19053_ (.Y(_04308_),
    .A(_05678_),
    .B(\soc_inst.cpu_core.id_is_compressed ));
 sg13g2_xor2_1 _19054_ (.B(\soc_inst.cpu_core.id_is_compressed ),
    .A(\soc_inst.cpu_core.id_pc[1] ),
    .X(_04309_));
 sg13g2_mux2_1 _19055_ (.A0(_04309_),
    .A1(_04307_),
    .S(_04276_),
    .X(_04310_));
 sg13g2_nor2_1 _19056_ (.A(_04289_),
    .B(_04306_),
    .Y(_04311_));
 sg13g2_a221oi_1 _19057_ (.B2(_04277_),
    .C1(_04311_),
    .B1(_04310_),
    .A1(_04291_),
    .Y(_04312_),
    .A2(_04309_));
 sg13g2_nor2_1 _19058_ (.A(_09224_),
    .B(_04312_),
    .Y(_04313_));
 sg13g2_a21oi_1 _19059_ (.A1(_04296_),
    .A2(_04309_),
    .Y(_04314_),
    .B1(net4107));
 sg13g2_o21ai_1 _19060_ (.B1(_04314_),
    .Y(_04315_),
    .A1(_04299_),
    .A2(_04306_));
 sg13g2_nor2_1 _19061_ (.A(_04313_),
    .B(_04315_),
    .Y(_04316_));
 sg13g2_nand2_1 _19062_ (.Y(_04317_),
    .A(\soc_inst.cpu_core.id_rs1_data[0] ),
    .B(\soc_inst.cpu_core.id_imm[0] ));
 sg13g2_nand2_1 _19063_ (.Y(_04318_),
    .A(\soc_inst.cpu_core.id_rs1_data[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xnor2_1 _19064_ (.Y(_04319_),
    .A(\soc_inst.cpu_core.id_rs1_data[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xor2_1 _19065_ (.B(_04319_),
    .A(_04317_),
    .X(_04320_));
 sg13g2_a221oi_1 _19066_ (.B2(net4217),
    .C1(net4110),
    .B1(_04320_),
    .A1(net4119),
    .Y(_04321_),
    .A2(_04307_));
 sg13g2_nor3_1 _19067_ (.A(net4935),
    .B(_04316_),
    .C(_04321_),
    .Y(_04322_));
 sg13g2_a21o_1 _19068_ (.A2(net2441),
    .A1(net4939),
    .B1(_04322_),
    .X(_01871_));
 sg13g2_nand2b_1 _19069_ (.Y(_04323_),
    .B(_04289_),
    .A_N(_04276_));
 sg13g2_o21ai_1 _19070_ (.B1(_04295_),
    .Y(_04324_),
    .A1(_09224_),
    .A2(_04323_));
 sg13g2_nand2_2 _19071_ (.Y(_04325_),
    .A(net4109),
    .B(_04324_));
 sg13g2_inv_1 _19072_ (.Y(_04326_),
    .A(_04325_));
 sg13g2_nand2_1 _19073_ (.Y(_04327_),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .B(_04308_));
 sg13g2_xnor2_1 _19074_ (.Y(_04328_),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .B(_04308_));
 sg13g2_and2_1 _19075_ (.A(\soc_inst.cpu_core.id_pc[2] ),
    .B(\soc_inst.cpu_core.id_imm[2] ),
    .X(_04329_));
 sg13g2_xor2_1 _19076_ (.B(\soc_inst.cpu_core.id_imm[2] ),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .X(_04330_));
 sg13g2_o21ai_1 _19077_ (.B1(_04304_),
    .Y(_04331_),
    .A1(_04278_),
    .A2(_04305_));
 sg13g2_xnor2_1 _19078_ (.Y(_04332_),
    .A(_04330_),
    .B(_04331_));
 sg13g2_nor2_2 _19079_ (.A(net4107),
    .B(_04324_),
    .Y(_04333_));
 sg13g2_or2_1 _19080_ (.X(_04334_),
    .B(_04324_),
    .A(net4107));
 sg13g2_and2_1 _19081_ (.A(\soc_inst.cpu_core.id_rs1_data[2] ),
    .B(\soc_inst.cpu_core.id_imm[2] ),
    .X(_04335_));
 sg13g2_xor2_1 _19082_ (.B(\soc_inst.cpu_core.id_imm[2] ),
    .A(\soc_inst.cpu_core.id_rs1_data[2] ),
    .X(_04336_));
 sg13g2_o21ai_1 _19083_ (.B1(_04318_),
    .Y(_04337_),
    .A1(_04317_),
    .A2(_04319_));
 sg13g2_nand2_1 _19084_ (.Y(_04338_),
    .A(_04336_),
    .B(_04337_));
 sg13g2_o21ai_1 _19085_ (.B1(net4217),
    .Y(_04339_),
    .A1(_04336_),
    .A2(_04337_));
 sg13g2_inv_1 _19086_ (.Y(_04340_),
    .A(_04339_));
 sg13g2_a21oi_1 _19087_ (.A1(_04338_),
    .A2(_04340_),
    .Y(_04341_),
    .B1(net4110));
 sg13g2_o21ai_1 _19088_ (.B1(_04341_),
    .Y(_04342_),
    .A1(_09232_),
    .A2(_04332_));
 sg13g2_a221oi_1 _19089_ (.B2(_04333_),
    .C1(net4935),
    .B1(_04332_),
    .A1(net3715),
    .Y(_04343_),
    .A2(_04328_));
 sg13g2_a22oi_1 _19090_ (.Y(_04344_),
    .B1(_04342_),
    .B2(_04343_),
    .A2(net1888),
    .A1(net4939));
 sg13g2_inv_1 _19091_ (.Y(_01872_),
    .A(net1889));
 sg13g2_xnor2_1 _19092_ (.Y(_04345_),
    .A(net2987),
    .B(_04327_));
 sg13g2_nand2_1 _19093_ (.Y(_04346_),
    .A(\soc_inst.cpu_core.id_pc[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_xnor2_1 _19094_ (.Y(_04347_),
    .A(\soc_inst.cpu_core.id_pc[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_a21oi_1 _19095_ (.A1(_04330_),
    .A2(_04331_),
    .Y(_04348_),
    .B1(_04329_));
 sg13g2_xor2_1 _19096_ (.B(_04348_),
    .A(_04347_),
    .X(_04349_));
 sg13g2_nor2_1 _19097_ (.A(_04334_),
    .B(_04349_),
    .Y(_04350_));
 sg13g2_nand2_1 _19098_ (.Y(_04351_),
    .A(\soc_inst.cpu_core.id_rs1_data[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_xnor2_1 _19099_ (.Y(_04352_),
    .A(\soc_inst.cpu_core.id_rs1_data[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_a21oi_1 _19100_ (.A1(_04336_),
    .A2(_04337_),
    .Y(_04353_),
    .B1(_04335_));
 sg13g2_nor2_1 _19101_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sg13g2_a21o_1 _19102_ (.A2(_04353_),
    .A1(_04352_),
    .B1(net4120),
    .X(_04355_));
 sg13g2_a21oi_1 _19103_ (.A1(net4119),
    .A2(_04349_),
    .Y(_04356_),
    .B1(net4110));
 sg13g2_o21ai_1 _19104_ (.B1(_04356_),
    .Y(_04357_),
    .A1(_04354_),
    .A2(_04355_));
 sg13g2_o21ai_1 _19105_ (.B1(_04357_),
    .Y(_04358_),
    .A1(_04325_),
    .A2(_04345_));
 sg13g2_nor3_1 _19106_ (.A(net4939),
    .B(_04350_),
    .C(_04358_),
    .Y(_04359_));
 sg13g2_a21o_1 _19107_ (.A2(net2384),
    .A1(net4938),
    .B1(_04359_),
    .X(_01873_));
 sg13g2_nand4_1 _19108_ (.B(\soc_inst.cpu_core.id_pc[3] ),
    .C(\soc_inst.cpu_core.id_pc[4] ),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .Y(_04360_),
    .D(_04308_));
 sg13g2_o21ai_1 _19109_ (.B1(_05681_),
    .Y(_04361_),
    .A1(_05680_),
    .A2(_04327_));
 sg13g2_a21oi_1 _19110_ (.A1(_04360_),
    .A2(_04361_),
    .Y(_04362_),
    .B1(_04325_));
 sg13g2_and2_1 _19111_ (.A(\soc_inst.cpu_core.id_pc[4] ),
    .B(\soc_inst.cpu_core.id_imm[4] ),
    .X(_04363_));
 sg13g2_xor2_1 _19112_ (.B(\soc_inst.cpu_core.id_imm[4] ),
    .A(\soc_inst.cpu_core.id_pc[4] ),
    .X(_04364_));
 sg13g2_o21ai_1 _19113_ (.B1(_04346_),
    .Y(_04365_),
    .A1(_04347_),
    .A2(_04348_));
 sg13g2_xor2_1 _19114_ (.B(_04365_),
    .A(_04364_),
    .X(_04366_));
 sg13g2_and2_1 _19115_ (.A(\soc_inst.cpu_core.id_rs1_data[4] ),
    .B(\soc_inst.cpu_core.id_imm[4] ),
    .X(_04367_));
 sg13g2_xor2_1 _19116_ (.B(\soc_inst.cpu_core.id_imm[4] ),
    .A(\soc_inst.cpu_core.id_rs1_data[4] ),
    .X(_04368_));
 sg13g2_o21ai_1 _19117_ (.B1(_04351_),
    .Y(_04369_),
    .A1(_04352_),
    .A2(_04353_));
 sg13g2_nand2_1 _19118_ (.Y(_04370_),
    .A(_04368_),
    .B(_04369_));
 sg13g2_nor2_1 _19119_ (.A(_04368_),
    .B(_04369_),
    .Y(_04371_));
 sg13g2_nor2_1 _19120_ (.A(net4120),
    .B(_04371_),
    .Y(_04372_));
 sg13g2_a221oi_1 _19121_ (.B2(_04372_),
    .C1(net4110),
    .B1(_04370_),
    .A1(net4119),
    .Y(_04373_),
    .A2(_04366_));
 sg13g2_nor3_1 _19122_ (.A(net4940),
    .B(_04362_),
    .C(_04373_),
    .Y(_04374_));
 sg13g2_o21ai_1 _19123_ (.B1(_04374_),
    .Y(_04375_),
    .A1(_04334_),
    .A2(_04366_));
 sg13g2_o21ai_1 _19124_ (.B1(_04375_),
    .Y(_01874_),
    .A1(net4752),
    .A2(_05709_));
 sg13g2_nor2_1 _19125_ (.A(_05682_),
    .B(_04360_),
    .Y(_04376_));
 sg13g2_xnor2_1 _19126_ (.Y(_04377_),
    .A(_05682_),
    .B(_04360_));
 sg13g2_a21oi_1 _19127_ (.A1(_04364_),
    .A2(_04365_),
    .Y(_04378_),
    .B1(_04363_));
 sg13g2_nor2_1 _19128_ (.A(\soc_inst.cpu_core.id_pc[5] ),
    .B(\soc_inst.cpu_core.id_imm[5] ),
    .Y(_04379_));
 sg13g2_xor2_1 _19129_ (.B(\soc_inst.cpu_core.id_imm[5] ),
    .A(\soc_inst.cpu_core.id_pc[5] ),
    .X(_04380_));
 sg13g2_xnor2_1 _19130_ (.Y(_04381_),
    .A(_04378_),
    .B(_04380_));
 sg13g2_a21oi_1 _19131_ (.A1(_04368_),
    .A2(_04369_),
    .Y(_04382_),
    .B1(_04367_));
 sg13g2_nor2_1 _19132_ (.A(\soc_inst.cpu_core.id_rs1_data[5] ),
    .B(\soc_inst.cpu_core.id_imm[5] ),
    .Y(_04383_));
 sg13g2_xnor2_1 _19133_ (.Y(_04384_),
    .A(\soc_inst.cpu_core.id_rs1_data[5] ),
    .B(\soc_inst.cpu_core.id_imm[5] ));
 sg13g2_a21oi_1 _19134_ (.A1(_04382_),
    .A2(_04384_),
    .Y(_04385_),
    .B1(net4120));
 sg13g2_o21ai_1 _19135_ (.B1(_04385_),
    .Y(_04386_),
    .A1(_04382_),
    .A2(_04384_));
 sg13g2_a21oi_1 _19136_ (.A1(net4119),
    .A2(_04381_),
    .Y(_04387_),
    .B1(net4109));
 sg13g2_a221oi_1 _19137_ (.B2(_04387_),
    .C1(net4940),
    .B1(_04386_),
    .A1(net3715),
    .Y(_04388_),
    .A2(_04377_));
 sg13g2_o21ai_1 _19138_ (.B1(_04388_),
    .Y(_04389_),
    .A1(_04334_),
    .A2(_04381_));
 sg13g2_o21ai_1 _19139_ (.B1(_04389_),
    .Y(_01875_),
    .A1(net4752),
    .A2(_05710_));
 sg13g2_nor3_2 _19140_ (.A(_05682_),
    .B(_05683_),
    .C(_04360_),
    .Y(_04390_));
 sg13g2_xnor2_1 _19141_ (.Y(_04391_),
    .A(\soc_inst.cpu_core.id_pc[6] ),
    .B(_04376_));
 sg13g2_xnor2_1 _19142_ (.Y(_04392_),
    .A(\soc_inst.cpu_core.id_pc[6] ),
    .B(\soc_inst.cpu_core.id_imm[6] ));
 sg13g2_a221oi_1 _19143_ (.B2(_04365_),
    .C1(_04363_),
    .B1(_04364_),
    .A1(\soc_inst.cpu_core.id_pc[5] ),
    .Y(_04393_),
    .A2(\soc_inst.cpu_core.id_imm[5] ));
 sg13g2_nor3_1 _19144_ (.A(_04379_),
    .B(_04392_),
    .C(_04393_),
    .Y(_04394_));
 sg13g2_o21ai_1 _19145_ (.B1(_04392_),
    .Y(_04395_),
    .A1(_04379_),
    .A2(_04393_));
 sg13g2_nand2b_1 _19146_ (.Y(_04396_),
    .B(_04395_),
    .A_N(_04394_));
 sg13g2_or2_1 _19147_ (.X(_04397_),
    .B(_04396_),
    .A(_09232_));
 sg13g2_and2_1 _19148_ (.A(\soc_inst.cpu_core.id_rs1_data[6] ),
    .B(\soc_inst.cpu_core.id_imm[6] ),
    .X(_04398_));
 sg13g2_xnor2_1 _19149_ (.Y(_04399_),
    .A(\soc_inst.cpu_core.id_rs1_data[6] ),
    .B(\soc_inst.cpu_core.id_imm[6] ));
 sg13g2_a221oi_1 _19150_ (.B2(_04369_),
    .C1(_04367_),
    .B1(_04368_),
    .A1(\soc_inst.cpu_core.id_rs1_data[5] ),
    .Y(_04400_),
    .A2(\soc_inst.cpu_core.id_imm[5] ));
 sg13g2_nor3_1 _19151_ (.A(_04383_),
    .B(_04399_),
    .C(_04400_),
    .Y(_04401_));
 sg13g2_o21ai_1 _19152_ (.B1(_04399_),
    .Y(_04402_),
    .A1(_04383_),
    .A2(_04400_));
 sg13g2_nand3b_1 _19153_ (.B(_04402_),
    .C(net4217),
    .Y(_04403_),
    .A_N(_04401_));
 sg13g2_nand3_1 _19154_ (.B(_04397_),
    .C(_04403_),
    .A(net4108),
    .Y(_04404_));
 sg13g2_a221oi_1 _19155_ (.B2(_04333_),
    .C1(net4937),
    .B1(_04396_),
    .A1(net3715),
    .Y(_04405_),
    .A2(_04391_));
 sg13g2_a22oi_1 _19156_ (.Y(_04406_),
    .B1(_04404_),
    .B2(_04405_),
    .A2(net2728),
    .A1(net4936));
 sg13g2_inv_1 _19157_ (.Y(_01876_),
    .A(net2729));
 sg13g2_nor2_2 _19158_ (.A(net4119),
    .B(_04333_),
    .Y(_04407_));
 sg13g2_nand2_2 _19159_ (.Y(_04408_),
    .A(_09232_),
    .B(_04334_));
 sg13g2_a21oi_1 _19160_ (.A1(\soc_inst.cpu_core.id_pc[6] ),
    .A2(\soc_inst.cpu_core.id_imm[6] ),
    .Y(_04409_),
    .B1(_04394_));
 sg13g2_nor2_1 _19161_ (.A(\soc_inst.cpu_core.id_pc[7] ),
    .B(\soc_inst.cpu_core.id_imm[7] ),
    .Y(_04410_));
 sg13g2_xor2_1 _19162_ (.B(net2036),
    .A(\soc_inst.cpu_core.id_pc[7] ),
    .X(_04411_));
 sg13g2_xnor2_1 _19163_ (.Y(_04412_),
    .A(_04409_),
    .B(_04411_));
 sg13g2_xnor2_1 _19164_ (.Y(_04413_),
    .A(\soc_inst.cpu_core.id_pc[7] ),
    .B(_04390_));
 sg13g2_nand2_1 _19165_ (.Y(_04414_),
    .A(\soc_inst.cpu_core.id_rs1_data[7] ),
    .B(\soc_inst.cpu_core.id_imm[7] ));
 sg13g2_xor2_1 _19166_ (.B(\soc_inst.cpu_core.id_imm[7] ),
    .A(\soc_inst.cpu_core.id_rs1_data[7] ),
    .X(_04415_));
 sg13g2_o21ai_1 _19167_ (.B1(_04415_),
    .Y(_04416_),
    .A1(_04398_),
    .A2(_04401_));
 sg13g2_nor3_1 _19168_ (.A(_04398_),
    .B(_04401_),
    .C(_04415_),
    .Y(_04417_));
 sg13g2_nor2_1 _19169_ (.A(_09230_),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_a21oi_1 _19170_ (.A1(_04416_),
    .A2(_04418_),
    .Y(_04419_),
    .B1(net4937));
 sg13g2_o21ai_1 _19171_ (.B1(_04419_),
    .Y(_04420_),
    .A1(_04325_),
    .A2(_04413_));
 sg13g2_a21oi_1 _19172_ (.A1(_04408_),
    .A2(_04412_),
    .Y(_04421_),
    .B1(_04420_));
 sg13g2_a21oi_1 _19173_ (.A1(net4972),
    .A2(_05711_),
    .Y(_01877_),
    .B1(_04421_));
 sg13g2_nand2_1 _19174_ (.Y(_04422_),
    .A(net4938),
    .B(net1461));
 sg13g2_nand2_1 _19175_ (.Y(_04423_),
    .A(\soc_inst.cpu_core.id_pc[8] ),
    .B(\soc_inst.cpu_core.id_imm[8] ));
 sg13g2_xor2_1 _19176_ (.B(\soc_inst.cpu_core.id_imm[8] ),
    .A(\soc_inst.cpu_core.id_pc[8] ),
    .X(_04424_));
 sg13g2_a221oi_1 _19177_ (.B2(\soc_inst.cpu_core.id_imm[7] ),
    .C1(_04394_),
    .B1(\soc_inst.cpu_core.id_pc[7] ),
    .A1(\soc_inst.cpu_core.id_pc[6] ),
    .Y(_04425_),
    .A2(\soc_inst.cpu_core.id_imm[6] ));
 sg13g2_nor2_1 _19178_ (.A(_04410_),
    .B(_04425_),
    .Y(_04426_));
 sg13g2_nand2_1 _19179_ (.Y(_04427_),
    .A(_04424_),
    .B(_04426_));
 sg13g2_xor2_1 _19180_ (.B(_04426_),
    .A(_04424_),
    .X(_04428_));
 sg13g2_nor2_1 _19181_ (.A(_04334_),
    .B(_04428_),
    .Y(_04429_));
 sg13g2_and3_2 _19182_ (.X(_04430_),
    .A(\soc_inst.cpu_core.id_pc[7] ),
    .B(\soc_inst.cpu_core.id_pc[8] ),
    .C(_04390_));
 sg13g2_a21oi_1 _19183_ (.A1(\soc_inst.cpu_core.id_pc[7] ),
    .A2(_04390_),
    .Y(_04431_),
    .B1(\soc_inst.cpu_core.id_pc[8] ));
 sg13g2_nor2_1 _19184_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 sg13g2_and2_1 _19185_ (.A(_04414_),
    .B(_04416_),
    .X(_04433_));
 sg13g2_nand2_1 _19186_ (.Y(_04434_),
    .A(\soc_inst.cpu_core.id_rs1_data[8] ),
    .B(\soc_inst.cpu_core.id_imm[8] ));
 sg13g2_xnor2_1 _19187_ (.Y(_04435_),
    .A(\soc_inst.cpu_core.id_rs1_data[8] ),
    .B(\soc_inst.cpu_core.id_imm[8] ));
 sg13g2_or2_1 _19188_ (.X(_04436_),
    .B(_04435_),
    .A(_04433_));
 sg13g2_nand2_1 _19189_ (.Y(_04437_),
    .A(net4217),
    .B(_04436_));
 sg13g2_a21oi_1 _19190_ (.A1(_04433_),
    .A2(_04435_),
    .Y(_04438_),
    .B1(_04437_));
 sg13g2_a21oi_1 _19191_ (.A1(_09231_),
    .A2(_04428_),
    .Y(_04439_),
    .B1(_04438_));
 sg13g2_a21oi_1 _19192_ (.A1(net4108),
    .A2(_04439_),
    .Y(_04440_),
    .B1(net4935));
 sg13g2_o21ai_1 _19193_ (.B1(_04440_),
    .Y(_04441_),
    .A1(_04325_),
    .A2(_04432_));
 sg13g2_o21ai_1 _19194_ (.B1(_04422_),
    .Y(_01878_),
    .A1(_04429_),
    .A2(_04441_));
 sg13g2_xnor2_1 _19195_ (.Y(_04442_),
    .A(\soc_inst.cpu_core.id_pc[9] ),
    .B(_04430_));
 sg13g2_nor2_1 _19196_ (.A(\soc_inst.cpu_core.id_pc[9] ),
    .B(\soc_inst.cpu_core.id_imm[9] ),
    .Y(_04443_));
 sg13g2_nand2_1 _19197_ (.Y(_04444_),
    .A(\soc_inst.cpu_core.id_pc[9] ),
    .B(\soc_inst.cpu_core.id_imm[9] ));
 sg13g2_nor2b_1 _19198_ (.A(_04443_),
    .B_N(_04444_),
    .Y(_04445_));
 sg13g2_nand2_1 _19199_ (.Y(_04446_),
    .A(_04423_),
    .B(_04427_));
 sg13g2_xnor2_1 _19200_ (.Y(_04447_),
    .A(_04445_),
    .B(_04446_));
 sg13g2_nand2_1 _19201_ (.Y(_04448_),
    .A(\soc_inst.cpu_core.id_rs1_data[9] ),
    .B(\soc_inst.cpu_core.id_imm[9] ));
 sg13g2_xnor2_1 _19202_ (.Y(_04449_),
    .A(\soc_inst.cpu_core.id_rs1_data[9] ),
    .B(\soc_inst.cpu_core.id_imm[9] ));
 sg13g2_and2_1 _19203_ (.A(_04434_),
    .B(_04436_),
    .X(_04450_));
 sg13g2_nor2_1 _19204_ (.A(_04449_),
    .B(_04450_),
    .Y(_04451_));
 sg13g2_o21ai_1 _19205_ (.B1(net4217),
    .Y(_04452_),
    .A1(_04449_),
    .A2(_04450_));
 sg13g2_a21oi_1 _19206_ (.A1(_04449_),
    .A2(_04450_),
    .Y(_04453_),
    .B1(_04452_));
 sg13g2_o21ai_1 _19207_ (.B1(net4107),
    .Y(_04454_),
    .A1(_09232_),
    .A2(_04447_));
 sg13g2_o21ai_1 _19208_ (.B1(net4752),
    .Y(_04455_),
    .A1(_04453_),
    .A2(_04454_));
 sg13g2_a221oi_1 _19209_ (.B2(_04333_),
    .C1(_04455_),
    .B1(_04447_),
    .A1(net3715),
    .Y(_04456_),
    .A2(_04442_));
 sg13g2_a21o_1 _19210_ (.A2(net2208),
    .A1(net4976),
    .B1(_04456_),
    .X(_01879_));
 sg13g2_xor2_1 _19211_ (.B(\soc_inst.cpu_core.id_imm[10] ),
    .A(\soc_inst.cpu_core.id_pc[10] ),
    .X(_04457_));
 sg13g2_o21ai_1 _19212_ (.B1(_04444_),
    .Y(_04458_),
    .A1(_04423_),
    .A2(_04443_));
 sg13g2_nand2_1 _19213_ (.Y(_04459_),
    .A(_04424_),
    .B(_04445_));
 sg13g2_nor3_1 _19214_ (.A(_04410_),
    .B(_04425_),
    .C(_04459_),
    .Y(_04460_));
 sg13g2_o21ai_1 _19215_ (.B1(_04457_),
    .Y(_04461_),
    .A1(_04458_),
    .A2(_04460_));
 sg13g2_or3_1 _19216_ (.A(_04457_),
    .B(_04458_),
    .C(_04460_),
    .X(_04462_));
 sg13g2_and2_1 _19217_ (.A(_04461_),
    .B(_04462_),
    .X(_04463_));
 sg13g2_inv_1 _19218_ (.Y(_04464_),
    .A(_04463_));
 sg13g2_nand2_1 _19219_ (.Y(_04465_),
    .A(\soc_inst.cpu_core.id_rs1_data[10] ),
    .B(\soc_inst.cpu_core.id_imm[10] ));
 sg13g2_xnor2_1 _19220_ (.Y(_04466_),
    .A(\soc_inst.cpu_core.id_rs1_data[10] ),
    .B(\soc_inst.cpu_core.id_imm[10] ));
 sg13g2_a21oi_1 _19221_ (.A1(\soc_inst.cpu_core.id_rs1_data[9] ),
    .A2(\soc_inst.cpu_core.id_imm[9] ),
    .Y(_04467_),
    .B1(_04451_));
 sg13g2_or2_1 _19222_ (.X(_04468_),
    .B(_04467_),
    .A(_04466_));
 sg13g2_a21oi_1 _19223_ (.A1(_04466_),
    .A2(_04467_),
    .Y(_04469_),
    .B1(net4120));
 sg13g2_a221oi_1 _19224_ (.B2(_04469_),
    .C1(net4109),
    .B1(_04468_),
    .A1(_09231_),
    .Y(_04470_),
    .A2(_04463_));
 sg13g2_nand3_1 _19225_ (.B(\soc_inst.cpu_core.id_pc[10] ),
    .C(_04430_),
    .A(\soc_inst.cpu_core.id_pc[9] ),
    .Y(_04471_));
 sg13g2_a21o_1 _19226_ (.A2(_04430_),
    .A1(\soc_inst.cpu_core.id_pc[9] ),
    .B1(\soc_inst.cpu_core.id_pc[10] ),
    .X(_04472_));
 sg13g2_nand2_1 _19227_ (.Y(_04473_),
    .A(_04471_),
    .B(_04472_));
 sg13g2_nand2b_1 _19228_ (.Y(_04474_),
    .B(_04473_),
    .A_N(_04323_));
 sg13g2_a21oi_1 _19229_ (.A1(_04323_),
    .A2(_04464_),
    .Y(_04475_),
    .B1(_09224_));
 sg13g2_o21ai_1 _19230_ (.B1(net4109),
    .Y(_04476_),
    .A1(_04295_),
    .A2(_04473_));
 sg13g2_a221oi_1 _19231_ (.B2(_04475_),
    .C1(_04476_),
    .B1(_04474_),
    .A1(_04300_),
    .Y(_04477_),
    .A2(_04463_));
 sg13g2_nor3_1 _19232_ (.A(net4935),
    .B(_04470_),
    .C(_04477_),
    .Y(_04478_));
 sg13g2_a21o_1 _19233_ (.A2(net2263),
    .A1(net4965),
    .B1(_04478_),
    .X(_01880_));
 sg13g2_nor2_1 _19234_ (.A(\soc_inst.cpu_core.id_rs1_data[11] ),
    .B(\soc_inst.cpu_core.id_imm[11] ),
    .Y(_04479_));
 sg13g2_xnor2_1 _19235_ (.Y(_04480_),
    .A(\soc_inst.cpu_core.id_rs1_data[11] ),
    .B(\soc_inst.cpu_core.id_imm[11] ));
 sg13g2_nand3_1 _19236_ (.B(_04468_),
    .C(_04480_),
    .A(_04465_),
    .Y(_04481_));
 sg13g2_a21oi_1 _19237_ (.A1(_04465_),
    .A2(_04468_),
    .Y(_04482_),
    .B1(_04480_));
 sg13g2_nor2_1 _19238_ (.A(net4120),
    .B(_04482_),
    .Y(_04483_));
 sg13g2_xor2_1 _19239_ (.B(\soc_inst.cpu_core.id_imm[11] ),
    .A(\soc_inst.cpu_core.id_pc[11] ),
    .X(_04484_));
 sg13g2_o21ai_1 _19240_ (.B1(_04461_),
    .Y(_04485_),
    .A1(_05687_),
    .A2(_05688_));
 sg13g2_xnor2_1 _19241_ (.Y(_04486_),
    .A(_04484_),
    .B(_04485_));
 sg13g2_o21ai_1 _19242_ (.B1(net4108),
    .Y(_04487_),
    .A1(_09232_),
    .A2(_04486_));
 sg13g2_a21oi_1 _19243_ (.A1(_04481_),
    .A2(_04483_),
    .Y(_04488_),
    .B1(_04487_));
 sg13g2_nor2_1 _19244_ (.A(_05689_),
    .B(_04471_),
    .Y(_04489_));
 sg13g2_xnor2_1 _19245_ (.Y(_04490_),
    .A(\soc_inst.cpu_core.id_pc[11] ),
    .B(_04471_));
 sg13g2_a21oi_1 _19246_ (.A1(_04333_),
    .A2(_04486_),
    .Y(_04491_),
    .B1(net4920));
 sg13g2_o21ai_1 _19247_ (.B1(_04491_),
    .Y(_04492_),
    .A1(_04325_),
    .A2(_04490_));
 sg13g2_nand2_1 _19248_ (.Y(_04493_),
    .A(net4924),
    .B(net1825));
 sg13g2_o21ai_1 _19249_ (.B1(_04493_),
    .Y(_01881_),
    .A1(_04488_),
    .A2(_04492_));
 sg13g2_nand2_1 _19250_ (.Y(_04494_),
    .A(net4924),
    .B(net1322));
 sg13g2_and2_1 _19251_ (.A(\soc_inst.cpu_core.id_pc[12] ),
    .B(\soc_inst.cpu_core.id_imm[12] ),
    .X(_04495_));
 sg13g2_xor2_1 _19252_ (.B(\soc_inst.cpu_core.id_imm[12] ),
    .A(\soc_inst.cpu_core.id_pc[12] ),
    .X(_04496_));
 sg13g2_a22oi_1 _19253_ (.Y(_04497_),
    .B1(\soc_inst.cpu_core.id_pc[11] ),
    .B2(\soc_inst.cpu_core.id_imm[11] ),
    .A2(\soc_inst.cpu_core.id_imm[10] ),
    .A1(\soc_inst.cpu_core.id_pc[10] ));
 sg13g2_a22oi_1 _19254_ (.Y(_04498_),
    .B1(_04461_),
    .B2(_04497_),
    .A2(_05690_),
    .A1(_05689_));
 sg13g2_xor2_1 _19255_ (.B(_04498_),
    .A(_04496_),
    .X(_04499_));
 sg13g2_nor2_1 _19256_ (.A(_04466_),
    .B(_04480_),
    .Y(_04500_));
 sg13g2_or4_1 _19257_ (.A(_04435_),
    .B(_04449_),
    .C(_04466_),
    .D(_04480_),
    .X(_04501_));
 sg13g2_a21oi_1 _19258_ (.A1(_04414_),
    .A2(_04416_),
    .Y(_04502_),
    .B1(_04501_));
 sg13g2_o21ai_1 _19259_ (.B1(_04448_),
    .Y(_04503_),
    .A1(_04434_),
    .A2(_04449_));
 sg13g2_a22oi_1 _19260_ (.Y(_04504_),
    .B1(_04500_),
    .B2(_04503_),
    .A2(\soc_inst.cpu_core.id_imm[11] ),
    .A1(\soc_inst.cpu_core.id_rs1_data[11] ));
 sg13g2_o21ai_1 _19261_ (.B1(_04504_),
    .Y(_04505_),
    .A1(_04465_),
    .A2(_04479_));
 sg13g2_nand2_1 _19262_ (.Y(_04506_),
    .A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .B(\soc_inst.cpu_core.id_imm[12] ));
 sg13g2_xnor2_1 _19263_ (.Y(_04507_),
    .A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .B(\soc_inst.cpu_core.id_imm[12] ));
 sg13g2_inv_1 _19264_ (.Y(_04508_),
    .A(_04507_));
 sg13g2_o21ai_1 _19265_ (.B1(_04508_),
    .Y(_04509_),
    .A1(_04502_),
    .A2(_04505_));
 sg13g2_nor3_1 _19266_ (.A(_04502_),
    .B(_04505_),
    .C(_04508_),
    .Y(_04510_));
 sg13g2_nor2_1 _19267_ (.A(net4120),
    .B(_04510_),
    .Y(_04511_));
 sg13g2_a22oi_1 _19268_ (.Y(_04512_),
    .B1(_04509_),
    .B2(_04511_),
    .A2(_04499_),
    .A1(net4119));
 sg13g2_nor2_1 _19269_ (.A(_04334_),
    .B(_04499_),
    .Y(_04513_));
 sg13g2_xnor2_1 _19270_ (.Y(_04514_),
    .A(_05691_),
    .B(_04489_));
 sg13g2_a21oi_1 _19271_ (.A1(net4107),
    .A2(_04512_),
    .Y(_04515_),
    .B1(net4920));
 sg13g2_o21ai_1 _19272_ (.B1(_04515_),
    .Y(_04516_),
    .A1(_04325_),
    .A2(_04514_));
 sg13g2_o21ai_1 _19273_ (.B1(_04494_),
    .Y(_01882_),
    .A1(_04513_),
    .A2(_04516_));
 sg13g2_nor2_1 _19274_ (.A(\soc_inst.cpu_core.id_pc[13] ),
    .B(\soc_inst.cpu_core.id_imm[13] ),
    .Y(_04517_));
 sg13g2_xor2_1 _19275_ (.B(\soc_inst.cpu_core.id_imm[13] ),
    .A(\soc_inst.cpu_core.id_pc[13] ),
    .X(_04518_));
 sg13g2_a21oi_1 _19276_ (.A1(_04496_),
    .A2(_04498_),
    .Y(_04519_),
    .B1(_04495_));
 sg13g2_xnor2_1 _19277_ (.Y(_04520_),
    .A(_04518_),
    .B(_04519_));
 sg13g2_nor2_1 _19278_ (.A(\soc_inst.cpu_core.id_rs1_data[13] ),
    .B(\soc_inst.cpu_core.id_imm[13] ),
    .Y(_04521_));
 sg13g2_nand2_1 _19279_ (.Y(_04522_),
    .A(\soc_inst.cpu_core.id_rs1_data[13] ),
    .B(\soc_inst.cpu_core.id_imm[13] ));
 sg13g2_nand2b_1 _19280_ (.Y(_04523_),
    .B(_04522_),
    .A_N(_04521_));
 sg13g2_nand3_1 _19281_ (.B(_04509_),
    .C(_04523_),
    .A(_04506_),
    .Y(_04524_));
 sg13g2_a21oi_1 _19282_ (.A1(_04506_),
    .A2(_04509_),
    .Y(_04525_),
    .B1(_04523_));
 sg13g2_nor2_1 _19283_ (.A(net4120),
    .B(_04525_),
    .Y(_04526_));
 sg13g2_a221oi_1 _19284_ (.B2(_04526_),
    .C1(net4109),
    .B1(_04524_),
    .A1(net4119),
    .Y(_04527_),
    .A2(_04520_));
 sg13g2_nor2_1 _19285_ (.A(_04334_),
    .B(_04520_),
    .Y(_04528_));
 sg13g2_nand3_1 _19286_ (.B(\soc_inst.cpu_core.id_pc[13] ),
    .C(_04489_),
    .A(\soc_inst.cpu_core.id_pc[12] ),
    .Y(_04529_));
 sg13g2_a21o_1 _19287_ (.A2(_04489_),
    .A1(\soc_inst.cpu_core.id_pc[12] ),
    .B1(\soc_inst.cpu_core.id_pc[13] ),
    .X(_04530_));
 sg13g2_a21oi_1 _19288_ (.A1(_04529_),
    .A2(_04530_),
    .Y(_04531_),
    .B1(_04325_));
 sg13g2_nor4_1 _19289_ (.A(net4924),
    .B(_04527_),
    .C(_04528_),
    .D(_04531_),
    .Y(_04532_));
 sg13g2_a21o_1 _19290_ (.A2(net2352),
    .A1(net4961),
    .B1(_04532_),
    .X(_01883_));
 sg13g2_nand2_1 _19291_ (.Y(_04533_),
    .A(net4920),
    .B(net1107));
 sg13g2_nor2_1 _19292_ (.A(\soc_inst.cpu_core.id_pc[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ),
    .Y(_04534_));
 sg13g2_nand2_1 _19293_ (.Y(_04535_),
    .A(\soc_inst.cpu_core.id_pc[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ));
 sg13g2_nor2b_1 _19294_ (.A(_04534_),
    .B_N(_04535_),
    .Y(_04536_));
 sg13g2_a21oi_1 _19295_ (.A1(\soc_inst.cpu_core.id_pc[13] ),
    .A2(\soc_inst.cpu_core.id_imm[13] ),
    .Y(_04537_),
    .B1(_04495_));
 sg13g2_nor2_1 _19296_ (.A(_04517_),
    .B(_04519_),
    .Y(_04538_));
 sg13g2_a21oi_1 _19297_ (.A1(\soc_inst.cpu_core.id_pc[13] ),
    .A2(\soc_inst.cpu_core.id_imm[13] ),
    .Y(_04539_),
    .B1(_04538_));
 sg13g2_xor2_1 _19298_ (.B(_04539_),
    .A(_04536_),
    .X(_04540_));
 sg13g2_nor2_2 _19299_ (.A(_05693_),
    .B(_04529_),
    .Y(_04541_));
 sg13g2_xnor2_1 _19300_ (.Y(_04542_),
    .A(_05693_),
    .B(_04529_));
 sg13g2_mux2_1 _19301_ (.A0(_04542_),
    .A1(_04540_),
    .S(_04276_),
    .X(_04543_));
 sg13g2_nor2_1 _19302_ (.A(_09223_),
    .B(_04543_),
    .Y(_04544_));
 sg13g2_a21oi_1 _19303_ (.A1(_04289_),
    .A2(_04299_),
    .Y(_04545_),
    .B1(_04540_));
 sg13g2_a21oi_1 _19304_ (.A1(_04292_),
    .A2(_04295_),
    .Y(_04546_),
    .B1(_04542_));
 sg13g2_nor4_1 _19305_ (.A(net4107),
    .B(_04544_),
    .C(_04545_),
    .D(_04546_),
    .Y(_04547_));
 sg13g2_nand2_1 _19306_ (.Y(_04548_),
    .A(\soc_inst.cpu_core.id_rs1_data[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ));
 sg13g2_xor2_1 _19307_ (.B(\soc_inst.cpu_core.id_imm[14] ),
    .A(\soc_inst.cpu_core.id_rs1_data[14] ),
    .X(_04549_));
 sg13g2_inv_1 _19308_ (.Y(_04550_),
    .A(_04549_));
 sg13g2_a21o_1 _19309_ (.A2(\soc_inst.cpu_core.id_imm[13] ),
    .A1(\soc_inst.cpu_core.id_rs1_data[13] ),
    .B1(_04525_),
    .X(_04551_));
 sg13g2_and2_1 _19310_ (.A(_04549_),
    .B(_04551_),
    .X(_04552_));
 sg13g2_nor2_1 _19311_ (.A(net4120),
    .B(_04552_),
    .Y(_04553_));
 sg13g2_o21ai_1 _19312_ (.B1(_04553_),
    .Y(_04554_),
    .A1(_04549_),
    .A2(_04551_));
 sg13g2_o21ai_1 _19313_ (.B1(_04554_),
    .Y(_04555_),
    .A1(_09232_),
    .A2(_04540_));
 sg13g2_o21ai_1 _19314_ (.B1(net4751),
    .Y(_04556_),
    .A1(net4109),
    .A2(_04555_));
 sg13g2_o21ai_1 _19315_ (.B1(_04533_),
    .Y(_01884_),
    .A1(_04547_),
    .A2(_04556_));
 sg13g2_nor2_1 _19316_ (.A(\soc_inst.cpu_core.id_pc[15] ),
    .B(\soc_inst.cpu_core.id_imm[15] ),
    .Y(_04557_));
 sg13g2_xor2_1 _19317_ (.B(\soc_inst.cpu_core.id_imm[15] ),
    .A(\soc_inst.cpu_core.id_pc[15] ),
    .X(_04558_));
 sg13g2_o21ai_1 _19318_ (.B1(_04535_),
    .Y(_04559_),
    .A1(_04534_),
    .A2(_04539_));
 sg13g2_xor2_1 _19319_ (.B(_04559_),
    .A(_04558_),
    .X(_04560_));
 sg13g2_xnor2_1 _19320_ (.Y(_04561_),
    .A(\soc_inst.cpu_core.id_rs1_data[15] ),
    .B(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_a21oi_1 _19321_ (.A1(\soc_inst.cpu_core.id_rs1_data[14] ),
    .A2(\soc_inst.cpu_core.id_imm[14] ),
    .Y(_04562_),
    .B1(_04552_));
 sg13g2_o21ai_1 _19322_ (.B1(net4216),
    .Y(_04563_),
    .A1(_04561_),
    .A2(_04562_));
 sg13g2_a21oi_1 _19323_ (.A1(_04561_),
    .A2(_04562_),
    .Y(_04564_),
    .B1(_04563_));
 sg13g2_xnor2_1 _19324_ (.Y(_04565_),
    .A(_05694_),
    .B(_04541_));
 sg13g2_nand2_1 _19325_ (.Y(_04566_),
    .A(net4965),
    .B(net508));
 sg13g2_a221oi_1 _19326_ (.B2(net3715),
    .C1(_04564_),
    .B1(_04565_),
    .A1(net3713),
    .Y(_04567_),
    .A2(_04560_));
 sg13g2_o21ai_1 _19327_ (.B1(_04566_),
    .Y(_01885_),
    .A1(net4965),
    .A2(_04567_));
 sg13g2_and2_1 _19328_ (.A(_04536_),
    .B(_04558_),
    .X(_04568_));
 sg13g2_nand3_1 _19329_ (.B(_04518_),
    .C(_04568_),
    .A(_04496_),
    .Y(_04569_));
 sg13g2_a221oi_1 _19330_ (.B2(_04497_),
    .C1(_04569_),
    .B1(_04461_),
    .A1(_05689_),
    .Y(_04570_),
    .A2(_05690_));
 sg13g2_nor2_1 _19331_ (.A(_04517_),
    .B(_04537_),
    .Y(_04571_));
 sg13g2_nand2_1 _19332_ (.Y(_04572_),
    .A(_04568_),
    .B(_04571_));
 sg13g2_a22oi_1 _19333_ (.Y(_04573_),
    .B1(\soc_inst.cpu_core.id_pc[15] ),
    .B2(\soc_inst.cpu_core.id_imm[15] ),
    .A2(\soc_inst.cpu_core.id_imm[14] ),
    .A1(\soc_inst.cpu_core.id_pc[14] ));
 sg13g2_o21ai_1 _19334_ (.B1(_04572_),
    .Y(_04574_),
    .A1(_04557_),
    .A2(_04573_));
 sg13g2_or2_1 _19335_ (.X(_04575_),
    .B(_04574_),
    .A(_04570_));
 sg13g2_nand2_1 _19336_ (.Y(_04576_),
    .A(\soc_inst.cpu_core.id_pc[16] ),
    .B(\soc_inst.cpu_core.id_imm[16] ));
 sg13g2_xor2_1 _19337_ (.B(\soc_inst.cpu_core.id_imm[16] ),
    .A(\soc_inst.cpu_core.id_pc[16] ),
    .X(_04577_));
 sg13g2_nand2_1 _19338_ (.Y(_04578_),
    .A(_04575_),
    .B(_04577_));
 sg13g2_or2_1 _19339_ (.X(_04579_),
    .B(_04577_),
    .A(_04575_));
 sg13g2_nand3_1 _19340_ (.B(_04578_),
    .C(_04579_),
    .A(net3712),
    .Y(_04580_));
 sg13g2_nor2_1 _19341_ (.A(_04550_),
    .B(_04561_),
    .Y(_04581_));
 sg13g2_nand2b_1 _19342_ (.Y(_04582_),
    .B(_04581_),
    .A_N(_04523_));
 sg13g2_o21ai_1 _19343_ (.B1(_04522_),
    .Y(_04583_),
    .A1(_04506_),
    .A2(_04521_));
 sg13g2_a21oi_1 _19344_ (.A1(_05658_),
    .A2(_05695_),
    .Y(_04584_),
    .B1(_04548_));
 sg13g2_a221oi_1 _19345_ (.B2(_04583_),
    .C1(_04584_),
    .B1(_04581_),
    .A1(\soc_inst.cpu_core.id_rs1_data[15] ),
    .Y(_04585_),
    .A2(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_o21ai_1 _19346_ (.B1(_04585_),
    .Y(_04586_),
    .A1(_04509_),
    .A2(_04582_));
 sg13g2_nand2_1 _19347_ (.Y(_04587_),
    .A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .B(\soc_inst.cpu_core.id_imm[16] ));
 sg13g2_xnor2_1 _19348_ (.Y(_04588_),
    .A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .B(\soc_inst.cpu_core.id_imm[16] ));
 sg13g2_nand2b_2 _19349_ (.Y(_04589_),
    .B(_04586_),
    .A_N(_04588_));
 sg13g2_nor2b_1 _19350_ (.A(_04586_),
    .B_N(_04588_),
    .Y(_04590_));
 sg13g2_nor2_1 _19351_ (.A(net4121),
    .B(_04590_),
    .Y(_04591_));
 sg13g2_nand3_1 _19352_ (.B(\soc_inst.cpu_core.id_pc[16] ),
    .C(_04541_),
    .A(\soc_inst.cpu_core.id_pc[15] ),
    .Y(_04592_));
 sg13g2_a21o_1 _19353_ (.A2(_04541_),
    .A1(\soc_inst.cpu_core.id_pc[15] ),
    .B1(\soc_inst.cpu_core.id_pc[16] ),
    .X(_04593_));
 sg13g2_and2_1 _19354_ (.A(_04592_),
    .B(_04593_),
    .X(_04594_));
 sg13g2_a221oi_1 _19355_ (.B2(net3714),
    .C1(net4912),
    .B1(_04594_),
    .A1(_04589_),
    .Y(_04595_),
    .A2(_04591_));
 sg13g2_a22oi_1 _19356_ (.Y(_01886_),
    .B1(_04580_),
    .B2(_04595_),
    .A2(_05712_),
    .A1(net4917));
 sg13g2_nor2_1 _19357_ (.A(net4751),
    .B(net1301),
    .Y(_04596_));
 sg13g2_nor2_1 _19358_ (.A(\soc_inst.cpu_core.id_pc[17] ),
    .B(\soc_inst.cpu_core.id_imm[17] ),
    .Y(_04597_));
 sg13g2_xor2_1 _19359_ (.B(\soc_inst.cpu_core.id_imm[17] ),
    .A(\soc_inst.cpu_core.id_pc[17] ),
    .X(_04598_));
 sg13g2_and2_1 _19360_ (.A(_04576_),
    .B(_04578_),
    .X(_04599_));
 sg13g2_xnor2_1 _19361_ (.Y(_04600_),
    .A(_04598_),
    .B(_04599_));
 sg13g2_nand2_1 _19362_ (.Y(_04601_),
    .A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .B(\soc_inst.cpu_core.id_imm[17] ));
 sg13g2_xnor2_1 _19363_ (.Y(_04602_),
    .A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .B(\soc_inst.cpu_core.id_imm[17] ));
 sg13g2_nand3_1 _19364_ (.B(_04589_),
    .C(_04602_),
    .A(_04587_),
    .Y(_04603_));
 sg13g2_or2_1 _19365_ (.X(_04604_),
    .B(_04602_),
    .A(_04589_));
 sg13g2_or2_1 _19366_ (.X(_04605_),
    .B(_04602_),
    .A(_04587_));
 sg13g2_and4_1 _19367_ (.A(net4216),
    .B(_04603_),
    .C(_04604_),
    .D(_04605_),
    .X(_04606_));
 sg13g2_nor2_1 _19368_ (.A(_05697_),
    .B(_04592_),
    .Y(_04607_));
 sg13g2_xnor2_1 _19369_ (.Y(_04608_),
    .A(\soc_inst.cpu_core.id_pc[17] ),
    .B(_04592_));
 sg13g2_a221oi_1 _19370_ (.B2(net3714),
    .C1(_04606_),
    .B1(_04608_),
    .A1(net3712),
    .Y(_04609_),
    .A2(_04600_));
 sg13g2_a21oi_1 _19371_ (.A1(net4751),
    .A2(_04609_),
    .Y(_01887_),
    .B1(_04596_));
 sg13g2_nand2_1 _19372_ (.Y(_04610_),
    .A(\soc_inst.cpu_core.id_pc[18] ),
    .B(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_xor2_1 _19373_ (.B(\soc_inst.cpu_core.id_imm[18] ),
    .A(\soc_inst.cpu_core.id_pc[18] ),
    .X(_04611_));
 sg13g2_a22oi_1 _19374_ (.Y(_04612_),
    .B1(\soc_inst.cpu_core.id_pc[17] ),
    .B2(\soc_inst.cpu_core.id_imm[17] ),
    .A2(\soc_inst.cpu_core.id_imm[16] ),
    .A1(\soc_inst.cpu_core.id_pc[16] ));
 sg13g2_a21oi_1 _19375_ (.A1(_04578_),
    .A2(_04612_),
    .Y(_04613_),
    .B1(_04597_));
 sg13g2_xor2_1 _19376_ (.B(_04613_),
    .A(_04611_),
    .X(_04614_));
 sg13g2_nand2_1 _19377_ (.Y(_04615_),
    .A(\soc_inst.cpu_core.id_rs1_data[18] ),
    .B(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_xnor2_1 _19378_ (.Y(_04616_),
    .A(\soc_inst.cpu_core.id_rs1_data[18] ),
    .B(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_nand2_1 _19379_ (.Y(_04617_),
    .A(_04601_),
    .B(_04605_));
 sg13g2_nand2b_1 _19380_ (.Y(_04618_),
    .B(_04604_),
    .A_N(_04617_));
 sg13g2_nand2b_1 _19381_ (.Y(_04619_),
    .B(_04618_),
    .A_N(_04616_));
 sg13g2_nand2b_1 _19382_ (.Y(_04620_),
    .B(_04616_),
    .A_N(_04618_));
 sg13g2_nand3_1 _19383_ (.B(_04619_),
    .C(_04620_),
    .A(net4216),
    .Y(_04621_));
 sg13g2_nor3_1 _19384_ (.A(_05697_),
    .B(_05698_),
    .C(_04592_),
    .Y(_04622_));
 sg13g2_xnor2_1 _19385_ (.Y(_04623_),
    .A(_05698_),
    .B(_04607_));
 sg13g2_a221oi_1 _19386_ (.B2(net3714),
    .C1(net4917),
    .B1(_04623_),
    .A1(net3712),
    .Y(_04624_),
    .A2(_04614_));
 sg13g2_a22oi_1 _19387_ (.Y(_01888_),
    .B1(_04621_),
    .B2(_04624_),
    .A2(_05713_),
    .A1(net4917));
 sg13g2_nor2_1 _19388_ (.A(\soc_inst.cpu_core.id_pc[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ),
    .Y(_04625_));
 sg13g2_nand2_1 _19389_ (.Y(_04626_),
    .A(\soc_inst.cpu_core.id_pc[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ));
 sg13g2_nor2b_2 _19390_ (.A(_04625_),
    .B_N(_04626_),
    .Y(_04627_));
 sg13g2_o21ai_1 _19391_ (.B1(_04613_),
    .Y(_04628_),
    .A1(\soc_inst.cpu_core.id_pc[18] ),
    .A2(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_nand2_1 _19392_ (.Y(_04629_),
    .A(_04610_),
    .B(_04628_));
 sg13g2_xor2_1 _19393_ (.B(_04629_),
    .A(_04627_),
    .X(_04630_));
 sg13g2_nor2_1 _19394_ (.A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ),
    .Y(_04631_));
 sg13g2_nand2_1 _19395_ (.Y(_04632_),
    .A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ));
 sg13g2_nand2b_1 _19396_ (.Y(_04633_),
    .B(_04632_),
    .A_N(_04631_));
 sg13g2_nand3_1 _19397_ (.B(_04619_),
    .C(_04633_),
    .A(_04615_),
    .Y(_04634_));
 sg13g2_a21o_1 _19398_ (.A2(_04619_),
    .A1(_04615_),
    .B1(_04633_),
    .X(_04635_));
 sg13g2_nand3_1 _19399_ (.B(_04634_),
    .C(_04635_),
    .A(net4216),
    .Y(_04636_));
 sg13g2_xnor2_1 _19400_ (.Y(_04637_),
    .A(_05699_),
    .B(_04622_));
 sg13g2_a221oi_1 _19401_ (.B2(net3714),
    .C1(net4910),
    .B1(_04637_),
    .A1(net3712),
    .Y(_04638_),
    .A2(_04630_));
 sg13g2_a22oi_1 _19402_ (.Y(_01889_),
    .B1(_04636_),
    .B2(_04638_),
    .A2(_05714_),
    .A1(net4912));
 sg13g2_nand2_1 _19403_ (.Y(_04639_),
    .A(_04611_),
    .B(_04627_));
 sg13g2_and4_1 _19404_ (.A(_04577_),
    .B(_04598_),
    .C(_04611_),
    .D(_04627_),
    .X(_04640_));
 sg13g2_o21ai_1 _19405_ (.B1(_04640_),
    .Y(_04641_),
    .A1(_04570_),
    .A2(_04574_));
 sg13g2_a21oi_1 _19406_ (.A1(_04610_),
    .A2(_04626_),
    .Y(_04642_),
    .B1(_04625_));
 sg13g2_nor3_1 _19407_ (.A(_04597_),
    .B(_04612_),
    .C(_04639_),
    .Y(_04643_));
 sg13g2_nor2_1 _19408_ (.A(_04642_),
    .B(_04643_),
    .Y(_04644_));
 sg13g2_nand2_1 _19409_ (.Y(_04645_),
    .A(_04641_),
    .B(_04644_));
 sg13g2_xnor2_1 _19410_ (.Y(_04646_),
    .A(\soc_inst.cpu_core.id_pc[20] ),
    .B(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_xnor2_1 _19411_ (.Y(_04647_),
    .A(_04645_),
    .B(_04646_));
 sg13g2_nand2_1 _19412_ (.Y(_04648_),
    .A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .B(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_xnor2_1 _19413_ (.Y(_04649_),
    .A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .B(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_nor2_1 _19414_ (.A(_04616_),
    .B(_04633_),
    .Y(_04650_));
 sg13g2_nor4_1 _19415_ (.A(_04588_),
    .B(_04602_),
    .C(_04616_),
    .D(_04633_),
    .Y(_04651_));
 sg13g2_o21ai_1 _19416_ (.B1(_04632_),
    .Y(_04652_),
    .A1(_04615_),
    .A2(_04631_));
 sg13g2_a221oi_1 _19417_ (.B2(_04586_),
    .C1(_04652_),
    .B1(_04651_),
    .A1(_04617_),
    .Y(_04653_),
    .A2(_04650_));
 sg13g2_or2_1 _19418_ (.X(_04654_),
    .B(_04653_),
    .A(_04649_));
 sg13g2_a21oi_1 _19419_ (.A1(_04649_),
    .A2(_04653_),
    .Y(_04655_),
    .B1(net4121));
 sg13g2_and3_2 _19420_ (.X(_04656_),
    .A(\soc_inst.cpu_core.id_pc[19] ),
    .B(\soc_inst.cpu_core.id_pc[20] ),
    .C(_04622_));
 sg13g2_a21oi_1 _19421_ (.A1(\soc_inst.cpu_core.id_pc[19] ),
    .A2(_04622_),
    .Y(_04657_),
    .B1(\soc_inst.cpu_core.id_pc[20] ));
 sg13g2_nor2_1 _19422_ (.A(_04656_),
    .B(_04657_),
    .Y(_04658_));
 sg13g2_a21oi_1 _19423_ (.A1(_04654_),
    .A2(_04655_),
    .Y(_04659_),
    .B1(net4900));
 sg13g2_a22oi_1 _19424_ (.Y(_04660_),
    .B1(_04658_),
    .B2(net3714),
    .A2(_04647_),
    .A1(net3712));
 sg13g2_a22oi_1 _19425_ (.Y(_01890_),
    .B1(_04659_),
    .B2(_04660_),
    .A2(_05715_),
    .A1(net4911));
 sg13g2_nor2_1 _19426_ (.A(\soc_inst.cpu_core.id_pc[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ),
    .Y(_04661_));
 sg13g2_xnor2_1 _19427_ (.Y(_04662_),
    .A(\soc_inst.cpu_core.id_pc[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_o21ai_1 _19428_ (.B1(_04645_),
    .Y(_04663_),
    .A1(\soc_inst.cpu_core.id_pc[20] ),
    .A2(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_o21ai_1 _19429_ (.B1(_04663_),
    .Y(_04664_),
    .A1(_05700_),
    .A2(_05701_));
 sg13g2_xnor2_1 _19430_ (.Y(_04665_),
    .A(_04662_),
    .B(_04664_));
 sg13g2_nand2_1 _19431_ (.Y(_04666_),
    .A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_xnor2_1 _19432_ (.Y(_04667_),
    .A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_nand3_1 _19433_ (.B(_04654_),
    .C(_04667_),
    .A(_04648_),
    .Y(_04668_));
 sg13g2_a21o_1 _19434_ (.A2(_04654_),
    .A1(_04648_),
    .B1(_04667_),
    .X(_04669_));
 sg13g2_nand3_1 _19435_ (.B(_04668_),
    .C(_04669_),
    .A(net4216),
    .Y(_04670_));
 sg13g2_xnor2_1 _19436_ (.Y(_04671_),
    .A(_05702_),
    .B(_04656_));
 sg13g2_a221oi_1 _19437_ (.B2(net3714),
    .C1(net4913),
    .B1(_04671_),
    .A1(net3712),
    .Y(_04672_),
    .A2(_04665_));
 sg13g2_a22oi_1 _19438_ (.Y(_01891_),
    .B1(_04670_),
    .B2(_04672_),
    .A2(_05716_),
    .A1(net4913));
 sg13g2_or2_1 _19439_ (.X(_04673_),
    .B(\soc_inst.cpu_core.id_imm[22] ),
    .A(\soc_inst.cpu_core.id_pc[22] ));
 sg13g2_and2_1 _19440_ (.A(\soc_inst.cpu_core.id_pc[22] ),
    .B(\soc_inst.cpu_core.id_imm[22] ),
    .X(_04674_));
 sg13g2_xor2_1 _19441_ (.B(\soc_inst.cpu_core.id_imm[22] ),
    .A(\soc_inst.cpu_core.id_pc[22] ),
    .X(_04675_));
 sg13g2_a22oi_1 _19442_ (.Y(_04676_),
    .B1(\soc_inst.cpu_core.id_pc[21] ),
    .B2(\soc_inst.cpu_core.id_imm[21] ),
    .A2(\soc_inst.cpu_core.id_imm[20] ),
    .A1(\soc_inst.cpu_core.id_pc[20] ));
 sg13g2_a21oi_1 _19443_ (.A1(_04663_),
    .A2(_04676_),
    .Y(_04677_),
    .B1(_04661_));
 sg13g2_xor2_1 _19444_ (.B(_04677_),
    .A(_04675_),
    .X(_04678_));
 sg13g2_nand2_1 _19445_ (.Y(_04679_),
    .A(\soc_inst.cpu_core.id_rs1_data[22] ),
    .B(\soc_inst.cpu_core.id_imm[22] ));
 sg13g2_xnor2_1 _19446_ (.Y(_04680_),
    .A(\soc_inst.cpu_core.id_rs1_data[22] ),
    .B(\soc_inst.cpu_core.id_imm[22] ));
 sg13g2_o21ai_1 _19447_ (.B1(_04666_),
    .Y(_04681_),
    .A1(_04648_),
    .A2(_04667_));
 sg13g2_a21o_1 _19448_ (.A2(_04669_),
    .A1(_04666_),
    .B1(_04680_),
    .X(_04682_));
 sg13g2_nand3_1 _19449_ (.B(_04669_),
    .C(_04680_),
    .A(_04666_),
    .Y(_04683_));
 sg13g2_nand3_1 _19450_ (.B(_04682_),
    .C(_04683_),
    .A(net4216),
    .Y(_04684_));
 sg13g2_nand3_1 _19451_ (.B(\soc_inst.cpu_core.id_pc[22] ),
    .C(_04656_),
    .A(\soc_inst.cpu_core.id_pc[21] ),
    .Y(_04685_));
 sg13g2_a21o_1 _19452_ (.A2(_04656_),
    .A1(\soc_inst.cpu_core.id_pc[21] ),
    .B1(\soc_inst.cpu_core.id_pc[22] ),
    .X(_04686_));
 sg13g2_and2_1 _19453_ (.A(_04685_),
    .B(_04686_),
    .X(_04687_));
 sg13g2_a221oi_1 _19454_ (.B2(net3714),
    .C1(net4910),
    .B1(_04687_),
    .A1(net3712),
    .Y(_04688_),
    .A2(_04678_));
 sg13g2_a22oi_1 _19455_ (.Y(_01892_),
    .B1(_04684_),
    .B2(_04688_),
    .A2(_05717_),
    .A1(net4914));
 sg13g2_nand2_1 _19456_ (.Y(_04689_),
    .A(_05704_),
    .B(_05705_));
 sg13g2_nor2_1 _19457_ (.A(_05704_),
    .B(_05705_),
    .Y(_04690_));
 sg13g2_xor2_1 _19458_ (.B(\soc_inst.cpu_core.id_imm[23] ),
    .A(\soc_inst.cpu_core.id_pc[23] ),
    .X(_04691_));
 sg13g2_a21oi_1 _19459_ (.A1(_04673_),
    .A2(_04677_),
    .Y(_04692_),
    .B1(_04674_));
 sg13g2_xor2_1 _19460_ (.B(_04692_),
    .A(_04691_),
    .X(_04693_));
 sg13g2_xnor2_1 _19461_ (.Y(_04694_),
    .A(\soc_inst.cpu_core.id_rs1_data[23] ),
    .B(\soc_inst.cpu_core.id_imm[23] ));
 sg13g2_nand3_1 _19462_ (.B(_04682_),
    .C(_04694_),
    .A(_04679_),
    .Y(_04695_));
 sg13g2_a21o_1 _19463_ (.A2(_04682_),
    .A1(_04679_),
    .B1(_04694_),
    .X(_04696_));
 sg13g2_nand3_1 _19464_ (.B(_04695_),
    .C(_04696_),
    .A(net4216),
    .Y(_04697_));
 sg13g2_o21ai_1 _19465_ (.B1(_04697_),
    .Y(_04698_),
    .A1(_09232_),
    .A2(_04693_));
 sg13g2_nor2_1 _19466_ (.A(_05704_),
    .B(_04685_),
    .Y(_04699_));
 sg13g2_xnor2_1 _19467_ (.Y(_04700_),
    .A(_05704_),
    .B(_04685_));
 sg13g2_a221oi_1 _19468_ (.B2(net3714),
    .C1(net4912),
    .B1(_04700_),
    .A1(_04333_),
    .Y(_04701_),
    .A2(_04693_));
 sg13g2_o21ai_1 _19469_ (.B1(_04701_),
    .Y(_04702_),
    .A1(net4109),
    .A2(_04698_));
 sg13g2_o21ai_1 _19470_ (.B1(_04702_),
    .Y(_01893_),
    .A1(net4751),
    .A2(_05718_));
 sg13g2_nor2_1 _19471_ (.A(_04646_),
    .B(_04662_),
    .Y(_04703_));
 sg13g2_and2_1 _19472_ (.A(_04675_),
    .B(_04691_),
    .X(_04704_));
 sg13g2_nand2_1 _19473_ (.Y(_04705_),
    .A(_04703_),
    .B(_04704_));
 sg13g2_a21o_1 _19474_ (.A2(_04644_),
    .A1(_04641_),
    .B1(_04705_),
    .X(_04706_));
 sg13g2_nor2_1 _19475_ (.A(_04661_),
    .B(_04676_),
    .Y(_04707_));
 sg13g2_a221oi_1 _19476_ (.B2(_04707_),
    .C1(_04690_),
    .B1(_04704_),
    .A1(_04674_),
    .Y(_04708_),
    .A2(_04689_));
 sg13g2_nand2_1 _19477_ (.Y(_04709_),
    .A(_04706_),
    .B(_04708_));
 sg13g2_a21o_1 _19478_ (.A2(_04699_),
    .A1(net4109),
    .B1(net3712),
    .X(_04710_));
 sg13g2_xor2_1 _19479_ (.B(_04709_),
    .A(\soc_inst.cpu_core.id_imm[24] ),
    .X(_04711_));
 sg13g2_nand2_1 _19480_ (.Y(_04712_),
    .A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .B(\soc_inst.cpu_core.id_imm[24] ));
 sg13g2_xnor2_1 _19481_ (.Y(_04713_),
    .A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .B(\soc_inst.cpu_core.id_imm[24] ));
 sg13g2_nor2_1 _19482_ (.A(_04680_),
    .B(_04694_),
    .Y(_04714_));
 sg13g2_or4_1 _19483_ (.A(_04649_),
    .B(_04667_),
    .C(_04680_),
    .D(_04694_),
    .X(_04715_));
 sg13g2_a21oi_1 _19484_ (.A1(_05668_),
    .A2(_05705_),
    .Y(_04716_),
    .B1(_04679_));
 sg13g2_a221oi_1 _19485_ (.B2(_04714_),
    .C1(_04716_),
    .B1(_04681_),
    .A1(\soc_inst.cpu_core.id_rs1_data[23] ),
    .Y(_04717_),
    .A2(\soc_inst.cpu_core.id_imm[23] ));
 sg13g2_o21ai_1 _19486_ (.B1(_04717_),
    .Y(_04718_),
    .A1(_04653_),
    .A2(_04715_));
 sg13g2_nand2b_1 _19487_ (.Y(_04719_),
    .B(_04718_),
    .A_N(_04713_));
 sg13g2_nand2b_1 _19488_ (.Y(_04720_),
    .B(_04713_),
    .A_N(_04718_));
 sg13g2_nand3_1 _19489_ (.B(_04719_),
    .C(_04720_),
    .A(net4216),
    .Y(_04721_));
 sg13g2_a221oi_1 _19490_ (.B2(_04711_),
    .C1(net4912),
    .B1(_04710_),
    .A1(net3715),
    .Y(_04722_),
    .A2(_04699_));
 sg13g2_a22oi_1 _19491_ (.Y(_01894_),
    .B1(_04721_),
    .B2(_04722_),
    .A2(_05774_),
    .A1(net4901));
 sg13g2_nor2_1 _19492_ (.A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .B(\soc_inst.cpu_core.id_imm[25] ),
    .Y(_04723_));
 sg13g2_nand2_1 _19493_ (.Y(_04724_),
    .A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .B(\soc_inst.cpu_core.id_imm[25] ));
 sg13g2_nand2b_1 _19494_ (.Y(_04725_),
    .B(_04724_),
    .A_N(_04723_));
 sg13g2_a21o_1 _19495_ (.A2(_04719_),
    .A1(_04712_),
    .B1(_04725_),
    .X(_04726_));
 sg13g2_nand3_1 _19496_ (.B(_04719_),
    .C(_04725_),
    .A(_04712_),
    .Y(_04727_));
 sg13g2_nand3_1 _19497_ (.B(_04726_),
    .C(_04727_),
    .A(net4217),
    .Y(_04728_));
 sg13g2_a21oi_1 _19498_ (.A1(\soc_inst.cpu_core.id_imm[24] ),
    .A2(_04709_),
    .Y(_04729_),
    .B1(\soc_inst.cpu_core.id_imm[25] ));
 sg13g2_nand2_1 _19499_ (.Y(_04730_),
    .A(\soc_inst.cpu_core.id_imm[24] ),
    .B(\soc_inst.cpu_core.id_imm[25] ));
 sg13g2_a21oi_1 _19500_ (.A1(_04706_),
    .A2(_04708_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_nor3_1 _19501_ (.A(_04407_),
    .B(_04729_),
    .C(_04731_),
    .Y(_04732_));
 sg13g2_nor2_1 _19502_ (.A(net4905),
    .B(_04732_),
    .Y(_04733_));
 sg13g2_a22oi_1 _19503_ (.Y(_01895_),
    .B1(_04728_),
    .B2(_04733_),
    .A2(_05776_),
    .A1(net4905));
 sg13g2_nor2_1 _19504_ (.A(net4751),
    .B(net936),
    .Y(_04734_));
 sg13g2_and2_1 _19505_ (.A(\soc_inst.cpu_core.id_imm[26] ),
    .B(_04731_),
    .X(_04735_));
 sg13g2_nor2_1 _19506_ (.A(\soc_inst.cpu_core.id_imm[26] ),
    .B(_04731_),
    .Y(_04736_));
 sg13g2_nor3_1 _19507_ (.A(_04407_),
    .B(_04735_),
    .C(_04736_),
    .Y(_04737_));
 sg13g2_nand2_1 _19508_ (.Y(_04738_),
    .A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .B(\soc_inst.cpu_core.id_imm[26] ));
 sg13g2_xnor2_1 _19509_ (.Y(_04739_),
    .A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .B(\soc_inst.cpu_core.id_imm[26] ));
 sg13g2_a21oi_1 _19510_ (.A1(_04724_),
    .A2(_04726_),
    .Y(_04740_),
    .B1(_04739_));
 sg13g2_nand3_1 _19511_ (.B(_04726_),
    .C(_04739_),
    .A(_04724_),
    .Y(_04741_));
 sg13g2_nor2_1 _19512_ (.A(net4121),
    .B(_04740_),
    .Y(_04742_));
 sg13g2_a21oi_1 _19513_ (.A1(_04741_),
    .A2(_04742_),
    .Y(_04743_),
    .B1(_04737_));
 sg13g2_a21oi_1 _19514_ (.A1(net4751),
    .A2(_04743_),
    .Y(_01896_),
    .B1(_04734_));
 sg13g2_nor2_1 _19515_ (.A(\soc_inst.cpu_core.id_rs1_data[27] ),
    .B(\soc_inst.cpu_core.id_imm[27] ),
    .Y(_04744_));
 sg13g2_nand2_1 _19516_ (.Y(_04745_),
    .A(\soc_inst.cpu_core.id_rs1_data[27] ),
    .B(\soc_inst.cpu_core.id_imm[27] ));
 sg13g2_nand2b_2 _19517_ (.Y(_04746_),
    .B(_04745_),
    .A_N(_04744_));
 sg13g2_a21oi_1 _19518_ (.A1(\soc_inst.cpu_core.id_rs1_data[26] ),
    .A2(\soc_inst.cpu_core.id_imm[26] ),
    .Y(_04747_),
    .B1(_04740_));
 sg13g2_a21oi_1 _19519_ (.A1(_04746_),
    .A2(_04747_),
    .Y(_04748_),
    .B1(net4121));
 sg13g2_o21ai_1 _19520_ (.B1(_04748_),
    .Y(_04749_),
    .A1(_04746_),
    .A2(_04747_));
 sg13g2_nor2_1 _19521_ (.A(\soc_inst.cpu_core.id_imm[27] ),
    .B(_04735_),
    .Y(_04750_));
 sg13g2_nand2_1 _19522_ (.Y(_04751_),
    .A(\soc_inst.cpu_core.id_imm[27] ),
    .B(_04735_));
 sg13g2_nor2_1 _19523_ (.A(_04407_),
    .B(_04750_),
    .Y(_04752_));
 sg13g2_a21oi_1 _19524_ (.A1(_04751_),
    .A2(_04752_),
    .Y(_04753_),
    .B1(net4905));
 sg13g2_a22oi_1 _19525_ (.Y(_01897_),
    .B1(_04749_),
    .B2(_04753_),
    .A2(_05777_),
    .A1(net4905));
 sg13g2_nand3_1 _19526_ (.B(\soc_inst.cpu_core.id_imm[28] ),
    .C(_04735_),
    .A(\soc_inst.cpu_core.id_imm[27] ),
    .Y(_04754_));
 sg13g2_nand2b_1 _19527_ (.Y(_04755_),
    .B(_04751_),
    .A_N(\soc_inst.cpu_core.id_imm[28] ));
 sg13g2_nor2_1 _19528_ (.A(_04739_),
    .B(_04746_),
    .Y(_04756_));
 sg13g2_o21ai_1 _19529_ (.B1(_04724_),
    .Y(_04757_),
    .A1(_04712_),
    .A2(_04723_));
 sg13g2_nor4_1 _19530_ (.A(_04713_),
    .B(_04725_),
    .C(_04739_),
    .D(_04746_),
    .Y(_04758_));
 sg13g2_o21ai_1 _19531_ (.B1(_04745_),
    .Y(_04759_),
    .A1(_04738_),
    .A2(_04744_));
 sg13g2_a221oi_1 _19532_ (.B2(_04718_),
    .C1(_04759_),
    .B1(_04758_),
    .A1(_04756_),
    .Y(_04760_),
    .A2(_04757_));
 sg13g2_and2_1 _19533_ (.A(\soc_inst.cpu_core.id_rs1_data[28] ),
    .B(\soc_inst.cpu_core.id_imm[28] ),
    .X(_04761_));
 sg13g2_xnor2_1 _19534_ (.Y(_04762_),
    .A(\soc_inst.cpu_core.id_rs1_data[28] ),
    .B(\soc_inst.cpu_core.id_imm[28] ));
 sg13g2_nor2_1 _19535_ (.A(_04760_),
    .B(_04762_),
    .Y(_04763_));
 sg13g2_a21o_1 _19536_ (.A2(_04762_),
    .A1(_04760_),
    .B1(net4121),
    .X(_04764_));
 sg13g2_nand3_1 _19537_ (.B(_04754_),
    .C(_04755_),
    .A(net3713),
    .Y(_04765_));
 sg13g2_o21ai_1 _19538_ (.B1(_04765_),
    .Y(_04766_),
    .A1(_04763_),
    .A2(_04764_));
 sg13g2_mux2_1 _19539_ (.A0(net1405),
    .A1(_04766_),
    .S(net4751),
    .X(_01898_));
 sg13g2_nand4_1 _19540_ (.B(\soc_inst.cpu_core.id_imm[28] ),
    .C(\soc_inst.cpu_core.id_imm[29] ),
    .A(\soc_inst.cpu_core.id_imm[27] ),
    .Y(_04767_),
    .D(_04735_));
 sg13g2_nand2b_1 _19541_ (.Y(_04768_),
    .B(_04754_),
    .A_N(\soc_inst.cpu_core.id_imm[29] ));
 sg13g2_nand3_1 _19542_ (.B(_04767_),
    .C(_04768_),
    .A(net3713),
    .Y(_04769_));
 sg13g2_xor2_1 _19543_ (.B(\soc_inst.cpu_core.id_imm[29] ),
    .A(\soc_inst.cpu_core.id_rs1_data[29] ),
    .X(_04770_));
 sg13g2_inv_1 _19544_ (.Y(_04771_),
    .A(_04770_));
 sg13g2_nor3_1 _19545_ (.A(_04760_),
    .B(_04762_),
    .C(_04771_),
    .Y(_04772_));
 sg13g2_nor3_1 _19546_ (.A(_04761_),
    .B(_04763_),
    .C(_04770_),
    .Y(_04773_));
 sg13g2_and2_1 _19547_ (.A(_04761_),
    .B(_04770_),
    .X(_04774_));
 sg13g2_nor4_1 _19548_ (.A(net4121),
    .B(_04772_),
    .C(_04773_),
    .D(_04774_),
    .Y(_04775_));
 sg13g2_nor2_1 _19549_ (.A(net4906),
    .B(_04775_),
    .Y(_04776_));
 sg13g2_a22oi_1 _19550_ (.Y(_01899_),
    .B1(_04769_),
    .B2(_04776_),
    .A2(_05780_),
    .A1(net4918));
 sg13g2_a21oi_1 _19551_ (.A1(\soc_inst.cpu_core.id_rs1_data[29] ),
    .A2(\soc_inst.cpu_core.id_imm[29] ),
    .Y(_04777_),
    .B1(_04774_));
 sg13g2_nor2b_1 _19552_ (.A(_04772_),
    .B_N(_04777_),
    .Y(_04778_));
 sg13g2_nand2_1 _19553_ (.Y(_04779_),
    .A(\soc_inst.cpu_core.id_rs1_data[30] ),
    .B(\soc_inst.cpu_core.id_imm[30] ));
 sg13g2_xnor2_1 _19554_ (.Y(_04780_),
    .A(\soc_inst.cpu_core.id_rs1_data[30] ),
    .B(\soc_inst.cpu_core.id_imm[30] ));
 sg13g2_or2_1 _19555_ (.X(_04781_),
    .B(_04780_),
    .A(_04778_));
 sg13g2_a21oi_1 _19556_ (.A1(_04778_),
    .A2(_04780_),
    .Y(_04782_),
    .B1(net4121));
 sg13g2_nor2_1 _19557_ (.A(_05706_),
    .B(_04767_),
    .Y(_04783_));
 sg13g2_a21oi_1 _19558_ (.A1(_05706_),
    .A2(_04767_),
    .Y(_04784_),
    .B1(_04407_));
 sg13g2_nand2b_1 _19559_ (.Y(_04785_),
    .B(_04784_),
    .A_N(_04783_));
 sg13g2_a21oi_1 _19560_ (.A1(_04781_),
    .A2(_04782_),
    .Y(_04786_),
    .B1(net4906));
 sg13g2_a22oi_1 _19561_ (.Y(_01900_),
    .B1(_04785_),
    .B2(_04786_),
    .A2(_05782_),
    .A1(net4906));
 sg13g2_xnor2_1 _19562_ (.Y(_04787_),
    .A(\soc_inst.cpu_core.id_rs1_data[31] ),
    .B(net993));
 sg13g2_a21o_1 _19563_ (.A2(_04781_),
    .A1(_04779_),
    .B1(_04787_),
    .X(_04788_));
 sg13g2_nand3_1 _19564_ (.B(_04781_),
    .C(_04787_),
    .A(_04779_),
    .Y(_04789_));
 sg13g2_nand3_1 _19565_ (.B(_04788_),
    .C(_04789_),
    .A(net4217),
    .Y(_04790_));
 sg13g2_xor2_1 _19566_ (.B(_04783_),
    .A(net993),
    .X(_04791_));
 sg13g2_a21oi_1 _19567_ (.A1(net3713),
    .A2(_04791_),
    .Y(_04792_),
    .B1(net4906));
 sg13g2_a22oi_1 _19568_ (.Y(_01901_),
    .B1(_04790_),
    .B2(_04792_),
    .A2(_05783_),
    .A1(net4918));
 sg13g2_nor3_2 _19569_ (.A(_09029_),
    .B(_09031_),
    .C(_09086_),
    .Y(_04793_));
 sg13g2_nand3_1 _19570_ (.B(net5078),
    .C(_04793_),
    .A(net4783),
    .Y(_04794_));
 sg13g2_a21oi_1 _19571_ (.A1(net5078),
    .A2(_04793_),
    .Y(_04795_),
    .B1(net4783));
 sg13g2_nor2b_1 _19572_ (.A(_09040_),
    .B_N(_06043_),
    .Y(_04796_));
 sg13g2_a21oi_1 _19573_ (.A1(_04793_),
    .A2(_04796_),
    .Y(_04797_),
    .B1(_04795_));
 sg13g2_and2_1 _19574_ (.A(_04794_),
    .B(_04797_),
    .X(_01902_));
 sg13g2_nand2_1 _19575_ (.Y(_04798_),
    .A(_09041_),
    .B(_09042_));
 sg13g2_a22oi_1 _19576_ (.Y(_01903_),
    .B1(_04798_),
    .B2(_04793_),
    .A2(_04794_),
    .A1(_05490_));
 sg13g2_nand2_1 _19577_ (.Y(_04799_),
    .A(_06718_),
    .B(_07217_));
 sg13g2_nand3_1 _19578_ (.B(net4090),
    .C(_07217_),
    .A(_06718_),
    .Y(_04800_));
 sg13g2_o21ai_1 _19579_ (.B1(_04800_),
    .Y(_04801_),
    .A1(net3797),
    .A2(net3786));
 sg13g2_nand2_1 _19580_ (.Y(_04802_),
    .A(net601),
    .B(net3744));
 sg13g2_a221oi_1 _19581_ (.B2(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .C1(net3993),
    .B1(net3990),
    .A1(\soc_inst.cpu_core.ex_alu_result[5] ),
    .Y(_04803_),
    .A2(net4052));
 sg13g2_nor2_1 _19582_ (.A(\soc_inst.cpu_core.ex_branch_target[5] ),
    .B(net4103),
    .Y(_04804_));
 sg13g2_nor2_1 _19583_ (.A(\soc_inst.cpu_core.ex_instr[5] ),
    .B(net4057),
    .Y(_04805_));
 sg13g2_nor4_2 _19584_ (.A(net3862),
    .B(_04803_),
    .C(_04804_),
    .Y(_04806_),
    .D(_04805_));
 sg13g2_nor2_1 _19585_ (.A(net3786),
    .B(_04806_),
    .Y(_04807_));
 sg13g2_a221oi_1 _19586_ (.B2(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .C1(net3842),
    .B1(net4170),
    .A1(net601),
    .Y(_04808_),
    .A2(_07605_));
 sg13g2_o21ai_1 _19587_ (.B1(_04802_),
    .Y(_01904_),
    .A1(_04807_),
    .A2(_04808_));
 sg13g2_nand2_1 _19588_ (.Y(_04809_),
    .A(net614),
    .B(net3744));
 sg13g2_a221oi_1 _19589_ (.B2(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .C1(net3993),
    .B1(net3989),
    .A1(\soc_inst.cpu_core.ex_alu_result[6] ),
    .Y(_04810_),
    .A2(net4052));
 sg13g2_nor2_1 _19590_ (.A(\soc_inst.cpu_core.ex_instr[6] ),
    .B(net4057),
    .Y(_04811_));
 sg13g2_nor2_1 _19591_ (.A(\soc_inst.cpu_core.ex_branch_target[6] ),
    .B(net4103),
    .Y(_04812_));
 sg13g2_nor4_2 _19592_ (.A(net3863),
    .B(_04810_),
    .C(_04811_),
    .Y(_04813_),
    .D(_04812_));
 sg13g2_nor2_1 _19593_ (.A(net3786),
    .B(_04813_),
    .Y(_04814_));
 sg13g2_a221oi_1 _19594_ (.B2(net614),
    .C1(net3842),
    .B1(_07612_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .Y(_04815_),
    .A2(net4169));
 sg13g2_o21ai_1 _19595_ (.B1(_04809_),
    .Y(_01905_),
    .A1(_04814_),
    .A2(_04815_));
 sg13g2_nand2_1 _19596_ (.Y(_04816_),
    .A(net578),
    .B(_04801_));
 sg13g2_a221oi_1 _19597_ (.B2(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .C1(net3994),
    .B1(net3990),
    .A1(\soc_inst.cpu_core.ex_alu_result[7] ),
    .Y(_04817_),
    .A2(net4052));
 sg13g2_a221oi_1 _19598_ (.B2(_05711_),
    .C1(_04817_),
    .B1(net4106),
    .A1(_05763_),
    .Y(_04818_),
    .A2(net4058));
 sg13g2_nor2_2 _19599_ (.A(net3785),
    .B(_04818_),
    .Y(_04819_));
 sg13g2_a221oi_1 _19600_ (.B2(net578),
    .C1(net3842),
    .B1(_08476_),
    .A1(net457),
    .Y(_04820_),
    .A2(net4172));
 sg13g2_o21ai_1 _19601_ (.B1(_04816_),
    .Y(_01906_),
    .A1(_04819_),
    .A2(_04820_));
 sg13g2_a221oi_1 _19602_ (.B2(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .C1(net3993),
    .B1(net3989),
    .A1(\soc_inst.cpu_core.ex_alu_result[8] ),
    .Y(_04821_),
    .A2(net4052));
 sg13g2_nand2b_1 _19603_ (.Y(_04822_),
    .B(net4106),
    .A_N(\soc_inst.cpu_core.ex_branch_target[8] ));
 sg13g2_o21ai_1 _19604_ (.B1(_04822_),
    .Y(_04823_),
    .A1(\soc_inst.cpu_core.ex_instr[8] ),
    .A2(net4057));
 sg13g2_or4_1 _19605_ (.A(net3861),
    .B(net3785),
    .C(_04821_),
    .D(_04823_),
    .X(_04824_));
 sg13g2_a22oi_1 _19606_ (.Y(_04825_),
    .B1(_07616_),
    .B2(net1431),
    .A2(net4170),
    .A1(\soc_inst.cpu_core.mem_rs1_data[8] ));
 sg13g2_o21ai_1 _19607_ (.B1(_04824_),
    .Y(_04826_),
    .A1(net3843),
    .A2(_04825_));
 sg13g2_a21o_1 _19608_ (.A2(net3744),
    .A1(net1431),
    .B1(_04826_),
    .X(_01907_));
 sg13g2_nand2_1 _19609_ (.Y(_04827_),
    .A(net476),
    .B(net3744));
 sg13g2_a221oi_1 _19610_ (.B2(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .C1(net3994),
    .B1(net3990),
    .A1(\soc_inst.cpu_core.ex_alu_result[9] ),
    .Y(_04828_),
    .A2(net4053));
 sg13g2_nor2_1 _19611_ (.A(\soc_inst.cpu_core.ex_instr[9] ),
    .B(net4057),
    .Y(_04829_));
 sg13g2_nor2_1 _19612_ (.A(\soc_inst.cpu_core.ex_branch_target[9] ),
    .B(net4102),
    .Y(_04830_));
 sg13g2_nor4_1 _19613_ (.A(net3861),
    .B(_04828_),
    .C(_04829_),
    .D(_04830_),
    .Y(_04831_));
 sg13g2_nor2_2 _19614_ (.A(net3785),
    .B(_04831_),
    .Y(_04832_));
 sg13g2_a221oi_1 _19615_ (.B2(net476),
    .C1(net3842),
    .B1(_07620_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .Y(_04833_),
    .A2(net4169));
 sg13g2_o21ai_1 _19616_ (.B1(_04827_),
    .Y(_01908_),
    .A1(_04832_),
    .A2(_04833_));
 sg13g2_a22oi_1 _19617_ (.Y(_04834_),
    .B1(net3989),
    .B2(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .A2(net4054),
    .A1(\soc_inst.cpu_core.ex_alu_result[10] ));
 sg13g2_nand2_1 _19618_ (.Y(_04835_),
    .A(\soc_inst.cpu_core.ex_instr[10] ),
    .B(net4102));
 sg13g2_a22oi_1 _19619_ (.Y(_04836_),
    .B1(_04835_),
    .B2(net3993),
    .A2(_04834_),
    .A1(net4057));
 sg13g2_and2_1 _19620_ (.A(\soc_inst.cpu_core.ex_branch_target[10] ),
    .B(net4106),
    .X(_04837_));
 sg13g2_o21ai_1 _19621_ (.B1(net3839),
    .Y(_04838_),
    .A1(_04836_),
    .A2(_04837_));
 sg13g2_a22oi_1 _19622_ (.Y(_04839_),
    .B1(_07624_),
    .B2(net1567),
    .A2(net4170),
    .A1(\soc_inst.cpu_core.mem_rs1_data[10] ));
 sg13g2_o21ai_1 _19623_ (.B1(_04838_),
    .Y(_04840_),
    .A1(net3843),
    .A2(_04839_));
 sg13g2_a21o_1 _19624_ (.A2(net3744),
    .A1(net1567),
    .B1(_04840_),
    .X(_01909_));
 sg13g2_nand2_1 _19625_ (.Y(_04841_),
    .A(net416),
    .B(net3744));
 sg13g2_a221oi_1 _19626_ (.B2(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .C1(net3994),
    .B1(net3990),
    .A1(\soc_inst.cpu_core.ex_alu_result[11] ),
    .Y(_04842_),
    .A2(net4054));
 sg13g2_nor2_1 _19627_ (.A(\soc_inst.cpu_core.ex_instr[11] ),
    .B(net4057),
    .Y(_04843_));
 sg13g2_nor2_1 _19628_ (.A(\soc_inst.cpu_core.ex_branch_target[11] ),
    .B(net4102),
    .Y(_04844_));
 sg13g2_nor4_1 _19629_ (.A(net3861),
    .B(_04842_),
    .C(_04843_),
    .D(_04844_),
    .Y(_04845_));
 sg13g2_nor2_2 _19630_ (.A(net3786),
    .B(_04845_),
    .Y(_04846_));
 sg13g2_a221oi_1 _19631_ (.B2(net416),
    .C1(net3842),
    .B1(_08487_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .Y(_04847_),
    .A2(net4171));
 sg13g2_o21ai_1 _19632_ (.B1(_04841_),
    .Y(_01910_),
    .A1(_04846_),
    .A2(_04847_));
 sg13g2_a22oi_1 _19633_ (.Y(_04848_),
    .B1(net3990),
    .B2(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .A2(net4053),
    .A1(\soc_inst.cpu_core.ex_alu_result[12] ));
 sg13g2_a21oi_1 _19634_ (.A1(\soc_inst.cpu_core.ex_funct3[0] ),
    .A2(net4058),
    .Y(_04849_),
    .B1(net4106));
 sg13g2_o21ai_1 _19635_ (.B1(_04849_),
    .Y(_04850_),
    .A1(net4058),
    .A2(_04848_));
 sg13g2_o21ai_1 _19636_ (.B1(_04850_),
    .Y(_04851_),
    .A1(\soc_inst.cpu_core.ex_branch_target[12] ),
    .A2(net4102));
 sg13g2_a221oi_1 _19637_ (.B2(net1520),
    .C1(net3842),
    .B1(_08491_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .Y(_04852_),
    .A2(net4171));
 sg13g2_a21oi_1 _19638_ (.A1(net3842),
    .A2(_04851_),
    .Y(_04853_),
    .B1(_04852_));
 sg13g2_a21o_1 _19639_ (.A2(net3744),
    .A1(net1520),
    .B1(_04853_),
    .X(_01911_));
 sg13g2_nand2_1 _19640_ (.Y(_04854_),
    .A(net458),
    .B(net3742));
 sg13g2_a221oi_1 _19641_ (.B2(\soc_inst.cpu_core.ex_exception_pc[13] ),
    .C1(net3995),
    .B1(net3991),
    .A1(\soc_inst.cpu_core.ex_alu_result[13] ),
    .Y(_04855_),
    .A2(net4050));
 sg13g2_nor2_1 _19642_ (.A(\soc_inst.cpu_core.ex_funct3[1] ),
    .B(_06640_),
    .Y(_04856_));
 sg13g2_nor2_1 _19643_ (.A(\soc_inst.cpu_core.ex_branch_target[13] ),
    .B(net4102),
    .Y(_04857_));
 sg13g2_nor4_1 _19644_ (.A(net3860),
    .B(_04855_),
    .C(_04856_),
    .D(_04857_),
    .Y(_04858_));
 sg13g2_nor2_1 _19645_ (.A(net3786),
    .B(_04858_),
    .Y(_04859_));
 sg13g2_a221oi_1 _19646_ (.B2(net458),
    .C1(net3844),
    .B1(_08495_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .Y(_04860_),
    .A2(net4172));
 sg13g2_o21ai_1 _19647_ (.B1(_04854_),
    .Y(_01912_),
    .A1(_04859_),
    .A2(_04860_));
 sg13g2_a22oi_1 _19648_ (.Y(_04861_),
    .B1(net3991),
    .B2(\soc_inst.cpu_core.ex_exception_pc[14] ),
    .A2(net4050),
    .A1(\soc_inst.cpu_core.ex_alu_result[14] ));
 sg13g2_nand2_1 _19649_ (.Y(_04862_),
    .A(\soc_inst.cpu_core.ex_funct3[2] ),
    .B(net4102));
 sg13g2_a22oi_1 _19650_ (.Y(_04863_),
    .B1(_04862_),
    .B2(net3994),
    .A2(_04861_),
    .A1(net4056));
 sg13g2_and2_1 _19651_ (.A(\soc_inst.cpu_core.ex_branch_target[14] ),
    .B(net4105),
    .X(_04864_));
 sg13g2_o21ai_1 _19652_ (.B1(net3839),
    .Y(_04865_),
    .A1(_04863_),
    .A2(_04864_));
 sg13g2_a22oi_1 _19653_ (.Y(_04866_),
    .B1(_08499_),
    .B2(net1445),
    .A2(net4171),
    .A1(\soc_inst.cpu_core.mem_rs1_data[14] ));
 sg13g2_o21ai_1 _19654_ (.B1(_04865_),
    .Y(_04867_),
    .A1(net3842),
    .A2(_04866_));
 sg13g2_a21o_1 _19655_ (.A2(net3744),
    .A1(net1445),
    .B1(_04867_),
    .X(_01913_));
 sg13g2_a22oi_1 _19656_ (.Y(_04868_),
    .B1(net3991),
    .B2(\soc_inst.cpu_core.ex_exception_pc[15] ),
    .A2(net4050),
    .A1(\soc_inst.cpu_core.ex_alu_result[15] ));
 sg13g2_nand2_1 _19657_ (.Y(_04869_),
    .A(\soc_inst.cpu_core.ex_instr[15] ),
    .B(net4102));
 sg13g2_a22oi_1 _19658_ (.Y(_04870_),
    .B1(_04869_),
    .B2(net3995),
    .A2(_04868_),
    .A1(net4056));
 sg13g2_and2_1 _19659_ (.A(\soc_inst.cpu_core.ex_branch_target[15] ),
    .B(net4105),
    .X(_04871_));
 sg13g2_o21ai_1 _19660_ (.B1(net3838),
    .Y(_04872_),
    .A1(_04870_),
    .A2(_04871_));
 sg13g2_a22oi_1 _19661_ (.Y(_04873_),
    .B1(_08503_),
    .B2(net2038),
    .A2(net4167),
    .A1(net932));
 sg13g2_o21ai_1 _19662_ (.B1(_04872_),
    .Y(_04874_),
    .A1(net3838),
    .A2(_04873_));
 sg13g2_a21o_1 _19663_ (.A2(net3742),
    .A1(net2038),
    .B1(_04874_),
    .X(_01914_));
 sg13g2_a221oi_1 _19664_ (.B2(\soc_inst.cpu_core.ex_exception_pc[16] ),
    .C1(net3992),
    .B1(net3988),
    .A1(\soc_inst.cpu_core.ex_alu_result[16] ),
    .Y(_04875_),
    .A2(net4049));
 sg13g2_nand2_1 _19665_ (.Y(_04876_),
    .A(_05712_),
    .B(net4104));
 sg13g2_o21ai_1 _19666_ (.B1(_04876_),
    .Y(_04877_),
    .A1(\soc_inst.cpu_core.ex_instr[16] ),
    .A2(net4055));
 sg13g2_or4_1 _19667_ (.A(net3860),
    .B(net3785),
    .C(_04875_),
    .D(_04877_),
    .X(_04878_));
 sg13g2_a22oi_1 _19668_ (.Y(_04879_),
    .B1(_08507_),
    .B2(net1271),
    .A2(net4168),
    .A1(\soc_inst.cpu_core.mem_rs1_data[16] ));
 sg13g2_o21ai_1 _19669_ (.B1(_04878_),
    .Y(_04880_),
    .A1(net3840),
    .A2(_04879_));
 sg13g2_a21o_1 _19670_ (.A2(net3743),
    .A1(net1271),
    .B1(_04880_),
    .X(_01915_));
 sg13g2_nand2_1 _19671_ (.Y(_04881_),
    .A(net509),
    .B(net3743));
 sg13g2_a221oi_1 _19672_ (.B2(\soc_inst.cpu_core.ex_exception_pc[17] ),
    .C1(net3992),
    .B1(net3988),
    .A1(\soc_inst.cpu_core.ex_alu_result[17] ),
    .Y(_04882_),
    .A2(net4049));
 sg13g2_nor2_1 _19673_ (.A(\soc_inst.cpu_core.ex_instr[17] ),
    .B(net4056),
    .Y(_04883_));
 sg13g2_nor2_1 _19674_ (.A(\soc_inst.cpu_core.ex_branch_target[17] ),
    .B(net4101),
    .Y(_04884_));
 sg13g2_nor4_1 _19675_ (.A(net3860),
    .B(_04882_),
    .C(_04883_),
    .D(_04884_),
    .Y(_04885_));
 sg13g2_nor2_2 _19676_ (.A(net3785),
    .B(_04885_),
    .Y(_04886_));
 sg13g2_a221oi_1 _19677_ (.B2(net509),
    .C1(net3840),
    .B1(_08511_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .Y(_04887_),
    .A2(net4167));
 sg13g2_o21ai_1 _19678_ (.B1(_04881_),
    .Y(_01916_),
    .A1(_04886_),
    .A2(_04887_));
 sg13g2_a221oi_1 _19679_ (.B2(net1246),
    .C1(net3992),
    .B1(net3988),
    .A1(\soc_inst.cpu_core.ex_alu_result[18] ),
    .Y(_04888_),
    .A2(net4049));
 sg13g2_nand2_1 _19680_ (.Y(_04889_),
    .A(_05713_),
    .B(net4104));
 sg13g2_o21ai_1 _19681_ (.B1(_04889_),
    .Y(_04890_),
    .A1(\soc_inst.cpu_core.ex_instr[18] ),
    .A2(net4055));
 sg13g2_or4_1 _19682_ (.A(net3860),
    .B(net3785),
    .C(_04888_),
    .D(_04890_),
    .X(_04891_));
 sg13g2_a22oi_1 _19683_ (.Y(_04892_),
    .B1(_08515_),
    .B2(net2022),
    .A2(net4167),
    .A1(\soc_inst.cpu_core.mem_rs1_data[18] ));
 sg13g2_o21ai_1 _19684_ (.B1(_04891_),
    .Y(_04893_),
    .A1(net3837),
    .A2(_04892_));
 sg13g2_a21o_1 _19685_ (.A2(net3742),
    .A1(net2022),
    .B1(_04893_),
    .X(_01917_));
 sg13g2_nand2_1 _19686_ (.Y(_04894_),
    .A(net576),
    .B(net3742));
 sg13g2_a221oi_1 _19687_ (.B2(\soc_inst.cpu_core.ex_exception_pc[19] ),
    .C1(net3992),
    .B1(net3988),
    .A1(\soc_inst.cpu_core.ex_alu_result[19] ),
    .Y(_04895_),
    .A2(net4049));
 sg13g2_nor2_1 _19688_ (.A(\soc_inst.cpu_core.ex_instr[19] ),
    .B(net4055),
    .Y(_04896_));
 sg13g2_nor2_1 _19689_ (.A(\soc_inst.cpu_core.ex_branch_target[19] ),
    .B(net4103),
    .Y(_04897_));
 sg13g2_nor4_1 _19690_ (.A(net3860),
    .B(_04895_),
    .C(_04896_),
    .D(_04897_),
    .Y(_04898_));
 sg13g2_nor2_1 _19691_ (.A(net3785),
    .B(_04898_),
    .Y(_04899_));
 sg13g2_a221oi_1 _19692_ (.B2(net576),
    .C1(net3838),
    .B1(_08519_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .Y(_04900_),
    .A2(net4167));
 sg13g2_o21ai_1 _19693_ (.B1(_04894_),
    .Y(_01918_),
    .A1(_04899_),
    .A2(_04900_));
 sg13g2_nand2_1 _19694_ (.Y(_04901_),
    .A(net455),
    .B(net3742));
 sg13g2_a221oi_1 _19695_ (.B2(\soc_inst.cpu_core.ex_exception_pc[20] ),
    .C1(net3992),
    .B1(net3988),
    .A1(\soc_inst.cpu_core.ex_alu_result[20] ),
    .Y(_04902_),
    .A2(net4049));
 sg13g2_nor2_1 _19696_ (.A(\soc_inst.cpu_core.ex_instr[20] ),
    .B(net4055),
    .Y(_04903_));
 sg13g2_nor2_1 _19697_ (.A(\soc_inst.cpu_core.ex_branch_target[20] ),
    .B(net4101),
    .Y(_04904_));
 sg13g2_nor4_1 _19698_ (.A(net3860),
    .B(_04902_),
    .C(_04903_),
    .D(_04904_),
    .Y(_04905_));
 sg13g2_nor2_1 _19699_ (.A(net3785),
    .B(_04905_),
    .Y(_04906_));
 sg13g2_a221oi_1 _19700_ (.B2(net455),
    .C1(net3843),
    .B1(_08523_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .Y(_04907_),
    .A2(net4167));
 sg13g2_o21ai_1 _19701_ (.B1(_04901_),
    .Y(_01919_),
    .A1(_04906_),
    .A2(_04907_));
 sg13g2_a22oi_1 _19702_ (.Y(_04908_),
    .B1(net3988),
    .B2(\soc_inst.cpu_core.ex_exception_pc[21] ),
    .A2(net4049),
    .A1(\soc_inst.cpu_core.ex_alu_result[21] ));
 sg13g2_nand2_1 _19703_ (.Y(_04909_),
    .A(\soc_inst.cpu_core.ex_instr[21] ),
    .B(net4101));
 sg13g2_a22oi_1 _19704_ (.Y(_04910_),
    .B1(_04909_),
    .B2(net3992),
    .A2(_04908_),
    .A1(net4055));
 sg13g2_nor2_1 _19705_ (.A(_05716_),
    .B(net4101),
    .Y(_04911_));
 sg13g2_o21ai_1 _19706_ (.B1(net3837),
    .Y(_04912_),
    .A1(_04910_),
    .A2(_04911_));
 sg13g2_a22oi_1 _19707_ (.Y(_04913_),
    .B1(_08527_),
    .B2(net1851),
    .A2(net4167),
    .A1(\soc_inst.cpu_core.mem_rs1_data[21] ));
 sg13g2_o21ai_1 _19708_ (.B1(_04912_),
    .Y(_04914_),
    .A1(net3837),
    .A2(_04913_));
 sg13g2_a21o_1 _19709_ (.A2(net3742),
    .A1(net1851),
    .B1(_04914_),
    .X(_01920_));
 sg13g2_a22oi_1 _19710_ (.Y(_04915_),
    .B1(net3988),
    .B2(\soc_inst.cpu_core.ex_exception_pc[22] ),
    .A2(net4049),
    .A1(\soc_inst.cpu_core.ex_alu_result[22] ));
 sg13g2_nand2_1 _19711_ (.Y(_04916_),
    .A(\soc_inst.cpu_core.ex_instr[22] ),
    .B(net4101));
 sg13g2_a22oi_1 _19712_ (.Y(_04917_),
    .B1(_04916_),
    .B2(net3992),
    .A2(_04915_),
    .A1(net4056));
 sg13g2_nor2_1 _19713_ (.A(_05717_),
    .B(net4101),
    .Y(_04918_));
 sg13g2_o21ai_1 _19714_ (.B1(net3837),
    .Y(_04919_),
    .A1(_04917_),
    .A2(_04918_));
 sg13g2_a22oi_1 _19715_ (.Y(_04920_),
    .B1(_08531_),
    .B2(net2076),
    .A2(net4167),
    .A1(\soc_inst.cpu_core.mem_rs1_data[22] ));
 sg13g2_o21ai_1 _19716_ (.B1(_04919_),
    .Y(_04921_),
    .A1(net3838),
    .A2(_04920_));
 sg13g2_a21o_1 _19717_ (.A2(net3742),
    .A1(net2076),
    .B1(_04921_),
    .X(_01921_));
 sg13g2_a22oi_1 _19718_ (.Y(_04922_),
    .B1(net3988),
    .B2(\soc_inst.cpu_core.ex_exception_pc[23] ),
    .A2(net4049),
    .A1(\soc_inst.cpu_core.ex_alu_result[23] ));
 sg13g2_nand2_1 _19719_ (.Y(_04923_),
    .A(\soc_inst.cpu_core.ex_instr[23] ),
    .B(net4101));
 sg13g2_a22oi_1 _19720_ (.Y(_04924_),
    .B1(_04923_),
    .B2(net3992),
    .A2(_04922_),
    .A1(net4056));
 sg13g2_and2_1 _19721_ (.A(net1069),
    .B(net4105),
    .X(_04925_));
 sg13g2_o21ai_1 _19722_ (.B1(net3837),
    .Y(_04926_),
    .A1(_04924_),
    .A2(_04925_));
 sg13g2_a22oi_1 _19723_ (.Y(_04927_),
    .B1(_08535_),
    .B2(net1940),
    .A2(net4167),
    .A1(\soc_inst.cpu_core.mem_rs1_data[23] ));
 sg13g2_o21ai_1 _19724_ (.B1(_04926_),
    .Y(_04928_),
    .A1(net3837),
    .A2(_04927_));
 sg13g2_a21o_1 _19725_ (.A2(net3742),
    .A1(net1940),
    .B1(_04928_),
    .X(_01922_));
 sg13g2_nor2_1 _19726_ (.A(_05774_),
    .B(net4103),
    .Y(_04929_));
 sg13g2_a221oi_1 _19727_ (.B2(\soc_inst.cpu_core.ex_alu_result[24] ),
    .C1(_04929_),
    .B1(net4051),
    .A1(\soc_inst.cpu_core.ex_instr[24] ),
    .Y(_04930_),
    .A2(net4058));
 sg13g2_a221oi_1 _19728_ (.B2(net1503),
    .C1(net3841),
    .B1(_08540_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .Y(_04931_),
    .A2(net4168));
 sg13g2_a21oi_1 _19729_ (.A1(net3841),
    .A2(_04930_),
    .Y(_04932_),
    .B1(_04931_));
 sg13g2_a21o_1 _19730_ (.A2(net3745),
    .A1(net1503),
    .B1(_04932_),
    .X(_01923_));
 sg13g2_or2_1 _19731_ (.X(_04933_),
    .B(net1005),
    .A(net2348));
 sg13g2_a22oi_1 _19732_ (.Y(_04934_),
    .B1(_08544_),
    .B2(_04933_),
    .A2(net4226),
    .A1(net1005));
 sg13g2_a22oi_1 _19733_ (.Y(_04935_),
    .B1(net4051),
    .B2(\soc_inst.cpu_core.ex_alu_result[25] ),
    .A2(net4104),
    .A1(\soc_inst.cpu_core.ex_branch_target[25] ));
 sg13g2_o21ai_1 _19734_ (.B1(_04935_),
    .Y(_04936_),
    .A1(_05775_),
    .A2(net4055));
 sg13g2_a22oi_1 _19735_ (.Y(_04937_),
    .B1(_04936_),
    .B2(net3840),
    .A2(net3743),
    .A1(net2348));
 sg13g2_o21ai_1 _19736_ (.B1(_04937_),
    .Y(_01924_),
    .A1(net3840),
    .A2(_04934_));
 sg13g2_or2_1 _19737_ (.X(_04938_),
    .B(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .A(net2594));
 sg13g2_a22oi_1 _19738_ (.Y(_04939_),
    .B1(_08548_),
    .B2(_04938_),
    .A2(net4227),
    .A1(\soc_inst.cpu_core.mem_rs1_data[26] ));
 sg13g2_nand2_1 _19739_ (.Y(_04940_),
    .A(\soc_inst.cpu_core.ex_alu_result[26] ),
    .B(net4054));
 sg13g2_a22oi_1 _19740_ (.Y(_04941_),
    .B1(net4104),
    .B2(\soc_inst.cpu_core.ex_branch_target[26] ),
    .A2(net4058),
    .A1(net2261));
 sg13g2_nand2_2 _19741_ (.Y(_04942_),
    .A(_04940_),
    .B(_04941_));
 sg13g2_a22oi_1 _19742_ (.Y(_04943_),
    .B1(_04942_),
    .B2(net3841),
    .A2(net3745),
    .A1(net2594));
 sg13g2_o21ai_1 _19743_ (.B1(net2595),
    .Y(_01925_),
    .A1(net3841),
    .A2(_04939_));
 sg13g2_or2_1 _19744_ (.X(_04944_),
    .B(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .A(net2398));
 sg13g2_a22oi_1 _19745_ (.Y(_04945_),
    .B1(_08552_),
    .B2(_04944_),
    .A2(net4226),
    .A1(\soc_inst.cpu_core.mem_rs1_data[27] ));
 sg13g2_nand2_1 _19746_ (.Y(_04946_),
    .A(\soc_inst.cpu_core.ex_alu_result[27] ),
    .B(net4051));
 sg13g2_a22oi_1 _19747_ (.Y(_04947_),
    .B1(net4104),
    .B2(\soc_inst.cpu_core.ex_branch_target[27] ),
    .A2(net4058),
    .A1(\soc_inst.cpu_core.ex_funct7[2] ));
 sg13g2_nand2_2 _19748_ (.Y(_04948_),
    .A(_04946_),
    .B(_04947_));
 sg13g2_a22oi_1 _19749_ (.Y(_04949_),
    .B1(_04948_),
    .B2(net3840),
    .A2(net3743),
    .A1(net2398));
 sg13g2_o21ai_1 _19750_ (.B1(net2399),
    .Y(_01926_),
    .A1(net3840),
    .A2(_04945_));
 sg13g2_nand2_1 _19751_ (.Y(_04950_),
    .A(\soc_inst.cpu_core.ex_funct7[3] ),
    .B(net4058));
 sg13g2_a22oi_1 _19752_ (.Y(_04951_),
    .B1(net4051),
    .B2(\soc_inst.cpu_core.ex_alu_result[28] ),
    .A2(net4104),
    .A1(\soc_inst.cpu_core.ex_branch_target[28] ));
 sg13g2_nor2_1 _19753_ (.A(net1669),
    .B(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .Y(_04952_));
 sg13g2_a21oi_1 _19754_ (.A1(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .A2(net4226),
    .Y(_04953_),
    .B1(_08556_));
 sg13g2_nand3_1 _19755_ (.B(_04950_),
    .C(_04951_),
    .A(net3837),
    .Y(_04954_));
 sg13g2_o21ai_1 _19756_ (.B1(net3786),
    .Y(_04955_),
    .A1(_04952_),
    .A2(_04953_));
 sg13g2_a22oi_1 _19757_ (.Y(_04956_),
    .B1(_04954_),
    .B2(_04955_),
    .A2(net3743),
    .A1(net1669));
 sg13g2_inv_1 _19758_ (.Y(_01927_),
    .A(net1670));
 sg13g2_or2_1 _19759_ (.X(_04957_),
    .B(net1095),
    .A(net2418));
 sg13g2_a22oi_1 _19760_ (.Y(_04958_),
    .B1(_08560_),
    .B2(_04957_),
    .A2(net4226),
    .A1(net1095));
 sg13g2_a22oi_1 _19761_ (.Y(_04959_),
    .B1(net4051),
    .B2(\soc_inst.cpu_core.ex_alu_result[29] ),
    .A2(net4104),
    .A1(\soc_inst.cpu_core.ex_branch_target[29] ));
 sg13g2_o21ai_1 _19762_ (.B1(_04959_),
    .Y(_04960_),
    .A1(_05778_),
    .A2(net4055));
 sg13g2_a22oi_1 _19763_ (.Y(_04961_),
    .B1(_04960_),
    .B2(net3840),
    .A2(net3743),
    .A1(net2418));
 sg13g2_o21ai_1 _19764_ (.B1(_04961_),
    .Y(_01928_),
    .A1(net3840),
    .A2(_04958_));
 sg13g2_or2_1 _19765_ (.X(_04962_),
    .B(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .A(net2546));
 sg13g2_a22oi_1 _19766_ (.Y(_04963_),
    .B1(_08564_),
    .B2(_04962_),
    .A2(net4227),
    .A1(\soc_inst.cpu_core.mem_rs1_data[30] ));
 sg13g2_a22oi_1 _19767_ (.Y(_04964_),
    .B1(net4051),
    .B2(\soc_inst.cpu_core.ex_alu_result[30] ),
    .A2(net4104),
    .A1(\soc_inst.cpu_core.ex_branch_target[30] ));
 sg13g2_o21ai_1 _19768_ (.B1(_04964_),
    .Y(_04965_),
    .A1(_05781_),
    .A2(net4056));
 sg13g2_a22oi_1 _19769_ (.Y(_04966_),
    .B1(_04965_),
    .B2(net3841),
    .A2(net3743),
    .A1(net2546));
 sg13g2_o21ai_1 _19770_ (.B1(_04966_),
    .Y(_01929_),
    .A1(net3841),
    .A2(_04963_));
 sg13g2_nor2_1 _19771_ (.A(net1933),
    .B(net4879),
    .Y(_04967_));
 sg13g2_a21oi_1 _19772_ (.A1(net4879),
    .A2(net4227),
    .Y(_04968_),
    .B1(_08568_));
 sg13g2_nand2_1 _19773_ (.Y(_04969_),
    .A(\soc_inst.cpu_core.ex_funct7[6] ),
    .B(net4058));
 sg13g2_a22oi_1 _19774_ (.Y(_04970_),
    .B1(net4051),
    .B2(\soc_inst.cpu_core.ex_alu_result[31] ),
    .A2(net4105),
    .A1(\soc_inst.cpu_core.ex_branch_target[31] ));
 sg13g2_nand3_1 _19775_ (.B(_04969_),
    .C(_04970_),
    .A(net3837),
    .Y(_04971_));
 sg13g2_o21ai_1 _19776_ (.B1(net3786),
    .Y(_04972_),
    .A1(_04967_),
    .A2(_04968_));
 sg13g2_a22oi_1 _19777_ (.Y(_04973_),
    .B1(_04971_),
    .B2(_04972_),
    .A2(net3743),
    .A1(net1933));
 sg13g2_inv_1 _19778_ (.Y(_01930_),
    .A(net1934));
 sg13g2_a21oi_1 _19779_ (.A1(_07609_),
    .A2(net3765),
    .Y(_04974_),
    .B1(net387));
 sg13g2_and2_1 _19780_ (.A(net4698),
    .B(net3762),
    .X(_04975_));
 sg13g2_a21oi_1 _19781_ (.A1(_08468_),
    .A2(net3740),
    .Y(_01931_),
    .B1(net388));
 sg13g2_nand2_1 _19782_ (.Y(_04976_),
    .A(_07614_),
    .B(net3765));
 sg13g2_a22oi_1 _19783_ (.Y(_01932_),
    .B1(_04976_),
    .B2(_05617_),
    .A2(net3740),
    .A1(_08472_));
 sg13g2_a21oi_1 _19784_ (.A1(net3765),
    .A2(_08473_),
    .Y(_04977_),
    .B1(net547));
 sg13g2_a21oi_1 _19785_ (.A1(_08477_),
    .A2(net3740),
    .Y(_01933_),
    .B1(_04977_));
 sg13g2_a21oi_1 _19786_ (.A1(_07618_),
    .A2(net3765),
    .Y(_04978_),
    .B1(net506));
 sg13g2_a21oi_1 _19787_ (.A1(_08479_),
    .A2(net3740),
    .Y(_01934_),
    .B1(net507));
 sg13g2_a21oi_1 _19788_ (.A1(_07622_),
    .A2(net3766),
    .Y(_04979_),
    .B1(net664));
 sg13g2_a21oi_1 _19789_ (.A1(_08481_),
    .A2(net3740),
    .Y(_01935_),
    .B1(net665));
 sg13g2_nand2_1 _19790_ (.Y(_04980_),
    .A(_07626_),
    .B(net3766));
 sg13g2_a22oi_1 _19791_ (.Y(_01936_),
    .B1(_04980_),
    .B2(_05622_),
    .A2(net3741),
    .A1(_08483_));
 sg13g2_a21oi_1 _19792_ (.A1(net3765),
    .A2(_08484_),
    .Y(_04981_),
    .B1(net450));
 sg13g2_a21oi_1 _19793_ (.A1(_08488_),
    .A2(net3740),
    .Y(_01937_),
    .B1(net451));
 sg13g2_nand2_1 _19794_ (.Y(_04982_),
    .A(net3763),
    .B(_08489_));
 sg13g2_a22oi_1 _19795_ (.Y(_01938_),
    .B1(_04982_),
    .B2(_05625_),
    .A2(net3740),
    .A1(_08492_));
 sg13g2_a21oi_1 _19796_ (.A1(net3762),
    .A2(_08493_),
    .Y(_04983_),
    .B1(net945));
 sg13g2_a21oi_1 _19797_ (.A1(_08496_),
    .A2(net3741),
    .Y(_01939_),
    .B1(_04983_));
 sg13g2_a21oi_1 _19798_ (.A1(net3766),
    .A2(_08497_),
    .Y(_04984_),
    .B1(net538));
 sg13g2_a21oi_1 _19799_ (.A1(_08500_),
    .A2(net3740),
    .Y(_01940_),
    .B1(net539));
 sg13g2_nand2_1 _19800_ (.Y(_04985_),
    .A(net3762),
    .B(_08501_));
 sg13g2_a22oi_1 _19801_ (.Y(_01941_),
    .B1(_04985_),
    .B2(_05630_),
    .A2(net3739),
    .A1(_08504_));
 sg13g2_nand2_1 _19802_ (.Y(_04986_),
    .A(net3763),
    .B(_08505_));
 sg13g2_a22oi_1 _19803_ (.Y(_01942_),
    .B1(_04986_),
    .B2(_05632_),
    .A2(net3741),
    .A1(_08508_));
 sg13g2_nand2_1 _19804_ (.Y(_04987_),
    .A(net3763),
    .B(_08509_));
 sg13g2_a22oi_1 _19805_ (.Y(_01943_),
    .B1(_04987_),
    .B2(_05634_),
    .A2(net3739),
    .A1(_08512_));
 sg13g2_nand2_1 _19806_ (.Y(_04988_),
    .A(net3762),
    .B(_08513_));
 sg13g2_a22oi_1 _19807_ (.Y(_01944_),
    .B1(_04988_),
    .B2(_05636_),
    .A2(net3739),
    .A1(_08516_));
 sg13g2_nand2_1 _19808_ (.Y(_04989_),
    .A(net3762),
    .B(_08517_));
 sg13g2_a22oi_1 _19809_ (.Y(_01945_),
    .B1(_04989_),
    .B2(_05638_),
    .A2(net3739),
    .A1(_08520_));
 sg13g2_nand2_1 _19810_ (.Y(_04990_),
    .A(net3763),
    .B(_08521_));
 sg13g2_a22oi_1 _19811_ (.Y(_01946_),
    .B1(_04990_),
    .B2(_05640_),
    .A2(net3739),
    .A1(_08524_));
 sg13g2_nand2_1 _19812_ (.Y(_04991_),
    .A(net3762),
    .B(_08525_));
 sg13g2_a22oi_1 _19813_ (.Y(_01947_),
    .B1(_04991_),
    .B2(_05642_),
    .A2(net3739),
    .A1(_08528_));
 sg13g2_nand2_1 _19814_ (.Y(_04992_),
    .A(net3762),
    .B(_08529_));
 sg13g2_a22oi_1 _19815_ (.Y(_01948_),
    .B1(_04992_),
    .B2(_05644_),
    .A2(net3739),
    .A1(_08532_));
 sg13g2_nand2_1 _19816_ (.Y(_04993_),
    .A(net3762),
    .B(_08533_));
 sg13g2_a22oi_1 _19817_ (.Y(_01949_),
    .B1(_04993_),
    .B2(_05646_),
    .A2(net3739),
    .A1(_08536_));
 sg13g2_nor2_2 _19818_ (.A(_06692_),
    .B(_04799_),
    .Y(_04994_));
 sg13g2_nand3_1 _19819_ (.B(_06718_),
    .C(_07217_),
    .A(net4192),
    .Y(_04995_));
 sg13g2_nand2_1 _19820_ (.Y(_04996_),
    .A(_06747_),
    .B(_04995_));
 sg13g2_nand2_1 _19821_ (.Y(_04997_),
    .A(net1090),
    .B(net3719));
 sg13g2_a221oi_1 _19822_ (.B2(\soc_inst.cpu_core.id_pc[5] ),
    .C1(net3788),
    .B1(net3752),
    .A1(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .Y(_04998_),
    .A2(net3859));
 sg13g2_a221oi_1 _19823_ (.B2(net812),
    .C1(net3852),
    .B1(net4172),
    .A1(net1090),
    .Y(_04999_),
    .A2(_07605_));
 sg13g2_o21ai_1 _19824_ (.B1(_04997_),
    .Y(_01950_),
    .A1(_04998_),
    .A2(_04999_));
 sg13g2_nand2_1 _19825_ (.Y(_05000_),
    .A(_05683_),
    .B(net3753));
 sg13g2_o21ai_1 _19826_ (.B1(_05000_),
    .Y(_05001_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .A2(net3861));
 sg13g2_a22oi_1 _19827_ (.Y(_05002_),
    .B1(_07612_),
    .B2(net1435),
    .A2(net4170),
    .A1(\soc_inst.cpu_core.mem_rs1_data[6] ));
 sg13g2_mux2_1 _19828_ (.A0(_05001_),
    .A1(_05002_),
    .S(net3788),
    .X(_05003_));
 sg13g2_a22oi_1 _19829_ (.Y(_01951_),
    .B1(_05003_),
    .B2(_04995_),
    .A2(net3719),
    .A1(_05616_));
 sg13g2_nand2_1 _19830_ (.Y(_05004_),
    .A(_05684_),
    .B(net3752));
 sg13g2_o21ai_1 _19831_ (.B1(_05004_),
    .Y(_05005_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .A2(net3862));
 sg13g2_o21ai_1 _19832_ (.B1(_04995_),
    .Y(_05006_),
    .A1(net3788),
    .A2(_05005_));
 sg13g2_o21ai_1 _19833_ (.B1(_05006_),
    .Y(_05007_),
    .A1(net2683),
    .A2(net3796));
 sg13g2_a21oi_1 _19834_ (.A1(net2683),
    .A2(net4622),
    .Y(_05008_),
    .B1(_08473_));
 sg13g2_nand2_1 _19835_ (.Y(_05009_),
    .A(net4192),
    .B(net4172));
 sg13g2_or4_1 _19836_ (.A(_05618_),
    .B(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .C(_06692_),
    .D(net4609),
    .X(_05010_));
 sg13g2_o21ai_1 _19837_ (.B1(_05010_),
    .Y(_05011_),
    .A1(_05008_),
    .A2(_05009_));
 sg13g2_nand3_1 _19838_ (.B(net3946),
    .C(_05011_),
    .A(net4710),
    .Y(_05012_));
 sg13g2_a22oi_1 _19839_ (.Y(_01952_),
    .B1(_05007_),
    .B2(_05012_),
    .A2(net3755),
    .A1(_05618_));
 sg13g2_a221oi_1 _19840_ (.B2(_05685_),
    .C1(net3788),
    .B1(net3753),
    .A1(_05742_),
    .Y(_05013_),
    .A2(_06655_));
 sg13g2_a22oi_1 _19841_ (.Y(_05014_),
    .B1(_07616_),
    .B2(net1016),
    .A2(net4169),
    .A1(\soc_inst.cpu_core.mem_rs1_data[8] ));
 sg13g2_o21ai_1 _19842_ (.B1(_04995_),
    .Y(_05015_),
    .A1(net3852),
    .A2(_05014_));
 sg13g2_nor2_1 _19843_ (.A(_05013_),
    .B(_05015_),
    .Y(_05016_));
 sg13g2_a21oi_1 _19844_ (.A1(_05619_),
    .A2(net3719),
    .Y(_01953_),
    .B1(_05016_));
 sg13g2_nand2_1 _19845_ (.Y(_05017_),
    .A(_05686_),
    .B(net3753));
 sg13g2_o21ai_1 _19846_ (.B1(_05017_),
    .Y(_05018_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .A2(net3862));
 sg13g2_a22oi_1 _19847_ (.Y(_05019_),
    .B1(_07620_),
    .B2(net999),
    .A2(net4172),
    .A1(\soc_inst.cpu_core.mem_rs1_data[9] ));
 sg13g2_mux2_1 _19848_ (.A0(_05018_),
    .A1(_05019_),
    .S(net3788),
    .X(_05020_));
 sg13g2_a22oi_1 _19849_ (.Y(_01954_),
    .B1(_05020_),
    .B2(_04995_),
    .A2(net3719),
    .A1(_05620_));
 sg13g2_nand2_1 _19850_ (.Y(_05021_),
    .A(_05687_),
    .B(net3753));
 sg13g2_o21ai_1 _19851_ (.B1(_05021_),
    .Y(_05022_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .A2(net3861));
 sg13g2_a22oi_1 _19852_ (.Y(_05023_),
    .B1(_07624_),
    .B2(net1208),
    .A2(net4169),
    .A1(\soc_inst.cpu_core.mem_rs1_data[10] ));
 sg13g2_mux2_1 _19853_ (.A0(_05022_),
    .A1(_05023_),
    .S(net3788),
    .X(_05024_));
 sg13g2_a22oi_1 _19854_ (.Y(_01955_),
    .B1(_05024_),
    .B2(_04995_),
    .A2(net3719),
    .A1(_05621_));
 sg13g2_nand2_1 _19855_ (.Y(_05025_),
    .A(_05689_),
    .B(net3752));
 sg13g2_o21ai_1 _19856_ (.B1(_05025_),
    .Y(_05026_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .A2(net3861));
 sg13g2_o21ai_1 _19857_ (.B1(_04995_),
    .Y(_05027_),
    .A1(net3789),
    .A2(_05026_));
 sg13g2_o21ai_1 _19858_ (.B1(_05027_),
    .Y(_05028_),
    .A1(net2484),
    .A2(net3795));
 sg13g2_a21oi_1 _19859_ (.A1(net2484),
    .A2(net4622),
    .Y(_05029_),
    .B1(_08484_));
 sg13g2_or4_1 _19860_ (.A(_05623_),
    .B(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .C(_06692_),
    .D(net4609),
    .X(_05030_));
 sg13g2_o21ai_1 _19861_ (.B1(_05030_),
    .Y(_05031_),
    .A1(_05009_),
    .A2(_05029_));
 sg13g2_nand3_1 _19862_ (.B(net3946),
    .C(_05031_),
    .A(net4710),
    .Y(_05032_));
 sg13g2_a22oi_1 _19863_ (.Y(_01956_),
    .B1(_05028_),
    .B2(_05032_),
    .A2(net3756),
    .A1(_05623_));
 sg13g2_nand2_1 _19864_ (.Y(_05033_),
    .A(_05691_),
    .B(net3752));
 sg13g2_o21ai_1 _19865_ (.B1(_05033_),
    .Y(_05034_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .A2(net3863));
 sg13g2_o21ai_1 _19866_ (.B1(_04995_),
    .Y(_05035_),
    .A1(net3789),
    .A2(_05034_));
 sg13g2_o21ai_1 _19867_ (.B1(_05035_),
    .Y(_05036_),
    .A1(net2559),
    .A2(net3792));
 sg13g2_or4_1 _19868_ (.A(_05624_),
    .B(net2201),
    .C(_06692_),
    .D(net4609),
    .X(_05037_));
 sg13g2_a21oi_1 _19869_ (.A1(net2559),
    .A2(net4622),
    .Y(_05038_),
    .B1(_08489_));
 sg13g2_o21ai_1 _19870_ (.B1(_05037_),
    .Y(_05039_),
    .A1(_05009_),
    .A2(_05038_));
 sg13g2_nand3_1 _19871_ (.B(net3946),
    .C(_05039_),
    .A(net4711),
    .Y(_05040_));
 sg13g2_a22oi_1 _19872_ (.Y(_01957_),
    .B1(_05036_),
    .B2(_05040_),
    .A2(net3756),
    .A1(_05624_));
 sg13g2_a221oi_1 _19873_ (.B2(_05692_),
    .C1(net3788),
    .B1(net3752),
    .A1(_05747_),
    .Y(_05041_),
    .A2(net3858));
 sg13g2_nand2_1 _19874_ (.Y(_05042_),
    .A(net4703),
    .B(_08493_));
 sg13g2_o21ai_1 _19875_ (.B1(_08495_),
    .Y(_05043_),
    .A1(net789),
    .A2(\soc_inst.cpu_core.mem_rs1_data[13] ));
 sg13g2_a21oi_1 _19876_ (.A1(_05042_),
    .A2(_05043_),
    .Y(_05044_),
    .B1(net3851));
 sg13g2_nor3_1 _19877_ (.A(net3755),
    .B(_05041_),
    .C(_05044_),
    .Y(_05045_));
 sg13g2_a21oi_1 _19878_ (.A1(_05626_),
    .A2(_04996_),
    .Y(_01958_),
    .B1(_05045_));
 sg13g2_a221oi_1 _19879_ (.B2(_05693_),
    .C1(net3788),
    .B1(net3752),
    .A1(_05748_),
    .Y(_05046_),
    .A2(net3858));
 sg13g2_nand2_1 _19880_ (.Y(_05047_),
    .A(net4703),
    .B(_08497_));
 sg13g2_o21ai_1 _19881_ (.B1(_08499_),
    .Y(_05048_),
    .A1(net1914),
    .A2(\soc_inst.cpu_core.mem_rs1_data[14] ));
 sg13g2_a21oi_1 _19882_ (.A1(_05047_),
    .A2(_05048_),
    .Y(_05049_),
    .B1(net3852));
 sg13g2_nor3_1 _19883_ (.A(net3756),
    .B(_05046_),
    .C(_05049_),
    .Y(_05050_));
 sg13g2_a21oi_1 _19884_ (.A1(_05627_),
    .A2(net3719),
    .Y(_01959_),
    .B1(_05050_));
 sg13g2_a221oi_1 _19885_ (.B2(_05694_),
    .C1(net3789),
    .B1(net3754),
    .A1(_05749_),
    .Y(_05051_),
    .A2(net3858));
 sg13g2_nand2_1 _19886_ (.Y(_05052_),
    .A(net4703),
    .B(_08501_));
 sg13g2_o21ai_1 _19887_ (.B1(_08503_),
    .Y(_05053_),
    .A1(net832),
    .A2(\soc_inst.cpu_core.mem_rs1_data[15] ));
 sg13g2_a21oi_1 _19888_ (.A1(_05052_),
    .A2(_05053_),
    .Y(_05054_),
    .B1(net3850));
 sg13g2_nor3_1 _19889_ (.A(net3755),
    .B(_05051_),
    .C(_05054_),
    .Y(_05055_));
 sg13g2_a21oi_1 _19890_ (.A1(_05629_),
    .A2(net3718),
    .Y(_01960_),
    .B1(_05055_));
 sg13g2_a221oi_1 _19891_ (.B2(_05696_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05750_),
    .Y(_05056_),
    .A2(net3857));
 sg13g2_nand2_1 _19892_ (.Y(_05057_),
    .A(net4706),
    .B(_08505_));
 sg13g2_o21ai_1 _19893_ (.B1(_08507_),
    .Y(_05058_),
    .A1(net2061),
    .A2(\soc_inst.cpu_core.mem_rs1_data[16] ));
 sg13g2_a21oi_1 _19894_ (.A1(_05057_),
    .A2(_05058_),
    .Y(_05059_),
    .B1(net3852));
 sg13g2_nor3_1 _19895_ (.A(net3756),
    .B(_05056_),
    .C(_05059_),
    .Y(_05060_));
 sg13g2_a21oi_1 _19896_ (.A1(_05631_),
    .A2(net3718),
    .Y(_01961_),
    .B1(_05060_));
 sg13g2_a221oi_1 _19897_ (.B2(_05697_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05751_),
    .Y(_05061_),
    .A2(net3857));
 sg13g2_nand2_1 _19898_ (.Y(_05062_),
    .A(net4706),
    .B(_08509_));
 sg13g2_o21ai_1 _19899_ (.B1(_08511_),
    .Y(_05063_),
    .A1(net2115),
    .A2(\soc_inst.cpu_core.mem_rs1_data[17] ));
 sg13g2_a21oi_1 _19900_ (.A1(_05062_),
    .A2(_05063_),
    .Y(_05064_),
    .B1(net3850));
 sg13g2_nor3_1 _19901_ (.A(net3756),
    .B(_05061_),
    .C(_05064_),
    .Y(_05065_));
 sg13g2_a21oi_1 _19902_ (.A1(_05633_),
    .A2(net3718),
    .Y(_01962_),
    .B1(_05065_));
 sg13g2_a221oi_1 _19903_ (.B2(_05698_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05752_),
    .Y(_05066_),
    .A2(net3857));
 sg13g2_nand2_1 _19904_ (.Y(_05067_),
    .A(net4703),
    .B(_08513_));
 sg13g2_o21ai_1 _19905_ (.B1(_08515_),
    .Y(_05068_),
    .A1(net1104),
    .A2(\soc_inst.cpu_core.mem_rs1_data[18] ));
 sg13g2_a21oi_1 _19906_ (.A1(_05067_),
    .A2(_05068_),
    .Y(_05069_),
    .B1(net3850));
 sg13g2_nor3_1 _19907_ (.A(net3755),
    .B(_05066_),
    .C(_05069_),
    .Y(_05070_));
 sg13g2_a21oi_1 _19908_ (.A1(_05635_),
    .A2(net3718),
    .Y(_01963_),
    .B1(_05070_));
 sg13g2_a221oi_1 _19909_ (.B2(_05699_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05753_),
    .Y(_05071_),
    .A2(net3857));
 sg13g2_nand2_1 _19910_ (.Y(_05072_),
    .A(net4703),
    .B(_08517_));
 sg13g2_o21ai_1 _19911_ (.B1(_08519_),
    .Y(_05073_),
    .A1(net1307),
    .A2(\soc_inst.cpu_core.mem_rs1_data[19] ));
 sg13g2_a21oi_1 _19912_ (.A1(_05072_),
    .A2(_05073_),
    .Y(_05074_),
    .B1(net3850));
 sg13g2_nor3_1 _19913_ (.A(net3755),
    .B(_05071_),
    .C(_05074_),
    .Y(_05075_));
 sg13g2_a21oi_1 _19914_ (.A1(_05637_),
    .A2(net3718),
    .Y(_01964_),
    .B1(_05075_));
 sg13g2_a221oi_1 _19915_ (.B2(_05700_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05754_),
    .Y(_05076_),
    .A2(net3857));
 sg13g2_nand2_1 _19916_ (.Y(_05077_),
    .A(net4706),
    .B(_08521_));
 sg13g2_o21ai_1 _19917_ (.B1(_08523_),
    .Y(_05078_),
    .A1(net1634),
    .A2(net1576));
 sg13g2_a21oi_1 _19918_ (.A1(_05077_),
    .A2(_05078_),
    .Y(_05079_),
    .B1(net3850));
 sg13g2_nor3_1 _19919_ (.A(net3756),
    .B(_05076_),
    .C(_05079_),
    .Y(_05080_));
 sg13g2_a21oi_1 _19920_ (.A1(_05639_),
    .A2(net3719),
    .Y(_01965_),
    .B1(_05080_));
 sg13g2_a221oi_1 _19921_ (.B2(_05702_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05755_),
    .Y(_05081_),
    .A2(net3857));
 sg13g2_nand2_1 _19922_ (.Y(_05082_),
    .A(net4703),
    .B(_08525_));
 sg13g2_o21ai_1 _19923_ (.B1(_08527_),
    .Y(_05083_),
    .A1(net1713),
    .A2(\soc_inst.cpu_core.mem_rs1_data[21] ));
 sg13g2_a21oi_1 _19924_ (.A1(_05082_),
    .A2(_05083_),
    .Y(_05084_),
    .B1(net3850));
 sg13g2_nor3_1 _19925_ (.A(net3755),
    .B(_05081_),
    .C(_05084_),
    .Y(_05085_));
 sg13g2_a21oi_1 _19926_ (.A1(_05641_),
    .A2(net3718),
    .Y(_01966_),
    .B1(_05085_));
 sg13g2_a221oi_1 _19927_ (.B2(_05703_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05756_),
    .Y(_05086_),
    .A2(net3857));
 sg13g2_nand2_1 _19928_ (.Y(_05087_),
    .A(net4703),
    .B(_08529_));
 sg13g2_o21ai_1 _19929_ (.B1(_08531_),
    .Y(_05088_),
    .A1(net925),
    .A2(\soc_inst.cpu_core.mem_rs1_data[22] ));
 sg13g2_a21oi_1 _19930_ (.A1(_05087_),
    .A2(_05088_),
    .Y(_05089_),
    .B1(net3850));
 sg13g2_nor3_1 _19931_ (.A(net3755),
    .B(_05086_),
    .C(_05089_),
    .Y(_05090_));
 sg13g2_a21oi_1 _19932_ (.A1(_05643_),
    .A2(net3718),
    .Y(_01967_),
    .B1(_05090_));
 sg13g2_a221oi_1 _19933_ (.B2(_05704_),
    .C1(net3787),
    .B1(net3751),
    .A1(_05757_),
    .Y(_05091_),
    .A2(net3857));
 sg13g2_nand2_1 _19934_ (.Y(_05092_),
    .A(net4703),
    .B(_08533_));
 sg13g2_o21ai_1 _19935_ (.B1(_08535_),
    .Y(_05093_),
    .A1(net1949),
    .A2(net2983));
 sg13g2_a21oi_1 _19936_ (.A1(_05092_),
    .A2(_05093_),
    .Y(_05094_),
    .B1(net3850));
 sg13g2_nor3_1 _19937_ (.A(net3755),
    .B(_05091_),
    .C(_05094_),
    .Y(_05095_));
 sg13g2_a21oi_1 _19938_ (.A1(_05645_),
    .A2(net3718),
    .Y(_01968_),
    .B1(_05095_));
 sg13g2_o21ai_1 _19939_ (.B1(net3860),
    .Y(_05096_),
    .A1(\soc_inst.cpu_core.id_int_is_interrupt ),
    .A2(\soc_inst.cpu_core.csr_file.mcause[31] ));
 sg13g2_a221oi_1 _19940_ (.B2(net2247),
    .C1(net3846),
    .B1(_08568_),
    .A1(net4879),
    .Y(_05097_),
    .A2(net4168));
 sg13g2_a21oi_1 _19941_ (.A1(net3846),
    .A2(_05096_),
    .Y(_05098_),
    .B1(_05097_));
 sg13g2_nand4_1 _19942_ (.B(_06731_),
    .C(_06797_),
    .A(net2247),
    .Y(_05099_),
    .D(_07217_));
 sg13g2_nand2b_1 _19943_ (.Y(_01969_),
    .B(net2248),
    .A_N(_05098_));
 sg13g2_nor2_1 _19944_ (.A(_06526_),
    .B(_07824_),
    .Y(_05100_));
 sg13g2_mux2_1 _19945_ (.A0(net2469),
    .A1(net5047),
    .S(_05100_),
    .X(_01970_));
 sg13g2_nor2_1 _19946_ (.A(_06526_),
    .B(_07120_),
    .Y(_05101_));
 sg13g2_mux2_1 _19947_ (.A0(net2488),
    .A1(net5047),
    .S(_05101_),
    .X(_01971_));
 sg13g2_o21ai_1 _19948_ (.B1(_07647_),
    .Y(_05102_),
    .A1(_06443_),
    .A2(_06980_));
 sg13g2_nand2_1 _19949_ (.Y(_05103_),
    .A(net90),
    .B(_05102_));
 sg13g2_o21ai_1 _19950_ (.B1(_07647_),
    .Y(_05104_),
    .A1(_05472_),
    .A2(net5128));
 sg13g2_o21ai_1 _19951_ (.B1(_05103_),
    .Y(_01972_),
    .A1(net280),
    .A2(_05104_));
 sg13g2_nor2b_1 _19952_ (.A(\soc_inst.gpio_inst.gpio_sync2[6] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[6] ),
    .Y(_05105_));
 sg13g2_a21oi_1 _19953_ (.A1(net80),
    .A2(_05105_),
    .Y(_05106_),
    .B1(net330));
 sg13g2_a21oi_1 _19954_ (.A1(net5031),
    .A2(_07131_),
    .Y(_01973_),
    .B1(net331));
 sg13g2_nor2b_1 _19955_ (.A(\soc_inst.gpio_inst.gpio_sync2[5] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[5] ),
    .Y(_05107_));
 sg13g2_a21oi_1 _19956_ (.A1(net88),
    .A2(_05107_),
    .Y(_05108_),
    .B1(net562));
 sg13g2_a21oi_1 _19957_ (.A1(net5034),
    .A2(_07131_),
    .Y(_01974_),
    .B1(net563));
 sg13g2_nor2b_1 _19958_ (.A(\soc_inst.gpio_inst.gpio_sync2[4] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[4] ),
    .Y(_05109_));
 sg13g2_a21oi_1 _19959_ (.A1(net83),
    .A2(_05109_),
    .Y(_05110_),
    .B1(net357));
 sg13g2_a21oi_1 _19960_ (.A1(net5037),
    .A2(_07131_),
    .Y(_01975_),
    .B1(net358));
 sg13g2_nor2b_1 _19961_ (.A(\soc_inst.gpio_inst.gpio_sync2[3] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[3] ),
    .Y(_05111_));
 sg13g2_a21oi_1 _19962_ (.A1(net86),
    .A2(_05111_),
    .Y(_05112_),
    .B1(net380));
 sg13g2_a21oi_1 _19963_ (.A1(net5039),
    .A2(_07131_),
    .Y(_01976_),
    .B1(net381));
 sg13g2_nor2b_1 _19964_ (.A(\soc_inst.gpio_inst.gpio_sync2[2] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[2] ),
    .Y(_05113_));
 sg13g2_a21oi_1 _19965_ (.A1(net84),
    .A2(_05113_),
    .Y(_05114_),
    .B1(net483));
 sg13g2_a21oi_1 _19966_ (.A1(net5043),
    .A2(_07131_),
    .Y(_01977_),
    .B1(net484));
 sg13g2_nor2b_1 _19967_ (.A(\soc_inst.gpio_inst.gpio_sync2[1] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[1] ),
    .Y(_05115_));
 sg13g2_a21oi_1 _19968_ (.A1(net82),
    .A2(_05115_),
    .Y(_05116_),
    .B1(net513));
 sg13g2_a21oi_1 _19969_ (.A1(net5045),
    .A2(_07131_),
    .Y(_01978_),
    .B1(net514));
 sg13g2_a21o_1 _19970_ (.A2(net2873),
    .A1(net4939),
    .B1(_02481_),
    .X(_01979_));
 sg13g2_a21o_1 _19971_ (.A2(net2838),
    .A1(net4971),
    .B1(_02483_),
    .X(_01980_));
 sg13g2_a21o_1 _19972_ (.A2(net2810),
    .A1(net4941),
    .B1(_02485_),
    .X(_01981_));
 sg13g2_a21o_1 _19973_ (.A2(net2878),
    .A1(net4970),
    .B1(_02487_),
    .X(_01982_));
 sg13g2_a21o_1 _19974_ (.A2(net2582),
    .A1(net4936),
    .B1(_02489_),
    .X(_01983_));
 sg13g2_a21o_1 _19975_ (.A2(net2805),
    .A1(net4941),
    .B1(_02491_),
    .X(_01984_));
 sg13g2_a21o_1 _19976_ (.A2(net2750),
    .A1(net4937),
    .B1(_02493_),
    .X(_01985_));
 sg13g2_a21o_1 _19977_ (.A2(net2910),
    .A1(net4970),
    .B1(_02495_),
    .X(_01986_));
 sg13g2_a21o_1 _19978_ (.A2(net2622),
    .A1(net4938),
    .B1(_02497_),
    .X(_01987_));
 sg13g2_a21o_1 _19979_ (.A2(net2763),
    .A1(net4938),
    .B1(_02499_),
    .X(_01988_));
 sg13g2_a21o_1 _19980_ (.A2(net2659),
    .A1(net4920),
    .B1(_02501_),
    .X(_01989_));
 sg13g2_a21o_1 _19981_ (.A2(net2660),
    .A1(net4920),
    .B1(_02503_),
    .X(_01990_));
 sg13g2_a21o_1 _19982_ (.A2(net2689),
    .A1(net4921),
    .B1(_02505_),
    .X(_01991_));
 sg13g2_a21o_1 _19983_ (.A2(net2806),
    .A1(net4925),
    .B1(_02507_),
    .X(_01992_));
 sg13g2_a21o_1 _19984_ (.A2(net2668),
    .A1(net4918),
    .B1(_02509_),
    .X(_01993_));
 sg13g2_a21o_1 _19985_ (.A2(net2790),
    .A1(net4918),
    .B1(_02511_),
    .X(_01994_));
 sg13g2_a21o_1 _19986_ (.A2(net2830),
    .A1(net4952),
    .B1(_02513_),
    .X(_01995_));
 sg13g2_a21o_1 _19987_ (.A2(net2772),
    .A1(net4910),
    .B1(_02515_),
    .X(_01996_));
 sg13g2_a21o_1 _19988_ (.A2(net2671),
    .A1(net4911),
    .B1(_02517_),
    .X(_01997_));
 sg13g2_a21o_1 _19989_ (.A2(net2628),
    .A1(net4910),
    .B1(_02519_),
    .X(_01998_));
 sg13g2_a21o_1 _19990_ (.A2(net2757),
    .A1(net4911),
    .B1(_02521_),
    .X(_01999_));
 sg13g2_a21o_1 _19991_ (.A2(net2765),
    .A1(net4911),
    .B1(_02523_),
    .X(_02000_));
 sg13g2_a21o_1 _19992_ (.A2(net2872),
    .A1(net4900),
    .B1(_02525_),
    .X(_02001_));
 sg13g2_a21o_1 _19993_ (.A2(net2560),
    .A1(net4900),
    .B1(_02527_),
    .X(_02002_));
 sg13g2_nand2_1 _19994_ (.Y(_05117_),
    .A(net4785),
    .B(_07861_));
 sg13g2_nor2_1 _19995_ (.A(_06296_),
    .B(_05117_),
    .Y(_05118_));
 sg13g2_nor2_1 _19996_ (.A(net1718),
    .B(net3968),
    .Y(_05119_));
 sg13g2_a21oi_1 _19997_ (.A1(net5049),
    .A2(net3968),
    .Y(_02003_),
    .B1(_05119_));
 sg13g2_nor2_1 _19998_ (.A(net1917),
    .B(net3968),
    .Y(_05120_));
 sg13g2_a21oi_1 _19999_ (.A1(net5044),
    .A2(net3967),
    .Y(_02004_),
    .B1(_05120_));
 sg13g2_nor2_1 _20000_ (.A(net1621),
    .B(net3967),
    .Y(_05121_));
 sg13g2_a21oi_1 _20001_ (.A1(net5043),
    .A2(net3967),
    .Y(_02005_),
    .B1(_05121_));
 sg13g2_nor2_1 _20002_ (.A(net1304),
    .B(net3969),
    .Y(_05122_));
 sg13g2_a21oi_1 _20003_ (.A1(net5040),
    .A2(net3967),
    .Y(_02006_),
    .B1(_05122_));
 sg13g2_nor2_1 _20004_ (.A(net1464),
    .B(net3968),
    .Y(_05123_));
 sg13g2_a21oi_1 _20005_ (.A1(net5037),
    .A2(net3968),
    .Y(_02007_),
    .B1(_05123_));
 sg13g2_nor2_1 _20006_ (.A(net1838),
    .B(net3969),
    .Y(_05124_));
 sg13g2_a21oi_1 _20007_ (.A1(net5034),
    .A2(net3969),
    .Y(_02008_),
    .B1(_05124_));
 sg13g2_nor2_1 _20008_ (.A(net1425),
    .B(net3968),
    .Y(_05125_));
 sg13g2_a21oi_1 _20009_ (.A1(net5031),
    .A2(net3969),
    .Y(_02009_),
    .B1(_05125_));
 sg13g2_nor2_1 _20010_ (.A(net1964),
    .B(net3968),
    .Y(_05126_));
 sg13g2_a21oi_1 _20011_ (.A1(net5028),
    .A2(net3968),
    .Y(_02010_),
    .B1(_05126_));
 sg13g2_nor2_1 _20012_ (.A(net1517),
    .B(net3967),
    .Y(_05127_));
 sg13g2_a21oi_1 _20013_ (.A1(net5026),
    .A2(net3967),
    .Y(_02011_),
    .B1(_05127_));
 sg13g2_nor2_1 _20014_ (.A(net1767),
    .B(net3967),
    .Y(_05128_));
 sg13g2_a21oi_1 _20015_ (.A1(net5024),
    .A2(net3967),
    .Y(_02012_),
    .B1(_05128_));
 sg13g2_nor2_1 _20016_ (.A(net1421),
    .B(net3966),
    .Y(_05129_));
 sg13g2_a21oi_1 _20017_ (.A1(net5023),
    .A2(net3966),
    .Y(_02013_),
    .B1(_05129_));
 sg13g2_nor2_1 _20018_ (.A(net1416),
    .B(net3965),
    .Y(_05130_));
 sg13g2_a21oi_1 _20019_ (.A1(net5022),
    .A2(net3965),
    .Y(_02014_),
    .B1(_05130_));
 sg13g2_nor2_1 _20020_ (.A(net1383),
    .B(net3965),
    .Y(_05131_));
 sg13g2_a21oi_1 _20021_ (.A1(net5021),
    .A2(net3965),
    .Y(_02015_),
    .B1(_05131_));
 sg13g2_nor2_1 _20022_ (.A(net1786),
    .B(net3965),
    .Y(_05132_));
 sg13g2_a21oi_1 _20023_ (.A1(net5020),
    .A2(net3965),
    .Y(_02016_),
    .B1(_05132_));
 sg13g2_nor2_1 _20024_ (.A(net2116),
    .B(net3965),
    .Y(_05133_));
 sg13g2_a21oi_1 _20025_ (.A1(net5019),
    .A2(net3965),
    .Y(_02017_),
    .B1(_05133_));
 sg13g2_nor2_1 _20026_ (.A(net1758),
    .B(net3966),
    .Y(_05134_));
 sg13g2_a21oi_1 _20027_ (.A1(net5018),
    .A2(net3966),
    .Y(_02018_),
    .B1(_05134_));
 sg13g2_nor3_1 _20028_ (.A(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .B(net3800),
    .C(_06733_),
    .Y(_05135_));
 sg13g2_a221oi_1 _20029_ (.B2(net2084),
    .C1(net3855),
    .B1(_08476_),
    .A1(net457),
    .Y(_05136_),
    .A2(net4172));
 sg13g2_nor4_1 _20030_ (.A(net5054),
    .B(net2084),
    .C(net3796),
    .D(_06733_),
    .Y(_05137_));
 sg13g2_nor3_1 _20031_ (.A(_05135_),
    .B(_05136_),
    .C(_05137_),
    .Y(_05138_));
 sg13g2_nor2_1 _20032_ (.A(_06672_),
    .B(_04799_),
    .Y(_05139_));
 sg13g2_a21o_1 _20033_ (.A2(_05139_),
    .A1(net2084),
    .B1(_05138_),
    .X(_02019_));
 sg13g2_o21ai_1 _20034_ (.B1(_06734_),
    .Y(_05140_),
    .A1(net2382),
    .A2(net5054));
 sg13g2_a22oi_1 _20035_ (.Y(_05141_),
    .B1(_08487_),
    .B2(_05398_),
    .A2(net4171),
    .A1(\soc_inst.cpu_core.mem_rs1_data[11] ));
 sg13g2_nand2b_1 _20036_ (.Y(_05142_),
    .B(_05141_),
    .A_N(net3855));
 sg13g2_a22oi_1 _20037_ (.Y(_02020_),
    .B1(_05140_),
    .B2(_05142_),
    .A2(_05139_),
    .A1(_05398_));
 sg13g2_o21ai_1 _20038_ (.B1(_06734_),
    .Y(_05143_),
    .A1(net2074),
    .A2(net5056));
 sg13g2_a22oi_1 _20039_ (.Y(_05144_),
    .B1(_08491_),
    .B2(_05397_),
    .A2(net4171),
    .A1(\soc_inst.cpu_core.mem_rs1_data[12] ));
 sg13g2_nand2b_1 _20040_ (.Y(_05145_),
    .B(_05144_),
    .A_N(net3855));
 sg13g2_a22oi_1 _20041_ (.Y(_02021_),
    .B1(_05143_),
    .B2(_05145_),
    .A2(_05139_),
    .A1(_05397_));
 sg13g2_nand2_1 _20042_ (.Y(_05146_),
    .A(net5060),
    .B(_09010_));
 sg13g2_nor2_2 _20043_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ),
    .B(_05146_),
    .Y(_05147_));
 sg13g2_nor2_1 _20044_ (.A(net4597),
    .B(net2739),
    .Y(_05148_));
 sg13g2_o21ai_1 _20045_ (.B1(net4596),
    .Y(_05149_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ),
    .A2(_05146_));
 sg13g2_and2_1 _20046_ (.A(net2240),
    .B(net4596),
    .X(_05150_));
 sg13g2_a21oi_1 _20047_ (.A1(net1712),
    .A2(net4597),
    .Y(_05151_),
    .B1(_05150_));
 sg13g2_o21ai_1 _20048_ (.B1(net5481),
    .Y(_05152_),
    .A1(net2405),
    .A2(net3964));
 sg13g2_a21oi_1 _20049_ (.A1(net3964),
    .A2(_05151_),
    .Y(_02022_),
    .B1(_05152_));
 sg13g2_and2_1 _20050_ (.A(net1979),
    .B(net4596),
    .X(_05153_));
 sg13g2_a21oi_1 _20051_ (.A1(net1156),
    .A2(net4597),
    .Y(_05154_),
    .B1(_05153_));
 sg13g2_o21ai_1 _20052_ (.B1(net5481),
    .Y(_05155_),
    .A1(net2240),
    .A2(net3964));
 sg13g2_a21oi_1 _20053_ (.A1(net3964),
    .A2(_05154_),
    .Y(_02023_),
    .B1(_05155_));
 sg13g2_and2_1 _20054_ (.A(net1962),
    .B(net4596),
    .X(_05156_));
 sg13g2_a21oi_1 _20055_ (.A1(net990),
    .A2(net4597),
    .Y(_05157_),
    .B1(_05156_));
 sg13g2_o21ai_1 _20056_ (.B1(net5481),
    .Y(_05158_),
    .A1(net1979),
    .A2(net3964));
 sg13g2_a21oi_1 _20057_ (.A1(net3964),
    .A2(_05157_),
    .Y(_02024_),
    .B1(_05158_));
 sg13g2_and2_1 _20058_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ),
    .B(net4596),
    .X(_05159_));
 sg13g2_a21oi_1 _20059_ (.A1(net1359),
    .A2(net4597),
    .Y(_05160_),
    .B1(_05159_));
 sg13g2_o21ai_1 _20060_ (.B1(net5482),
    .Y(_05161_),
    .A1(net1962),
    .A2(net3964));
 sg13g2_a21oi_1 _20061_ (.A1(net3964),
    .A2(_05160_),
    .Y(_02025_),
    .B1(_05161_));
 sg13g2_nand2_1 _20062_ (.Y(_05162_),
    .A(net374),
    .B(net4596));
 sg13g2_a21oi_1 _20063_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ),
    .A2(net4597),
    .Y(_05163_),
    .B1(_05148_));
 sg13g2_o21ai_1 _20064_ (.B1(net5482),
    .Y(_05164_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ),
    .A2(_05149_));
 sg13g2_a21oi_1 _20065_ (.A1(net375),
    .A2(_05163_),
    .Y(_02026_),
    .B1(_05164_));
 sg13g2_nor2_1 _20066_ (.A(net2739),
    .B(_05162_),
    .Y(_05165_));
 sg13g2_a21oi_1 _20067_ (.A1(net1154),
    .A2(net4597),
    .Y(_05166_),
    .B1(_05165_));
 sg13g2_nand2_1 _20068_ (.Y(_05167_),
    .A(net2528),
    .B(net4596));
 sg13g2_o21ai_1 _20069_ (.B1(_05166_),
    .Y(_05168_),
    .A1(_05148_),
    .A2(_05167_));
 sg13g2_and2_1 _20070_ (.A(net5482),
    .B(_05168_),
    .X(_02027_));
 sg13g2_nor2_1 _20071_ (.A(_05147_),
    .B(_05167_),
    .Y(_05169_));
 sg13g2_and2_1 _20072_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[7] ),
    .B(_08991_),
    .X(_05170_));
 sg13g2_a221oi_1 _20073_ (.B2(_05170_),
    .C1(net2529),
    .B1(_05147_),
    .A1(net842),
    .Y(_05171_),
    .A2(net4597));
 sg13g2_nor2b_1 _20074_ (.A(net2530),
    .B_N(net5482),
    .Y(_02028_));
 sg13g2_mux2_1 _20075_ (.A0(net5044),
    .A1(net1532),
    .S(_07013_),
    .X(_02029_));
 sg13g2_nor2_2 _20076_ (.A(net4268),
    .B(_05117_),
    .Y(_05172_));
 sg13g2_nor2_1 _20077_ (.A(net1033),
    .B(net3958),
    .Y(_05173_));
 sg13g2_a21oi_1 _20078_ (.A1(net5047),
    .A2(net3958),
    .Y(_02030_),
    .B1(_05173_));
 sg13g2_nor2_1 _20079_ (.A(net1182),
    .B(net3962),
    .Y(_05174_));
 sg13g2_a21oi_1 _20080_ (.A1(net5044),
    .A2(net3962),
    .Y(_02031_),
    .B1(_05174_));
 sg13g2_nor2_1 _20081_ (.A(net1480),
    .B(net3962),
    .Y(_05175_));
 sg13g2_a21oi_1 _20082_ (.A1(net5041),
    .A2(net3958),
    .Y(_02032_),
    .B1(_05175_));
 sg13g2_nor2_1 _20083_ (.A(net1492),
    .B(net3962),
    .Y(_05176_));
 sg13g2_a21oi_1 _20084_ (.A1(net5038),
    .A2(net3962),
    .Y(_02033_),
    .B1(_05176_));
 sg13g2_nor2_1 _20085_ (.A(net1234),
    .B(net3962),
    .Y(_05177_));
 sg13g2_a21oi_1 _20086_ (.A1(net5035),
    .A2(net3962),
    .Y(_02034_),
    .B1(_05177_));
 sg13g2_nor2_1 _20087_ (.A(net1347),
    .B(net3962),
    .Y(_05178_));
 sg13g2_a21oi_1 _20088_ (.A1(net5033),
    .A2(net3963),
    .Y(_02035_),
    .B1(_05178_));
 sg13g2_nor2_1 _20089_ (.A(net1814),
    .B(net3963),
    .Y(_05179_));
 sg13g2_a21oi_1 _20090_ (.A1(net5032),
    .A2(net3963),
    .Y(_02036_),
    .B1(_05179_));
 sg13g2_nor2_1 _20091_ (.A(net1861),
    .B(net3961),
    .Y(_05180_));
 sg13g2_a21oi_1 _20092_ (.A1(net5028),
    .A2(net3961),
    .Y(_02037_),
    .B1(_05180_));
 sg13g2_nor2_1 _20093_ (.A(net1487),
    .B(net3957),
    .Y(_05181_));
 sg13g2_a21oi_1 _20094_ (.A1(net5026),
    .A2(net3957),
    .Y(_02038_),
    .B1(_05181_));
 sg13g2_nor2_1 _20095_ (.A(net1187),
    .B(net3957),
    .Y(_05182_));
 sg13g2_a21oi_1 _20096_ (.A1(net5024),
    .A2(net3957),
    .Y(_02039_),
    .B1(_05182_));
 sg13g2_nor2_1 _20097_ (.A(net1608),
    .B(net3958),
    .Y(_05183_));
 sg13g2_a21oi_1 _20098_ (.A1(net5023),
    .A2(net3958),
    .Y(_02040_),
    .B1(_05183_));
 sg13g2_nor2_1 _20099_ (.A(net1686),
    .B(net3958),
    .Y(_05184_));
 sg13g2_a21oi_1 _20100_ (.A1(net5022),
    .A2(net3955),
    .Y(_02041_),
    .B1(_05184_));
 sg13g2_nor2_1 _20101_ (.A(net1361),
    .B(net3954),
    .Y(_05185_));
 sg13g2_a21oi_1 _20102_ (.A1(\soc_inst.core_mem_wdata[12] ),
    .A2(net3954),
    .Y(_02042_),
    .B1(_05185_));
 sg13g2_nor2_1 _20103_ (.A(net2008),
    .B(net3958),
    .Y(_05186_));
 sg13g2_a21oi_1 _20104_ (.A1(net5020),
    .A2(net3954),
    .Y(_02043_),
    .B1(_05186_));
 sg13g2_nor2_1 _20105_ (.A(net1132),
    .B(net3954),
    .Y(_05187_));
 sg13g2_a21oi_1 _20106_ (.A1(net5019),
    .A2(net3955),
    .Y(_02044_),
    .B1(_05187_));
 sg13g2_nor2_1 _20107_ (.A(net1455),
    .B(net3955),
    .Y(_05188_));
 sg13g2_a21oi_1 _20108_ (.A1(net770),
    .A2(net3955),
    .Y(_02045_),
    .B1(_05188_));
 sg13g2_nor2_1 _20109_ (.A(net1217),
    .B(net3953),
    .Y(_05189_));
 sg13g2_a21oi_1 _20110_ (.A1(\soc_inst.core_mem_wdata[16] ),
    .A2(net3953),
    .Y(_02046_),
    .B1(_05189_));
 sg13g2_nor2_1 _20111_ (.A(net1739),
    .B(net3953),
    .Y(_05190_));
 sg13g2_a21oi_1 _20112_ (.A1(\soc_inst.core_mem_wdata[17] ),
    .A2(net3953),
    .Y(_02047_),
    .B1(_05190_));
 sg13g2_nor2_1 _20113_ (.A(net1596),
    .B(net3954),
    .Y(_05191_));
 sg13g2_a21oi_1 _20114_ (.A1(net1170),
    .A2(net3953),
    .Y(_02048_),
    .B1(_05191_));
 sg13g2_nor2_1 _20115_ (.A(_00314_),
    .B(net3956),
    .Y(_05192_));
 sg13g2_a21oi_1 _20116_ (.A1(net1021),
    .A2(net3956),
    .Y(_02049_),
    .B1(_05192_));
 sg13g2_nor2_1 _20117_ (.A(net1496),
    .B(net3954),
    .Y(_05193_));
 sg13g2_a21oi_1 _20118_ (.A1(\soc_inst.core_mem_wdata[20] ),
    .A2(net3953),
    .Y(_02050_),
    .B1(_05193_));
 sg13g2_nor2_1 _20119_ (.A(net1925),
    .B(net3954),
    .Y(_05194_));
 sg13g2_a21oi_1 _20120_ (.A1(\soc_inst.core_mem_wdata[21] ),
    .A2(net3954),
    .Y(_02051_),
    .B1(_05194_));
 sg13g2_nor2_1 _20121_ (.A(net1389),
    .B(net3957),
    .Y(_05195_));
 sg13g2_a21oi_1 _20122_ (.A1(\soc_inst.core_mem_wdata[22] ),
    .A2(net3957),
    .Y(_02052_),
    .B1(_05195_));
 sg13g2_nor2_1 _20123_ (.A(net1856),
    .B(net3953),
    .Y(_05196_));
 sg13g2_a21oi_1 _20124_ (.A1(\soc_inst.core_mem_wdata[23] ),
    .A2(net3953),
    .Y(_02053_),
    .B1(_05196_));
 sg13g2_nor2_1 _20125_ (.A(net2221),
    .B(net3960),
    .Y(_05197_));
 sg13g2_a21oi_1 _20126_ (.A1(net962),
    .A2(net3960),
    .Y(_02054_),
    .B1(_05197_));
 sg13g2_nor2_1 _20127_ (.A(net2304),
    .B(net3960),
    .Y(_05198_));
 sg13g2_a21oi_1 _20128_ (.A1(\soc_inst.core_mem_wdata[25] ),
    .A2(net3960),
    .Y(_02055_),
    .B1(_05198_));
 sg13g2_nor2_1 _20129_ (.A(_00321_),
    .B(net3959),
    .Y(_05199_));
 sg13g2_a21oi_1 _20130_ (.A1(net532),
    .A2(net3960),
    .Y(_02056_),
    .B1(_05199_));
 sg13g2_nor2_1 _20131_ (.A(_00322_),
    .B(net3959),
    .Y(_05200_));
 sg13g2_a21oi_1 _20132_ (.A1(net480),
    .A2(net3960),
    .Y(_02057_),
    .B1(_05200_));
 sg13g2_nor2_1 _20133_ (.A(_00323_),
    .B(net3959),
    .Y(_05201_));
 sg13g2_a21oi_1 _20134_ (.A1(net610),
    .A2(net3960),
    .Y(_02058_),
    .B1(_05201_));
 sg13g2_nor2_1 _20135_ (.A(net2311),
    .B(net3961),
    .Y(_05202_));
 sg13g2_a21oi_1 _20136_ (.A1(\soc_inst.core_mem_wdata[29] ),
    .A2(net3959),
    .Y(_02059_),
    .B1(_05202_));
 sg13g2_nor2_1 _20137_ (.A(_00325_),
    .B(net3959),
    .Y(_05203_));
 sg13g2_a21oi_1 _20138_ (.A1(net383),
    .A2(net3959),
    .Y(_02060_),
    .B1(_05203_));
 sg13g2_nor2_1 _20139_ (.A(_00326_),
    .B(net3959),
    .Y(_05204_));
 sg13g2_a21oi_1 _20140_ (.A1(net422),
    .A2(net3959),
    .Y(_02061_),
    .B1(_05204_));
 sg13g2_nor2_2 _20141_ (.A(_07011_),
    .B(_07120_),
    .Y(_05205_));
 sg13g2_mux2_1 _20142_ (.A0(net1712),
    .A1(net5048),
    .S(_05205_),
    .X(_02062_));
 sg13g2_mux2_1 _20143_ (.A0(net1156),
    .A1(net5045),
    .S(_05205_),
    .X(_02063_));
 sg13g2_mux2_1 _20144_ (.A0(net990),
    .A1(net5042),
    .S(_05205_),
    .X(_02064_));
 sg13g2_mux2_1 _20145_ (.A0(net1359),
    .A1(net5039),
    .S(_05205_),
    .X(_02065_));
 sg13g2_mux2_1 _20146_ (.A0(net1483),
    .A1(net5035),
    .S(_05205_),
    .X(_02066_));
 sg13g2_mux2_1 _20147_ (.A0(net1154),
    .A1(net5033),
    .S(_05205_),
    .X(_02067_));
 sg13g2_mux2_1 _20148_ (.A0(net842),
    .A1(net5031),
    .S(_05205_),
    .X(_02068_));
 sg13g2_mux2_1 _20149_ (.A0(net572),
    .A1(net5029),
    .S(_05205_),
    .X(_02069_));
 sg13g2_a21oi_1 _20150_ (.A1(net572),
    .A2(_08990_),
    .Y(_05206_),
    .B1(_05170_));
 sg13g2_nor2b_1 _20151_ (.A(net573),
    .B_N(net5483),
    .Y(_02070_));
 sg13g2_a21oi_1 _20152_ (.A1(net5060),
    .A2(_09010_),
    .Y(_05207_),
    .B1(net517));
 sg13g2_nand4_1 _20153_ (.B(_05393_),
    .C(_05410_),
    .A(net869),
    .Y(_05208_),
    .D(_08987_));
 sg13g2_nand3_1 _20154_ (.B(net5480),
    .C(_05208_),
    .A(net5060),
    .Y(_05209_));
 sg13g2_nor2_1 _20155_ (.A(_05393_),
    .B(_05146_),
    .Y(_05210_));
 sg13g2_nor3_1 _20156_ (.A(net518),
    .B(_05209_),
    .C(_05210_),
    .Y(_02071_));
 sg13g2_nor2_1 _20157_ (.A(net1801),
    .B(_05210_),
    .Y(_05211_));
 sg13g2_and2_1 _20158_ (.A(net1801),
    .B(_05210_),
    .X(_05212_));
 sg13g2_nor3_1 _20159_ (.A(_05209_),
    .B(_05211_),
    .C(_05212_),
    .Y(_02072_));
 sg13g2_xnor2_1 _20160_ (.Y(_05213_),
    .A(net2059),
    .B(_05212_));
 sg13g2_nor2_1 _20161_ (.A(_05209_),
    .B(_05213_),
    .Y(_02073_));
 sg13g2_a21oi_1 _20162_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ),
    .A2(_05212_),
    .Y(_05214_),
    .B1(net869));
 sg13g2_and3_1 _20163_ (.X(_05215_),
    .A(net869),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ),
    .C(_05212_));
 sg13g2_nor3_1 _20164_ (.A(_05209_),
    .B(net870),
    .C(_05215_),
    .Y(_02074_));
 sg13g2_nor3_1 _20165_ (.A(net2892),
    .B(net2738),
    .C(net5060),
    .Y(_05216_));
 sg13g2_nor2_1 _20166_ (.A(_05392_),
    .B(_07850_),
    .Y(_05217_));
 sg13g2_nor3_1 _20167_ (.A(_09011_),
    .B(_05216_),
    .C(_05217_),
    .Y(_02075_));
 sg13g2_and2_1 _20168_ (.A(net1840),
    .B(_05217_),
    .X(_05218_));
 sg13g2_nor2_1 _20169_ (.A(net1840),
    .B(_05217_),
    .Y(_05219_));
 sg13g2_nor3_1 _20170_ (.A(_09011_),
    .B(_05218_),
    .C(net1841),
    .Y(_02076_));
 sg13g2_and2_1 _20171_ (.A(net1448),
    .B(_05218_),
    .X(_05220_));
 sg13g2_nor2_1 _20172_ (.A(net1448),
    .B(_05218_),
    .Y(_05221_));
 sg13g2_nor3_1 _20173_ (.A(net4023),
    .B(_05220_),
    .C(net1449),
    .Y(_02077_));
 sg13g2_and2_1 _20174_ (.A(net1842),
    .B(_05220_),
    .X(_05222_));
 sg13g2_nor2_1 _20175_ (.A(net1842),
    .B(_05220_),
    .Y(_05223_));
 sg13g2_nor3_1 _20176_ (.A(net4023),
    .B(_05222_),
    .C(_05223_),
    .Y(_02078_));
 sg13g2_and2_1 _20177_ (.A(net1364),
    .B(_05222_),
    .X(_05224_));
 sg13g2_nor2_1 _20178_ (.A(net1364),
    .B(_05222_),
    .Y(_05225_));
 sg13g2_nor3_1 _20179_ (.A(net4023),
    .B(_05224_),
    .C(net1365),
    .Y(_02079_));
 sg13g2_xnor2_1 _20180_ (.Y(_05226_),
    .A(net2199),
    .B(_05224_));
 sg13g2_nor2_1 _20181_ (.A(net4023),
    .B(_05226_),
    .Y(_02080_));
 sg13g2_a21oi_1 _20182_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .A2(_05224_),
    .Y(_05227_),
    .B1(net1311));
 sg13g2_and3_1 _20183_ (.X(_05228_),
    .A(net1311),
    .B(net2981),
    .C(_05224_));
 sg13g2_nor3_1 _20184_ (.A(net4023),
    .B(net1312),
    .C(_05228_),
    .Y(_02081_));
 sg13g2_nor2_1 _20185_ (.A(net2142),
    .B(_05228_),
    .Y(_05229_));
 sg13g2_and2_1 _20186_ (.A(net2142),
    .B(_05228_),
    .X(_05230_));
 sg13g2_nor3_1 _20187_ (.A(net4023),
    .B(net2143),
    .C(_05230_),
    .Y(_02082_));
 sg13g2_nor2_1 _20188_ (.A(net2167),
    .B(_05230_),
    .Y(_05231_));
 sg13g2_and2_1 _20189_ (.A(net2167),
    .B(_05230_),
    .X(_05232_));
 sg13g2_nor3_1 _20190_ (.A(net4023),
    .B(net2168),
    .C(_05232_),
    .Y(_02083_));
 sg13g2_a21oi_1 _20191_ (.A1(net2500),
    .A2(_05232_),
    .Y(_05233_),
    .B1(net4023));
 sg13g2_o21ai_1 _20192_ (.B1(_05233_),
    .Y(_05234_),
    .A1(net2500),
    .A2(_05232_));
 sg13g2_inv_1 _20193_ (.Y(_02084_),
    .A(_05234_));
 sg13g2_nor2_1 _20194_ (.A(_07011_),
    .B(_07824_),
    .Y(_05235_));
 sg13g2_mux2_1 _20195_ (.A0(net2525),
    .A1(net5048),
    .S(net3951),
    .X(_02085_));
 sg13g2_nand2_1 _20196_ (.Y(_05236_),
    .A(net5044),
    .B(net3951));
 sg13g2_o21ai_1 _20197_ (.B1(_05236_),
    .Y(_02086_),
    .A1(_05412_),
    .A2(net3950));
 sg13g2_nor2_1 _20198_ (.A(net2652),
    .B(net3950),
    .Y(_05237_));
 sg13g2_a21oi_1 _20199_ (.A1(net5041),
    .A2(net3950),
    .Y(_02087_),
    .B1(_05237_));
 sg13g2_nor2_1 _20200_ (.A(net2766),
    .B(net3950),
    .Y(_05238_));
 sg13g2_a21oi_1 _20201_ (.A1(net5038),
    .A2(net3950),
    .Y(_02088_),
    .B1(_05238_));
 sg13g2_mux2_1 _20202_ (.A0(net2839),
    .A1(net5035),
    .S(net3950),
    .X(_02089_));
 sg13g2_nor2_1 _20203_ (.A(net2654),
    .B(net3950),
    .Y(_05239_));
 sg13g2_a21oi_1 _20204_ (.A1(net5033),
    .A2(net3950),
    .Y(_02090_),
    .B1(_05239_));
 sg13g2_mux2_1 _20205_ (.A0(net2103),
    .A1(net5032),
    .S(net3951),
    .X(_02091_));
 sg13g2_mux2_1 _20206_ (.A0(net2803),
    .A1(net5029),
    .S(net3951),
    .X(_02092_));
 sg13g2_mux2_1 _20207_ (.A0(net2894),
    .A1(net5026),
    .S(net3952),
    .X(_02093_));
 sg13g2_nor2_1 _20208_ (.A(net4758),
    .B(net3952),
    .Y(_05240_));
 sg13g2_a21oi_1 _20209_ (.A1(net5024),
    .A2(net3952),
    .Y(_02094_),
    .B1(_05240_));
 sg13g2_o21ai_1 _20210_ (.B1(_08995_),
    .Y(_05241_),
    .A1(net2405),
    .A2(_09012_));
 sg13g2_nand2_1 _20211_ (.Y(_02095_),
    .A(net5482),
    .B(_05241_));
 sg13g2_o21ai_1 _20212_ (.B1(net4700),
    .Y(_05242_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .A2(net4609));
 sg13g2_nand3_1 _20213_ (.B(net4251),
    .C(_05242_),
    .A(net2414),
    .Y(_05243_));
 sg13g2_o21ai_1 _20214_ (.B1(net4618),
    .Y(_05244_),
    .A1(net2414),
    .A2(net928));
 sg13g2_nand3_1 _20215_ (.B(_05243_),
    .C(_05244_),
    .A(_05042_),
    .Y(_05245_));
 sg13g2_mux2_1 _20216_ (.A0(_05245_),
    .A1(net2414),
    .S(net3855),
    .X(_02096_));
 sg13g2_o21ai_1 _20217_ (.B1(net4699),
    .Y(_05246_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .A2(net4610));
 sg13g2_nand3_1 _20218_ (.B(net4257),
    .C(_05246_),
    .A(net2047),
    .Y(_05247_));
 sg13g2_o21ai_1 _20219_ (.B1(net4621),
    .Y(_05248_),
    .A1(net2047),
    .A2(\soc_inst.cpu_core.mem_rs1_data[14] ));
 sg13g2_nand3_1 _20220_ (.B(_05247_),
    .C(_05248_),
    .A(_05047_),
    .Y(_05249_));
 sg13g2_mux2_1 _20221_ (.A0(_05249_),
    .A1(net2047),
    .S(net3856),
    .X(_02097_));
 sg13g2_o21ai_1 _20222_ (.B1(net4700),
    .Y(_05250_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .A2(net4608));
 sg13g2_nand3_1 _20223_ (.B(net4251),
    .C(_05250_),
    .A(net2370),
    .Y(_05251_));
 sg13g2_o21ai_1 _20224_ (.B1(net4618),
    .Y(_05252_),
    .A1(net2370),
    .A2(net932));
 sg13g2_nand3_1 _20225_ (.B(_05251_),
    .C(_05252_),
    .A(_05052_),
    .Y(_05253_));
 sg13g2_mux2_1 _20226_ (.A0(_05253_),
    .A1(net2370),
    .S(net3854),
    .X(_02098_));
 sg13g2_o21ai_1 _20227_ (.B1(net4698),
    .Y(_05254_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .A2(net4606));
 sg13g2_nand3_1 _20228_ (.B(net4252),
    .C(_05254_),
    .A(net2099),
    .Y(_05255_));
 sg13g2_o21ai_1 _20229_ (.B1(net4617),
    .Y(_05256_),
    .A1(net2099),
    .A2(\soc_inst.cpu_core.mem_rs1_data[16] ));
 sg13g2_nand3_1 _20230_ (.B(_05255_),
    .C(_05256_),
    .A(_05057_),
    .Y(_05257_));
 sg13g2_mux2_1 _20231_ (.A0(_05257_),
    .A1(net2099),
    .S(net3853),
    .X(_02099_));
 sg13g2_o21ai_1 _20232_ (.B1(net4698),
    .Y(_05258_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .A2(net4605));
 sg13g2_nand3_1 _20233_ (.B(net4252),
    .C(_05258_),
    .A(net2002),
    .Y(_05259_));
 sg13g2_o21ai_1 _20234_ (.B1(net4617),
    .Y(_05260_),
    .A1(net2002),
    .A2(\soc_inst.cpu_core.mem_rs1_data[17] ));
 sg13g2_nand3_1 _20235_ (.B(_05259_),
    .C(_05260_),
    .A(_05062_),
    .Y(_05261_));
 sg13g2_mux2_1 _20236_ (.A0(_05261_),
    .A1(net2002),
    .S(net3853),
    .X(_02100_));
 sg13g2_o21ai_1 _20237_ (.B1(net4700),
    .Y(_05262_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .A2(net4603));
 sg13g2_nand3_1 _20238_ (.B(net4249),
    .C(_05262_),
    .A(net2070),
    .Y(_05263_));
 sg13g2_o21ai_1 _20239_ (.B1(net4618),
    .Y(_05264_),
    .A1(net2070),
    .A2(\soc_inst.cpu_core.mem_rs1_data[18] ));
 sg13g2_nand3_1 _20240_ (.B(_05263_),
    .C(_05264_),
    .A(_05067_),
    .Y(_05265_));
 sg13g2_mux2_1 _20241_ (.A0(_05265_),
    .A1(net2070),
    .S(net3854),
    .X(_02101_));
 sg13g2_o21ai_1 _20242_ (.B1(net4700),
    .Y(_05266_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .A2(net4603));
 sg13g2_nand3_1 _20243_ (.B(net4249),
    .C(_05266_),
    .A(net2012),
    .Y(_05267_));
 sg13g2_o21ai_1 _20244_ (.B1(net4618),
    .Y(_05268_),
    .A1(net2012),
    .A2(\soc_inst.cpu_core.mem_rs1_data[19] ));
 sg13g2_nand3_1 _20245_ (.B(_05267_),
    .C(_05268_),
    .A(_05072_),
    .Y(_05269_));
 sg13g2_mux2_1 _20246_ (.A0(_05269_),
    .A1(net2012),
    .S(net3854),
    .X(_02102_));
 sg13g2_o21ai_1 _20247_ (.B1(net4700),
    .Y(_05270_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .A2(net4604));
 sg13g2_nand3_1 _20248_ (.B(net4250),
    .C(_05270_),
    .A(net2212),
    .Y(_05271_));
 sg13g2_o21ai_1 _20249_ (.B1(net4618),
    .Y(_05272_),
    .A1(net2212),
    .A2(net1576));
 sg13g2_nand3_1 _20250_ (.B(_05271_),
    .C(_05272_),
    .A(_05077_),
    .Y(_05273_));
 sg13g2_mux2_1 _20251_ (.A0(_05273_),
    .A1(net2212),
    .S(net3854),
    .X(_02103_));
 sg13g2_o21ai_1 _20252_ (.B1(net4700),
    .Y(_05274_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .A2(net4603));
 sg13g2_nand3_1 _20253_ (.B(net4249),
    .C(_05274_),
    .A(net2329),
    .Y(_05275_));
 sg13g2_o21ai_1 _20254_ (.B1(net4618),
    .Y(_05276_),
    .A1(net2329),
    .A2(net2253));
 sg13g2_nand3_1 _20255_ (.B(_05275_),
    .C(_05276_),
    .A(_05082_),
    .Y(_05277_));
 sg13g2_mux2_1 _20256_ (.A0(_05277_),
    .A1(net2329),
    .S(net3854),
    .X(_02104_));
 sg13g2_o21ai_1 _20257_ (.B1(net4700),
    .Y(_05278_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .A2(net4604));
 sg13g2_nand3_1 _20258_ (.B(net4249),
    .C(_05278_),
    .A(net2231),
    .Y(_05279_));
 sg13g2_o21ai_1 _20259_ (.B1(net4618),
    .Y(_05280_),
    .A1(net2231),
    .A2(\soc_inst.cpu_core.mem_rs1_data[22] ));
 sg13g2_nand3_1 _20260_ (.B(_05279_),
    .C(_05280_),
    .A(_05087_),
    .Y(_05281_));
 sg13g2_mux2_1 _20261_ (.A0(_05281_),
    .A1(net2231),
    .S(net3854),
    .X(_02105_));
 sg13g2_o21ai_1 _20262_ (.B1(net4700),
    .Y(_05282_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .A2(net4603));
 sg13g2_nand3_1 _20263_ (.B(net4249),
    .C(_05282_),
    .A(net2120),
    .Y(_05283_));
 sg13g2_o21ai_1 _20264_ (.B1(net4618),
    .Y(_05284_),
    .A1(net2120),
    .A2(\soc_inst.cpu_core.mem_rs1_data[23] ));
 sg13g2_nand3_1 _20265_ (.B(_05283_),
    .C(_05284_),
    .A(_05092_),
    .Y(_05285_));
 sg13g2_mux2_1 _20266_ (.A0(_05285_),
    .A1(net2120),
    .S(net3854),
    .X(_02106_));
 sg13g2_nor3_1 _20267_ (.A(net3853),
    .B(_07217_),
    .C(_08540_),
    .Y(_05286_));
 sg13g2_nand3_1 _20268_ (.B(_06733_),
    .C(net4168),
    .A(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .Y(_05287_));
 sg13g2_o21ai_1 _20269_ (.B1(_05287_),
    .Y(_02107_),
    .A1(_05647_),
    .A2(_05286_));
 sg13g2_nor2_1 _20270_ (.A(net2057),
    .B(net1005),
    .Y(_05288_));
 sg13g2_a21oi_1 _20271_ (.A1(net1005),
    .A2(net4226),
    .Y(_05289_),
    .B1(net4617));
 sg13g2_o21ai_1 _20272_ (.B1(net4698),
    .Y(_05290_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[25] ),
    .A2(net4605));
 sg13g2_nand3_1 _20273_ (.B(net4253),
    .C(_05290_),
    .A(net2057),
    .Y(_05291_));
 sg13g2_o21ai_1 _20274_ (.B1(_05291_),
    .Y(_05292_),
    .A1(_05288_),
    .A2(_05289_));
 sg13g2_mux2_1 _20275_ (.A0(_05292_),
    .A1(net2057),
    .S(net3853),
    .X(_02108_));
 sg13g2_o21ai_1 _20276_ (.B1(net4699),
    .Y(_05293_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .A2(net4611));
 sg13g2_nand3_1 _20277_ (.B(net4257),
    .C(_05293_),
    .A(net2109),
    .Y(_05294_));
 sg13g2_or2_1 _20278_ (.X(_05295_),
    .B(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .A(\soc_inst.cpu_core.csr_file.mstatus[26] ));
 sg13g2_a22oi_1 _20279_ (.Y(_05296_),
    .B1(net4617),
    .B2(_05295_),
    .A2(net4227),
    .A1(\soc_inst.cpu_core.mem_rs1_data[26] ));
 sg13g2_a21oi_1 _20280_ (.A1(_05294_),
    .A2(_05296_),
    .Y(_05297_),
    .B1(net3856));
 sg13g2_a21o_1 _20281_ (.A2(net3856),
    .A1(net2109),
    .B1(_05297_),
    .X(_02109_));
 sg13g2_nor2_1 _20282_ (.A(net2063),
    .B(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .Y(_05298_));
 sg13g2_a21oi_1 _20283_ (.A1(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .A2(net4226),
    .Y(_05299_),
    .B1(net4617));
 sg13g2_o21ai_1 _20284_ (.B1(net4699),
    .Y(_05300_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .A2(net4605));
 sg13g2_nand3_1 _20285_ (.B(net4252),
    .C(_05300_),
    .A(net2063),
    .Y(_05301_));
 sg13g2_o21ai_1 _20286_ (.B1(_05301_),
    .Y(_05302_),
    .A1(_05298_),
    .A2(_05299_));
 sg13g2_mux2_1 _20287_ (.A0(_05302_),
    .A1(net2063),
    .S(net3853),
    .X(_02110_));
 sg13g2_nor2_1 _20288_ (.A(net2436),
    .B(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .Y(_05303_));
 sg13g2_a21oi_1 _20289_ (.A1(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .A2(net4226),
    .Y(_05304_),
    .B1(net4617));
 sg13g2_o21ai_1 _20290_ (.B1(net4698),
    .Y(_05305_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .A2(net4605));
 sg13g2_nand3_1 _20291_ (.B(net4253),
    .C(_05305_),
    .A(net2436),
    .Y(_05306_));
 sg13g2_o21ai_1 _20292_ (.B1(_05306_),
    .Y(_05307_),
    .A1(_05303_),
    .A2(_05304_));
 sg13g2_mux2_1 _20293_ (.A0(_05307_),
    .A1(net2436),
    .S(net3853),
    .X(_02111_));
 sg13g2_nor2_1 _20294_ (.A(net1937),
    .B(net1095),
    .Y(_05308_));
 sg13g2_a21oi_1 _20295_ (.A1(net1095),
    .A2(net4226),
    .Y(_05309_),
    .B1(net4617));
 sg13g2_o21ai_1 _20296_ (.B1(net4698),
    .Y(_05310_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[29] ),
    .A2(net4605));
 sg13g2_nand3_1 _20297_ (.B(net4253),
    .C(_05310_),
    .A(net1937),
    .Y(_05311_));
 sg13g2_o21ai_1 _20298_ (.B1(_05311_),
    .Y(_05312_),
    .A1(_05308_),
    .A2(_05309_));
 sg13g2_mux2_1 _20299_ (.A0(_05312_),
    .A1(net1937),
    .S(net3853),
    .X(_02112_));
 sg13g2_nor2_1 _20300_ (.A(net2410),
    .B(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .Y(_05313_));
 sg13g2_a21oi_1 _20301_ (.A1(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .A2(net4227),
    .Y(_05314_),
    .B1(net4623));
 sg13g2_o21ai_1 _20302_ (.B1(net4699),
    .Y(_05315_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .A2(net4607));
 sg13g2_nand3_1 _20303_ (.B(net4254),
    .C(_05315_),
    .A(net2410),
    .Y(_05316_));
 sg13g2_o21ai_1 _20304_ (.B1(_05316_),
    .Y(_05317_),
    .A1(_05313_),
    .A2(_05314_));
 sg13g2_mux2_1 _20305_ (.A0(_05317_),
    .A1(net2410),
    .S(net3856),
    .X(_02113_));
 sg13g2_nor2_1 _20306_ (.A(net2233),
    .B(net4879),
    .Y(_05318_));
 sg13g2_a21oi_1 _20307_ (.A1(net4879),
    .A2(net4227),
    .Y(_05319_),
    .B1(net4617));
 sg13g2_o21ai_1 _20308_ (.B1(net4699),
    .Y(_05320_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .A2(net4607));
 sg13g2_nand3_1 _20309_ (.B(net4254),
    .C(_05320_),
    .A(net2233),
    .Y(_05321_));
 sg13g2_o21ai_1 _20310_ (.B1(_05321_),
    .Y(_05322_),
    .A1(_05318_),
    .A2(_05319_));
 sg13g2_mux2_1 _20311_ (.A0(_05322_),
    .A1(net2233),
    .S(net3853),
    .X(_02114_));
 sg13g2_o21ai_1 _20312_ (.B1(net5465),
    .Y(_05323_),
    .A1(net4760),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ));
 sg13g2_a21oi_1 _20313_ (.A1(_05385_),
    .A2(net4760),
    .Y(_02115_),
    .B1(_05323_));
 sg13g2_o21ai_1 _20314_ (.B1(net5465),
    .Y(_05324_),
    .A1(net4760),
    .A2(net658));
 sg13g2_a21oi_1 _20315_ (.A1(_05384_),
    .A2(net4760),
    .Y(_02116_),
    .B1(_05324_));
 sg13g2_o21ai_1 _20316_ (.B1(net5465),
    .Y(_05325_),
    .A1(net4761),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ));
 sg13g2_a21oi_1 _20317_ (.A1(_05383_),
    .A2(net4760),
    .Y(_02117_),
    .B1(_05325_));
 sg13g2_o21ai_1 _20318_ (.B1(net5464),
    .Y(_05326_),
    .A1(net4761),
    .A2(net661));
 sg13g2_a21oi_1 _20319_ (.A1(_05382_),
    .A2(net4761),
    .Y(_02118_),
    .B1(net662));
 sg13g2_o21ai_1 _20320_ (.B1(net5435),
    .Y(_05327_),
    .A1(net4760),
    .A2(net679));
 sg13g2_a21oi_1 _20321_ (.A1(_05381_),
    .A2(net4761),
    .Y(_02119_),
    .B1(_05327_));
 sg13g2_o21ai_1 _20322_ (.B1(net5435),
    .Y(_05328_),
    .A1(net4760),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ));
 sg13g2_a21oi_1 _20323_ (.A1(_05380_),
    .A2(net4760),
    .Y(_02120_),
    .B1(_05328_));
 sg13g2_o21ai_1 _20324_ (.B1(net5464),
    .Y(_05329_),
    .A1(net4761),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ));
 sg13g2_a21oi_1 _20325_ (.A1(_05379_),
    .A2(net4761),
    .Y(_02121_),
    .B1(_05329_));
 sg13g2_o21ai_1 _20326_ (.B1(net5464),
    .Y(_05330_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ),
    .A2(net4762));
 sg13g2_a21oi_1 _20327_ (.A1(_05378_),
    .A2(net4762),
    .Y(_02122_),
    .B1(_05330_));
 sg13g2_nor2_2 _20328_ (.A(_05503_),
    .B(_06111_),
    .Y(_05331_));
 sg13g2_nand2_1 _20329_ (.Y(_05332_),
    .A(net1120),
    .B(_06110_));
 sg13g2_nor2b_2 _20330_ (.A(net1114),
    .B_N(net5473),
    .Y(_05333_));
 sg13g2_o21ai_1 _20331_ (.B1(net4658),
    .Y(_05334_),
    .A1(net620),
    .A2(net3948));
 sg13g2_a21oi_1 _20332_ (.A1(_05385_),
    .A2(net3948),
    .Y(_02123_),
    .B1(net621));
 sg13g2_o21ai_1 _20333_ (.B1(net4658),
    .Y(_05335_),
    .A1(net620),
    .A2(_05331_));
 sg13g2_a21oi_1 _20334_ (.A1(_05383_),
    .A2(_05331_),
    .Y(_02124_),
    .B1(net1115));
 sg13g2_o21ai_1 _20335_ (.B1(net4658),
    .Y(_05336_),
    .A1(net655),
    .A2(net3948));
 sg13g2_a21oi_1 _20336_ (.A1(_05383_),
    .A2(net3948),
    .Y(_02125_),
    .B1(_05336_));
 sg13g2_o21ai_1 _20337_ (.B1(net4658),
    .Y(_05337_),
    .A1(net655),
    .A2(_05331_));
 sg13g2_a21oi_1 _20338_ (.A1(_05381_),
    .A2(_05331_),
    .Y(_02126_),
    .B1(net656));
 sg13g2_o21ai_1 _20339_ (.B1(net4658),
    .Y(_05338_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ),
    .A2(net3948));
 sg13g2_a21oi_1 _20340_ (.A1(_05381_),
    .A2(net3948),
    .Y(_02127_),
    .B1(_05338_));
 sg13g2_o21ai_1 _20341_ (.B1(net4658),
    .Y(_05339_),
    .A1(net1299),
    .A2(net3948));
 sg13g2_a21oi_1 _20342_ (.A1(_05380_),
    .A2(net3948),
    .Y(_02128_),
    .B1(_05339_));
 sg13g2_o21ai_1 _20343_ (.B1(net4658),
    .Y(_05340_),
    .A1(net1276),
    .A2(net3949));
 sg13g2_a21oi_1 _20344_ (.A1(_05379_),
    .A2(net3949),
    .Y(_02129_),
    .B1(_05340_));
 sg13g2_o21ai_1 _20345_ (.B1(_05333_),
    .Y(_05341_),
    .A1(net1454),
    .A2(net3949));
 sg13g2_a21oi_1 _20346_ (.A1(_05378_),
    .A2(net3949),
    .Y(_02130_),
    .B1(_05341_));
 sg13g2_nor2_1 _20347_ (.A(net4762),
    .B(net938),
    .Y(_05342_));
 sg13g2_nand2_2 _20348_ (.Y(_05343_),
    .A(net4658),
    .B(_05342_));
 sg13g2_inv_1 _20349_ (.Y(_05344_),
    .A(_05343_));
 sg13g2_xor2_1 _20350_ (.B(_05332_),
    .A(net2124),
    .X(_05345_));
 sg13g2_nor2_1 _20351_ (.A(_05343_),
    .B(_05345_),
    .Y(_02131_));
 sg13g2_a21oi_1 _20352_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ),
    .A2(_05331_),
    .Y(_05346_),
    .B1(net522));
 sg13g2_and3_1 _20353_ (.X(_05347_),
    .A(net522),
    .B(net2124),
    .C(_05331_));
 sg13g2_nor3_1 _20354_ (.A(_05343_),
    .B(net523),
    .C(_05347_),
    .Y(_02132_));
 sg13g2_nand2_1 _20355_ (.Y(_05348_),
    .A(net2613),
    .B(_05347_));
 sg13g2_o21ai_1 _20356_ (.B1(_05344_),
    .Y(_05349_),
    .A1(net2613),
    .A2(_05347_));
 sg13g2_nor2b_1 _20357_ (.A(_05349_),
    .B_N(_05348_),
    .Y(_02133_));
 sg13g2_xnor2_1 _20358_ (.Y(_05350_),
    .A(_05377_),
    .B(_05348_));
 sg13g2_nor2_1 _20359_ (.A(_05343_),
    .B(net2598),
    .Y(_02134_));
 sg13g2_o21ai_1 _20360_ (.B1(net5438),
    .Y(_05351_),
    .A1(net1454),
    .A2(_06100_));
 sg13g2_a21oi_1 _20361_ (.A1(_05373_),
    .A2(_06073_),
    .Y(_02135_),
    .B1(_05351_));
 sg13g2_nor4_1 _20362_ (.A(net2577),
    .B(net4762),
    .C(net938),
    .D(net1120),
    .Y(_05352_));
 sg13g2_a21oi_1 _20363_ (.A1(_05503_),
    .A2(_05342_),
    .Y(_05353_),
    .B1(_05376_));
 sg13g2_nor3_1 _20364_ (.A(_06112_),
    .B(_05352_),
    .C(_05353_),
    .Y(_02136_));
 sg13g2_and2_1 _20365_ (.A(net2180),
    .B(_05353_),
    .X(_05354_));
 sg13g2_nor2_1 _20366_ (.A(net2180),
    .B(_05353_),
    .Y(_05355_));
 sg13g2_nor3_1 _20367_ (.A(net3947),
    .B(_05354_),
    .C(net2181),
    .Y(_02137_));
 sg13g2_and2_1 _20368_ (.A(net2430),
    .B(_05354_),
    .X(_05356_));
 sg13g2_nor2_1 _20369_ (.A(net2430),
    .B(_05354_),
    .Y(_05357_));
 sg13g2_nor3_1 _20370_ (.A(net3947),
    .B(_05356_),
    .C(_05357_),
    .Y(_02138_));
 sg13g2_and2_1 _20371_ (.A(net2112),
    .B(_05356_),
    .X(_05358_));
 sg13g2_nor2_1 _20372_ (.A(net2112),
    .B(_05356_),
    .Y(_05359_));
 sg13g2_nor3_1 _20373_ (.A(net3947),
    .B(net2113),
    .C(_05359_),
    .Y(_02139_));
 sg13g2_and2_1 _20374_ (.A(net1896),
    .B(_05358_),
    .X(_05360_));
 sg13g2_nor2_1 _20375_ (.A(net1896),
    .B(_05358_),
    .Y(_05361_));
 sg13g2_nor3_1 _20376_ (.A(net3947),
    .B(_05360_),
    .C(net2114),
    .Y(_02140_));
 sg13g2_and2_1 _20377_ (.A(net2198),
    .B(_05360_),
    .X(_05362_));
 sg13g2_nor2_1 _20378_ (.A(net2198),
    .B(_05360_),
    .Y(_05363_));
 sg13g2_nor3_1 _20379_ (.A(net3947),
    .B(_05362_),
    .C(_05363_),
    .Y(_02141_));
 sg13g2_and2_1 _20380_ (.A(net2132),
    .B(_05362_),
    .X(_05364_));
 sg13g2_nor2_1 _20381_ (.A(net2132),
    .B(_05362_),
    .Y(_05365_));
 sg13g2_nor3_1 _20382_ (.A(net3947),
    .B(_05364_),
    .C(net2133),
    .Y(_02142_));
 sg13g2_xnor2_1 _20383_ (.Y(_05366_),
    .A(net2679),
    .B(_05364_));
 sg13g2_nor2_1 _20384_ (.A(net3947),
    .B(_05366_),
    .Y(_02143_));
 sg13g2_nand3_1 _20385_ (.B(net2679),
    .C(_05364_),
    .A(net2929),
    .Y(_05367_));
 sg13g2_a21o_1 _20386_ (.A2(_05364_),
    .A1(net2679),
    .B1(net2929),
    .X(_05368_));
 sg13g2_and3_1 _20387_ (.X(_02144_),
    .A(_06113_),
    .B(_05367_),
    .C(_05368_));
 sg13g2_xor2_1 _20388_ (.B(_05367_),
    .A(net2795),
    .X(_05369_));
 sg13g2_nor2_1 _20389_ (.A(net3947),
    .B(net2796),
    .Y(_02145_));
 sg13g2_nand2b_1 _20390_ (.Y(_05370_),
    .B(net570),
    .A_N(net1532));
 sg13g2_nand2_1 _20391_ (.Y(_05371_),
    .A(net1532),
    .B(net1));
 sg13g2_nand3_1 _20392_ (.B(_05370_),
    .C(_05371_),
    .A(net5469),
    .Y(_02146_));
 sg13g2_o21ai_1 _20393_ (.B1(net5470),
    .Y(_05372_),
    .A1(_05373_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ));
 sg13g2_a21o_1 _20394_ (.A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .A1(net570),
    .B1(_05372_),
    .X(_02147_));
 sg13g2_xor2_1 _20395_ (.B(\soc_inst.spi_inst.state[0] ),
    .A(net520),
    .X(\soc_inst.spi_inst.next_state[1] ));
 sg13g2_dfrbpq_1 _20396_ (.RESET_B(net5436),
    .D(_00333_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][0] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _20397_ (.RESET_B(net5436),
    .D(_00334_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][1] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _20398_ (.RESET_B(net5437),
    .D(_00335_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][2] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _20399_ (.RESET_B(net5437),
    .D(_00336_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][3] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _20400_ (.RESET_B(net5428),
    .D(_00337_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][4] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _20401_ (.RESET_B(net5430),
    .D(_00338_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][5] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _20402_ (.RESET_B(net5425),
    .D(net1868),
    .Q(\soc_inst.pwm_inst.channel_duty[1][6] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _20403_ (.RESET_B(net5425),
    .D(_00340_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][7] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20404_ (.RESET_B(net5426),
    .D(_00341_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][8] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _20405_ (.RESET_B(net5408),
    .D(_00342_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][9] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _20406_ (.RESET_B(net5407),
    .D(net1189),
    .Q(\soc_inst.pwm_inst.channel_duty[1][10] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _20407_ (.RESET_B(net5411),
    .D(_00344_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][11] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20408_ (.RESET_B(net5411),
    .D(_00345_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][12] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _20409_ (.RESET_B(net5419),
    .D(net2314),
    .Q(\soc_inst.pwm_inst.channel_duty[1][13] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _20410_ (.RESET_B(net5432),
    .D(net2408),
    .Q(\soc_inst.pwm_inst.channel_duty[1][14] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _20411_ (.RESET_B(net5433),
    .D(_00348_),
    .Q(\soc_inst.pwm_inst.channel_duty[1][15] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _20412_ (.RESET_B(net5461),
    .D(net2279),
    .Q(\soc_inst.spi_inst.spi_sclk ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _20413_ (.RESET_B(net5459),
    .D(net750),
    .Q(\soc_inst.spi_inst.spi_mosi ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _20414_ (.RESET_B(net5456),
    .D(_00133_),
    .Q(\soc_inst.spi_inst.start_pending ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _20415_ (.RESET_B(net5452),
    .D(_00134_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[0] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20416_ (.RESET_B(net5454),
    .D(net225),
    .Q(\soc_inst.spi_inst.tx_shift_reg[1] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _20417_ (.RESET_B(net5454),
    .D(net324),
    .Q(\soc_inst.spi_inst.tx_shift_reg[2] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _20418_ (.RESET_B(net5454),
    .D(net274),
    .Q(\soc_inst.spi_inst.tx_shift_reg[3] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _20419_ (.RESET_B(net5454),
    .D(net239),
    .Q(\soc_inst.spi_inst.tx_shift_reg[4] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _20420_ (.RESET_B(net5452),
    .D(net560),
    .Q(\soc_inst.spi_inst.tx_shift_reg[5] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20421_ (.RESET_B(net5450),
    .D(net244),
    .Q(\soc_inst.spi_inst.tx_shift_reg[6] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20422_ (.RESET_B(net5450),
    .D(net171),
    .Q(\soc_inst.spi_inst.tx_shift_reg[7] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20423_ (.RESET_B(net5449),
    .D(net326),
    .Q(\soc_inst.spi_inst.tx_shift_reg[8] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20424_ (.RESET_B(net5449),
    .D(net302),
    .Q(\soc_inst.spi_inst.tx_shift_reg[9] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20425_ (.RESET_B(net5449),
    .D(net443),
    .Q(\soc_inst.spi_inst.tx_shift_reg[10] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20426_ (.RESET_B(net5449),
    .D(net216),
    .Q(\soc_inst.spi_inst.tx_shift_reg[11] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20427_ (.RESET_B(net5449),
    .D(net150),
    .Q(\soc_inst.spi_inst.tx_shift_reg[12] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20428_ (.RESET_B(net5449),
    .D(net439),
    .Q(\soc_inst.spi_inst.tx_shift_reg[13] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20429_ (.RESET_B(net5449),
    .D(net386),
    .Q(\soc_inst.spi_inst.tx_shift_reg[14] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20430_ (.RESET_B(net5454),
    .D(net270),
    .Q(\soc_inst.spi_inst.tx_shift_reg[15] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _20431_ (.RESET_B(net5461),
    .D(net119),
    .Q(\soc_inst.spi_inst.tx_shift_reg[16] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _20432_ (.RESET_B(net5476),
    .D(net188),
    .Q(\soc_inst.spi_inst.tx_shift_reg[17] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20433_ (.RESET_B(net5476),
    .D(net394),
    .Q(\soc_inst.spi_inst.tx_shift_reg[18] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20434_ (.RESET_B(net5476),
    .D(net166),
    .Q(\soc_inst.spi_inst.tx_shift_reg[19] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _20435_ (.RESET_B(net5476),
    .D(net114),
    .Q(\soc_inst.spi_inst.tx_shift_reg[20] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20436_ (.RESET_B(net5478),
    .D(net138),
    .Q(\soc_inst.spi_inst.tx_shift_reg[21] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20437_ (.RESET_B(net5477),
    .D(_00148_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[22] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20438_ (.RESET_B(net5477),
    .D(_00149_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[23] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _20439_ (.RESET_B(net5477),
    .D(net308),
    .Q(\soc_inst.spi_inst.tx_shift_reg[24] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _20440_ (.RESET_B(net5477),
    .D(net342),
    .Q(\soc_inst.spi_inst.tx_shift_reg[25] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _20441_ (.RESET_B(net5477),
    .D(_00152_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[26] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _20442_ (.RESET_B(net5477),
    .D(net233),
    .Q(\soc_inst.spi_inst.tx_shift_reg[27] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _20443_ (.RESET_B(net5477),
    .D(_00154_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[28] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20444_ (.RESET_B(net5477),
    .D(net340),
    .Q(\soc_inst.spi_inst.tx_shift_reg[29] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _20445_ (.RESET_B(net5478),
    .D(net349),
    .Q(\soc_inst.spi_inst.tx_shift_reg[30] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _20446_ (.RESET_B(net5478),
    .D(net367),
    .Q(\soc_inst.spi_inst.tx_shift_reg[31] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _20447_ (.RESET_B(net5462),
    .D(_00350_),
    .Q(\soc_inst.spi_inst.bit_counter[0] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20448_ (.RESET_B(net5457),
    .D(net819),
    .Q(\soc_inst.spi_inst.bit_counter[1] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20449_ (.RESET_B(net5457),
    .D(_00352_),
    .Q(\soc_inst.spi_inst.bit_counter[2] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _20450_ (.RESET_B(net5457),
    .D(net1985),
    .Q(\soc_inst.spi_inst.bit_counter[3] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _20451_ (.RESET_B(net5462),
    .D(_00354_),
    .Q(\soc_inst.spi_inst.bit_counter[4] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _20452_ (.RESET_B(net5457),
    .D(_00355_),
    .Q(\soc_inst.spi_inst.bit_counter[5] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _20453_ (.RESET_B(net5456),
    .D(net345),
    .Q(\soc_inst.spi_inst.state[0] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _20454_ (.RESET_B(net5456),
    .D(net521),
    .Q(\soc_inst.spi_inst.state[1] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _20455_ (.RESET_B(net5449),
    .D(_00356_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _20456_ (.RESET_B(net5446),
    .D(_00357_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _20457_ (.RESET_B(net5443),
    .D(_00358_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _20458_ (.RESET_B(net5440),
    .D(_00359_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _20459_ (.RESET_B(net5440),
    .D(_00360_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _20460_ (.RESET_B(net5439),
    .D(_00361_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _20461_ (.RESET_B(net5440),
    .D(_00362_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _20462_ (.RESET_B(net5439),
    .D(_00363_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _20463_ (.RESET_B(net5414),
    .D(_00364_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _20464_ (.RESET_B(net5415),
    .D(_00365_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _20465_ (.RESET_B(net5415),
    .D(_00366_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _20466_ (.RESET_B(net5415),
    .D(_00367_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _20467_ (.RESET_B(net5415),
    .D(_00368_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _20468_ (.RESET_B(net5415),
    .D(_00369_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _20469_ (.RESET_B(net5439),
    .D(_00370_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _20470_ (.RESET_B(net5440),
    .D(_00371_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _20471_ (.RESET_B(net5442),
    .D(_00372_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[16] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _20472_ (.RESET_B(net5446),
    .D(_00373_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[17] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _20473_ (.RESET_B(net5443),
    .D(_00374_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[18] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _20474_ (.RESET_B(net5443),
    .D(_00375_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[19] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _20475_ (.RESET_B(net5439),
    .D(_00376_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[20] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _20476_ (.RESET_B(net5439),
    .D(_00377_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[21] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _20477_ (.RESET_B(net5439),
    .D(_00378_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[22] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _20478_ (.RESET_B(net5439),
    .D(_00379_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[23] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _20479_ (.RESET_B(net5439),
    .D(_00380_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[24] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _20480_ (.RESET_B(net5445),
    .D(_00381_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[25] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _20481_ (.RESET_B(net5446),
    .D(_00382_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[26] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _20482_ (.RESET_B(net5446),
    .D(_00383_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[27] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _20483_ (.RESET_B(net5446),
    .D(_00384_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[28] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _20484_ (.RESET_B(net5446),
    .D(_00385_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[29] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _20485_ (.RESET_B(net5446),
    .D(_00386_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[30] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _20486_ (.RESET_B(net5446),
    .D(_00387_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[31] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _20487_ (.RESET_B(net5447),
    .D(_00388_),
    .Q(\soc_inst.spi_inst.cpha ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _20488_ (.RESET_B(net5454),
    .D(_00389_),
    .Q(\soc_inst.spi_ena ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _20489_ (.RESET_B(net5475),
    .D(_00390_),
    .Q(_00217_),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _20490_ (.RESET_B(net5475),
    .D(_00391_),
    .Q(_00218_),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _20491_ (.RESET_B(net5468),
    .D(net1684),
    .Q(_00219_),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _20492_ (.RESET_B(net5468),
    .D(net1434),
    .Q(_00220_),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _20493_ (.RESET_B(net5468),
    .D(_00394_),
    .Q(_00221_),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _20494_ (.RESET_B(net5468),
    .D(_00395_),
    .Q(\soc_inst.spi_inst.clock_divider[5] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _20495_ (.RESET_B(net5468),
    .D(_00396_),
    .Q(\soc_inst.spi_inst.clock_divider[6] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _20496_ (.RESET_B(net5447),
    .D(_00397_),
    .Q(\soc_inst.spi_inst.clock_divider[7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _20497_ (.RESET_B(net5456),
    .D(_00398_),
    .Q(\soc_inst.spi_inst.done ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _20498_ (.RESET_B(net5447),
    .D(_00399_),
    .Q(\soc_inst.spi_inst.cpol ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _20499_ (.RESET_B(net5462),
    .D(_10279_[0]),
    .Q(\soc_inst.spi_inst.spi_clk_en ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _20500_ (.RESET_B(net5456),
    .D(_00123_),
    .Q(\soc_inst.spi_inst.busy ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _20501_ (.RESET_B(net5473),
    .D(_00070_),
    .Q(\soc_inst.i2c_inst.clk_cnt[0] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _20502_ (.RESET_B(net5472),
    .D(_00071_),
    .Q(\soc_inst.i2c_inst.clk_cnt[1] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _20503_ (.RESET_B(net5472),
    .D(net712),
    .Q(\soc_inst.i2c_inst.clk_cnt[2] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _20504_ (.RESET_B(net5473),
    .D(_00073_),
    .Q(\soc_inst.i2c_inst.clk_cnt[3] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _20505_ (.RESET_B(net5473),
    .D(_00074_),
    .Q(\soc_inst.i2c_inst.clk_cnt[4] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _20506_ (.RESET_B(net5472),
    .D(_00075_),
    .Q(\soc_inst.i2c_inst.clk_cnt[5] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _20507_ (.RESET_B(net5472),
    .D(_00076_),
    .Q(\soc_inst.i2c_inst.clk_cnt[6] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _20508_ (.RESET_B(net5472),
    .D(_00077_),
    .Q(\soc_inst.i2c_inst.clk_cnt[7] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _20509_ (.RESET_B(net5460),
    .D(net469),
    .Q(\soc_inst.gpio_inst.int_pend_reg[0] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _20510_ (.RESET_B(net5466),
    .D(_00401_),
    .Q(\soc_inst.i2c_inst.ctrl_reg[2] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _20511_ (.RESET_B(net5466),
    .D(_00402_),
    .Q(\soc_inst.i2c_inst.ack_enable ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _20512_ (.RESET_B(net5468),
    .D(_00403_),
    .Q(\soc_inst.i2c_inst.ctrl_reg[4] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _20513_ (.RESET_B(net5466),
    .D(net160),
    .Q(\soc_inst.i2c_inst.arb_lost ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _20514_ (.RESET_B(net5474),
    .D(_10278_[0]),
    .Q(\soc_inst.i2c_inst.start_pending ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _20515_ (.RESET_B(net5466),
    .D(net670),
    .Q(\soc_inst.i2c_inst.data_reg[0] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _20516_ (.RESET_B(net5469),
    .D(net546),
    .Q(\soc_inst.i2c_inst.data_reg[1] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _20517_ (.RESET_B(net5469),
    .D(net1524),
    .Q(\soc_inst.i2c_inst.data_reg[2] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _20518_ (.RESET_B(net5464),
    .D(net653),
    .Q(\soc_inst.i2c_inst.data_reg[3] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _20519_ (.RESET_B(net5464),
    .D(net493),
    .Q(\soc_inst.i2c_inst.data_reg[4] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _20520_ (.RESET_B(net5464),
    .D(net537),
    .Q(\soc_inst.i2c_inst.data_reg[5] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _20521_ (.RESET_B(net5464),
    .D(net1693),
    .Q(\soc_inst.i2c_inst.data_reg[6] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _20522_ (.RESET_B(net5467),
    .D(_00085_),
    .Q(\soc_inst.i2c_inst.data_reg[7] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _20523_ (.RESET_B(net5471),
    .D(_00405_),
    .Q(_00222_),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _20524_ (.RESET_B(net5471),
    .D(net1726),
    .Q(_00223_),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _20525_ (.RESET_B(net5471),
    .D(net1619),
    .Q(_00224_),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _20526_ (.RESET_B(net5471),
    .D(net1953),
    .Q(_00225_),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _20527_ (.RESET_B(net5471),
    .D(_00409_),
    .Q(_00226_),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _20528_ (.RESET_B(net5471),
    .D(_00410_),
    .Q(\soc_inst.i2c_inst.prescale_reg[5] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _20529_ (.RESET_B(net5471),
    .D(net2138),
    .Q(\soc_inst.i2c_inst.prescale_reg[6] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _20530_ (.RESET_B(net5471),
    .D(_00412_),
    .Q(_00227_),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _20531_ (.RESET_B(net5479),
    .D(_10277_[0]),
    .Q(\soc_inst.i2c_inst.restart_pending ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _20532_ (.RESET_B(net5466),
    .D(_02148_),
    .Q(\soc_inst.i2c_inst.shift_reg[0] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _20533_ (.RESET_B(net5470),
    .D(net2148),
    .Q(\soc_inst.i2c_inst.shift_reg[1] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _20534_ (.RESET_B(net5470),
    .D(_02150_),
    .Q(\soc_inst.i2c_inst.shift_reg[2] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _20535_ (.RESET_B(net5465),
    .D(_02151_),
    .Q(\soc_inst.i2c_inst.shift_reg[3] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _20536_ (.RESET_B(net5465),
    .D(net2310),
    .Q(\soc_inst.i2c_inst.shift_reg[4] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _20537_ (.RESET_B(net5464),
    .D(net2157),
    .Q(\soc_inst.i2c_inst.shift_reg[5] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _20538_ (.RESET_B(net5465),
    .D(_02154_),
    .Q(\soc_inst.i2c_inst.shift_reg[6] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _20539_ (.RESET_B(net5466),
    .D(_02155_),
    .Q(\soc_inst.i2c_inst.shift_reg[7] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _20540_ (.RESET_B(net5480),
    .D(_00413_),
    .Q(\soc_inst.i2c_inst.bit_cnt[0] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _20541_ (.RESET_B(net5480),
    .D(_00414_),
    .Q(\soc_inst.i2c_inst.bit_cnt[1] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _20542_ (.RESET_B(net5480),
    .D(_00415_),
    .Q(\soc_inst.i2c_inst.bit_cnt[2] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _20543_ (.RESET_B(net5480),
    .D(net1123),
    .Q(\soc_inst.i2c_inst.bit_cnt[3] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _20544_ (.RESET_B(net5474),
    .D(_00417_),
    .Q(_00228_),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _20545_ (.RESET_B(net5479),
    .D(net825),
    .Q(\soc_inst.i2c_inst.stop_pending ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _20546_ (.RESET_B(net5459),
    .D(_00418_),
    .Q(_00229_),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _20547_ (.RESET_B(net5467),
    .D(_00087_),
    .Q(\soc_inst.i2c_inst.transfer_done ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _20548_ (.RESET_B(net5434),
    .D(_00107_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][0] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _20549_ (.RESET_B(net5434),
    .D(_00114_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][1] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _20550_ (.RESET_B(net5435),
    .D(net912),
    .Q(\soc_inst.pwm_inst.channel_counter[1][2] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _20551_ (.RESET_B(net5428),
    .D(_00116_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][3] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _20552_ (.RESET_B(net5427),
    .D(_00117_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][4] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _20553_ (.RESET_B(net5428),
    .D(_00118_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][5] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _20554_ (.RESET_B(net5428),
    .D(net2448),
    .Q(\soc_inst.pwm_inst.channel_counter[1][6] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _20555_ (.RESET_B(net5425),
    .D(_00120_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][7] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _20556_ (.RESET_B(net5427),
    .D(_00121_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][8] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20557_ (.RESET_B(net5426),
    .D(_00122_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20558_ (.RESET_B(net5411),
    .D(net2273),
    .Q(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20559_ (.RESET_B(net5411),
    .D(_00109_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][11] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20560_ (.RESET_B(net5411),
    .D(net2394),
    .Q(\soc_inst.pwm_inst.channel_counter[1][12] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _20561_ (.RESET_B(net5432),
    .D(net2302),
    .Q(\soc_inst.pwm_inst.channel_counter[1][13] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _20562_ (.RESET_B(net5432),
    .D(_00112_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _20563_ (.RESET_B(net5432),
    .D(_00113_),
    .Q(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _20564_ (.RESET_B(net5437),
    .D(_00091_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _20565_ (.RESET_B(net5437),
    .D(_00098_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _20566_ (.RESET_B(net5437),
    .D(net1590),
    .Q(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _20567_ (.RESET_B(net5430),
    .D(_00100_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _20568_ (.RESET_B(net5430),
    .D(net2473),
    .Q(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _20569_ (.RESET_B(net5430),
    .D(net2297),
    .Q(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _20570_ (.RESET_B(net5425),
    .D(net2319),
    .Q(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _20571_ (.RESET_B(net5425),
    .D(_00104_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20572_ (.RESET_B(net5426),
    .D(_00105_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _20573_ (.RESET_B(net5407),
    .D(_00106_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _20574_ (.RESET_B(net5407),
    .D(net1381),
    .Q(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _20575_ (.RESET_B(net5411),
    .D(_00093_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _20576_ (.RESET_B(net5427),
    .D(_00094_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _20577_ (.RESET_B(net5427),
    .D(_00095_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _20578_ (.RESET_B(net5427),
    .D(_00096_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _20579_ (.RESET_B(net5432),
    .D(_00097_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _20580_ (.RESET_B(net5224),
    .D(_00419_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.ram_in_quad_mode ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _20581_ (.RESET_B(net5434),
    .D(_00420_),
    .Q(_00230_),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _20582_ (.RESET_B(net5437),
    .D(_00421_),
    .Q(_00231_),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _20583_ (.RESET_B(net5437),
    .D(_00422_),
    .Q(_00232_),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _20584_ (.RESET_B(net5430),
    .D(net1377),
    .Q(_00233_),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _20585_ (.RESET_B(net5430),
    .D(_00424_),
    .Q(_00234_),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _20586_ (.RESET_B(net5430),
    .D(_00425_),
    .Q(_00235_),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _20587_ (.RESET_B(net5425),
    .D(net1830),
    .Q(_00236_),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _20588_ (.RESET_B(net5426),
    .D(_00427_),
    .Q(_00237_),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _20589_ (.RESET_B(net5407),
    .D(_00428_),
    .Q(_00238_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20590_ (.RESET_B(net5407),
    .D(_00429_),
    .Q(_00239_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20591_ (.RESET_B(net5408),
    .D(net1672),
    .Q(_00240_),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _20592_ (.RESET_B(net5408),
    .D(net1564),
    .Q(_00241_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20593_ (.RESET_B(net5411),
    .D(net1486),
    .Q(_00242_),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _20594_ (.RESET_B(net5427),
    .D(net1766),
    .Q(_00243_),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _20595_ (.RESET_B(net5432),
    .D(net1832),
    .Q(_00244_),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _20596_ (.RESET_B(net5433),
    .D(_00435_),
    .Q(_00245_),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _20597_ (.RESET_B(net5435),
    .D(_00436_),
    .Q(_00246_),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _20598_ (.RESET_B(net5434),
    .D(_00437_),
    .Q(_00247_),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _20599_ (.RESET_B(net5434),
    .D(_00438_),
    .Q(_00248_),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _20600_ (.RESET_B(net5434),
    .D(net1746),
    .Q(_00249_),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _20601_ (.RESET_B(net5427),
    .D(_00440_),
    .Q(_00250_),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _20602_ (.RESET_B(net5430),
    .D(_00441_),
    .Q(_00251_),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _20603_ (.RESET_B(net5429),
    .D(net1696),
    .Q(_00252_),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _20604_ (.RESET_B(net5426),
    .D(_00443_),
    .Q(_00253_),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _20605_ (.RESET_B(net5426),
    .D(net1604),
    .Q(_00254_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20606_ (.RESET_B(net5407),
    .D(_00445_),
    .Q(_00255_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20607_ (.RESET_B(net5408),
    .D(net2025),
    .Q(_00256_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20608_ (.RESET_B(net5407),
    .D(_00447_),
    .Q(_00257_),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _20609_ (.RESET_B(net5419),
    .D(net1331),
    .Q(_00258_),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _20610_ (.RESET_B(net5427),
    .D(net1645),
    .Q(_00259_),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _20611_ (.RESET_B(net5432),
    .D(net1555),
    .Q(_00260_),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _20612_ (.RESET_B(net5433),
    .D(_00451_),
    .Q(_00261_),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _20613_ (.RESET_B(net5436),
    .D(_00452_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _20614_ (.RESET_B(net5436),
    .D(_00453_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][1] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _20615_ (.RESET_B(net5436),
    .D(_00454_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][2] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _20616_ (.RESET_B(net5431),
    .D(_00455_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _20617_ (.RESET_B(net5431),
    .D(_00456_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][4] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _20618_ (.RESET_B(net5431),
    .D(_00457_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _20619_ (.RESET_B(net5425),
    .D(net2323),
    .Q(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _20620_ (.RESET_B(net5425),
    .D(net883),
    .Q(\soc_inst.pwm_inst.channel_duty[0][7] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _20621_ (.RESET_B(net5426),
    .D(_00460_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _20622_ (.RESET_B(net5407),
    .D(_00461_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _20623_ (.RESET_B(net5408),
    .D(net2081),
    .Q(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _20624_ (.RESET_B(net5411),
    .D(_00463_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _20625_ (.RESET_B(net5412),
    .D(_00464_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][12] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _20626_ (.RESET_B(net5412),
    .D(net2294),
    .Q(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _20627_ (.RESET_B(net5432),
    .D(net2095),
    .Q(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _20628_ (.RESET_B(net5433),
    .D(_00467_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _20629_ (.RESET_B(net5414),
    .D(net2960),
    .Q(\soc_inst.cpu_core.csr_file.timer_interrupt ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _20630_ (.RESET_B(net5447),
    .D(net2483),
    .Q(\soc_inst.spi_inst.len_sel[0] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _20631_ (.RESET_B(net5447),
    .D(net2964),
    .Q(\soc_inst.spi_inst.len_sel[1] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _20632_ (.RESET_B(net5460),
    .D(net87),
    .Q(\soc_inst.gpio_inst.gpio_sync2[0] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _20633_ (.RESET_B(net5460),
    .D(net82),
    .Q(\soc_inst.gpio_inst.gpio_sync2[1] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _20634_ (.RESET_B(net5458),
    .D(net84),
    .Q(\soc_inst.gpio_inst.gpio_sync2[2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _20635_ (.RESET_B(net5479),
    .D(net86),
    .Q(\soc_inst.gpio_inst.gpio_sync2[3] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _20636_ (.RESET_B(net5459),
    .D(net83),
    .Q(\soc_inst.gpio_inst.gpio_sync2[4] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20637_ (.RESET_B(net5457),
    .D(net88),
    .Q(\soc_inst.gpio_inst.gpio_sync2[5] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _20638_ (.RESET_B(net5457),
    .D(net80),
    .Q(\soc_inst.gpio_inst.gpio_sync2[6] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _20639_ (.RESET_B(net5182),
    .D(_00470_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _20640_ (.RESET_B(net5192),
    .D(_00471_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _20641_ (.RESET_B(net5183),
    .D(_00472_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _20642_ (.RESET_B(net5191),
    .D(_00473_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _20643_ (.RESET_B(net5219),
    .D(_00474_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _20644_ (.RESET_B(net5200),
    .D(_00475_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _20645_ (.RESET_B(net5219),
    .D(_00476_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _20646_ (.RESET_B(net5201),
    .D(_00477_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _20647_ (.RESET_B(net5148),
    .D(_00478_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _20648_ (.RESET_B(net5206),
    .D(_00479_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][9] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _20649_ (.RESET_B(net5175),
    .D(_00480_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _20650_ (.RESET_B(net5180),
    .D(_00481_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _20651_ (.RESET_B(net5208),
    .D(_00482_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _20652_ (.RESET_B(net5145),
    .D(_00483_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _20653_ (.RESET_B(net5206),
    .D(_00484_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _20654_ (.RESET_B(net5168),
    .D(_00485_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _20655_ (.RESET_B(net5144),
    .D(_00486_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _20656_ (.RESET_B(net5159),
    .D(_00487_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _20657_ (.RESET_B(net5129),
    .D(_00488_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _20658_ (.RESET_B(net5137),
    .D(_00489_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _20659_ (.RESET_B(net5131),
    .D(_00490_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _20660_ (.RESET_B(net5159),
    .D(_00491_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _20661_ (.RESET_B(net5142),
    .D(_00492_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][22] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _20662_ (.RESET_B(net5132),
    .D(_00493_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _20663_ (.RESET_B(net5154),
    .D(_00494_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _20664_ (.RESET_B(net5207),
    .D(_00495_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _20665_ (.RESET_B(net5184),
    .D(_00496_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _20666_ (.RESET_B(net5151),
    .D(_00497_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _20667_ (.RESET_B(net5141),
    .D(_00498_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][28] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _20668_ (.RESET_B(net5167),
    .D(_00499_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _20669_ (.RESET_B(net5186),
    .D(_00500_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _20670_ (.RESET_B(net5152),
    .D(_00501_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _20671_ (.RESET_B(net5459),
    .D(_00502_),
    .Q(\soc_inst.gpio_bidir_oe [0]),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _20672_ (.RESET_B(net5455),
    .D(_00503_),
    .Q(\soc_inst.gpio_bidir_out [0]),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _20673_ (.RESET_B(net5458),
    .D(_00504_),
    .Q(\soc_inst.gpio_inst.gpio_out[0] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _20674_ (.RESET_B(net5455),
    .D(net2593),
    .Q(\soc_inst.gpio_inst.gpio_out[1] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _20675_ (.RESET_B(net5458),
    .D(net1828),
    .Q(\soc_inst.gpio_inst.gpio_out[2] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _20676_ (.RESET_B(net5454),
    .D(_00507_),
    .Q(\soc_inst.gpio_inst.gpio_out[3] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _20677_ (.RESET_B(net5456),
    .D(_00508_),
    .Q(\soc_inst.gpio_inst.gpio_out[4] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _20678_ (.RESET_B(net5456),
    .D(_00509_),
    .Q(\soc_inst.gpio_inst.gpio_out[5] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _20679_ (.RESET_B(net5460),
    .D(net13),
    .Q(\soc_inst.gpio_inst.gpio_sync1[0] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _20680_ (.RESET_B(net5460),
    .D(net3),
    .Q(\soc_inst.gpio_inst.gpio_sync1[1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _20681_ (.RESET_B(net5455),
    .D(net4),
    .Q(\soc_inst.gpio_inst.gpio_sync1[2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _20682_ (.RESET_B(net5461),
    .D(net5),
    .Q(\soc_inst.gpio_inst.gpio_sync1[3] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _20683_ (.RESET_B(net5458),
    .D(net6),
    .Q(\soc_inst.gpio_inst.gpio_sync1[4] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20684_ (.RESET_B(net5451),
    .D(net7),
    .Q(\soc_inst.gpio_inst.gpio_sync1[5] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _20685_ (.RESET_B(net5457),
    .D(net8),
    .Q(\soc_inst.gpio_inst.gpio_sync1[6] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _20686_ (.RESET_B(net5476),
    .D(_00069_),
    .Q(\soc_inst.cpu_core.csr_file.external_interrupt ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _20687_ (.RESET_B(net5461),
    .D(_00510_),
    .Q(\soc_inst.gpio_inst.int_en_reg[0] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _20688_ (.RESET_B(net5460),
    .D(_00511_),
    .Q(\soc_inst.gpio_inst.int_en_reg[1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _20689_ (.RESET_B(net5458),
    .D(net2102),
    .Q(\soc_inst.gpio_inst.int_en_reg[2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _20690_ (.RESET_B(net5461),
    .D(_00513_),
    .Q(\soc_inst.gpio_inst.int_en_reg[3] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _20691_ (.RESET_B(net5458),
    .D(_00514_),
    .Q(\soc_inst.gpio_inst.int_en_reg[4] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _20692_ (.RESET_B(net5459),
    .D(_00515_),
    .Q(\soc_inst.gpio_inst.int_en_reg[5] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _20693_ (.RESET_B(net5461),
    .D(_00516_),
    .Q(\soc_inst.gpio_inst.int_en_reg[6] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _20694_ (.RESET_B(net5374),
    .D(_00517_),
    .Q(\soc_inst.mem_ctrl.spi_data_len[3] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _20695_ (.RESET_B(net5374),
    .D(net2742),
    .Q(\soc_inst.mem_ctrl.spi_data_len[4] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _20696_ (.RESET_B(net5374),
    .D(net2724),
    .Q(\soc_inst.mem_ctrl.spi_data_len[5] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _20697_ (.RESET_B(net5371),
    .D(net405),
    .Q(\soc_inst.mem_ctrl.next_instr_ready_reg ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _20698_ (.RESET_B(net5453),
    .D(net697),
    .Q(\soc_inst.mem_ctrl.spi_data_in[0] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20699_ (.RESET_B(net5453),
    .D(net466),
    .Q(\soc_inst.mem_ctrl.spi_data_in[1] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20700_ (.RESET_B(net5452),
    .D(net390),
    .Q(\soc_inst.mem_ctrl.spi_data_in[2] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20701_ (.RESET_B(net5453),
    .D(_00524_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[3] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20702_ (.RESET_B(net5453),
    .D(net531),
    .Q(\soc_inst.mem_ctrl.spi_data_in[4] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20703_ (.RESET_B(net5393),
    .D(net428),
    .Q(\soc_inst.mem_ctrl.spi_data_in[5] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _20704_ (.RESET_B(net5393),
    .D(_00527_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[6] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _20705_ (.RESET_B(net5450),
    .D(net413),
    .Q(\soc_inst.mem_ctrl.spi_data_in[7] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _20706_ (.RESET_B(net5452),
    .D(net672),
    .Q(\soc_inst.mem_ctrl.spi_data_in[8] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20707_ (.RESET_B(net5454),
    .D(net566),
    .Q(\soc_inst.mem_ctrl.spi_data_in[9] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20708_ (.RESET_B(net5450),
    .D(net779),
    .Q(\soc_inst.mem_ctrl.spi_data_in[10] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _20709_ (.RESET_B(net5450),
    .D(net361),
    .Q(\soc_inst.mem_ctrl.spi_data_in[11] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _20710_ (.RESET_B(net5451),
    .D(net581),
    .Q(\soc_inst.mem_ctrl.spi_data_in[12] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _20711_ (.RESET_B(net5450),
    .D(net558),
    .Q(\soc_inst.mem_ctrl.spi_data_in[13] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _20712_ (.RESET_B(net5451),
    .D(net535),
    .Q(\soc_inst.mem_ctrl.spi_data_in[14] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _20713_ (.RESET_B(net5450),
    .D(net489),
    .Q(\soc_inst.mem_ctrl.spi_data_in[15] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20714_ (.RESET_B(net5452),
    .D(net701),
    .Q(\soc_inst.mem_ctrl.spi_data_in[16] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20715_ (.RESET_B(net5394),
    .D(net693),
    .Q(\soc_inst.mem_ctrl.spi_data_in[17] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _20716_ (.RESET_B(net5452),
    .D(net407),
    .Q(\soc_inst.mem_ctrl.spi_data_in[18] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _20717_ (.RESET_B(net5452),
    .D(net415),
    .Q(\soc_inst.mem_ctrl.spi_data_in[19] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _20718_ (.RESET_B(net5395),
    .D(net613),
    .Q(\soc_inst.mem_ctrl.spi_data_in[20] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _20719_ (.RESET_B(net5452),
    .D(net437),
    .Q(\soc_inst.mem_ctrl.spi_data_in[21] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _20720_ (.RESET_B(net5396),
    .D(net378),
    .Q(\soc_inst.mem_ctrl.spi_data_in[22] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _20721_ (.RESET_B(net5390),
    .D(net347),
    .Q(\soc_inst.mem_ctrl.spi_data_in[23] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _20722_ (.RESET_B(net5389),
    .D(net297),
    .Q(\soc_inst.mem_ctrl.spi_data_in[24] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _20723_ (.RESET_B(net5390),
    .D(net328),
    .Q(\soc_inst.mem_ctrl.spi_data_in[25] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _20724_ (.RESET_B(net5390),
    .D(net314),
    .Q(\soc_inst.mem_ctrl.spi_data_in[26] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _20725_ (.RESET_B(net5389),
    .D(net214),
    .Q(\soc_inst.mem_ctrl.spi_data_in[27] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _20726_ (.RESET_B(net5389),
    .D(net265),
    .Q(\soc_inst.mem_ctrl.spi_data_in[28] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _20727_ (.RESET_B(net5389),
    .D(net227),
    .Q(\soc_inst.mem_ctrl.spi_data_in[29] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _20728_ (.RESET_B(net5376),
    .D(net278),
    .Q(\soc_inst.mem_ctrl.spi_data_in[30] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _20729_ (.RESET_B(net5376),
    .D(net355),
    .Q(\soc_inst.mem_ctrl.spi_data_in[31] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _20730_ (.RESET_B(net5302),
    .D(_00089_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.stop ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _20731_ (.RESET_B(net5378),
    .D(net471),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[5] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20732_ (.RESET_B(net5381),
    .D(net447),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[6] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20733_ (.RESET_B(net5345),
    .D(net435),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[8] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _20734_ (.RESET_B(net5345),
    .D(net479),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[9] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _20735_ (.RESET_B(net5382),
    .D(net464),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[10] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _20736_ (.RESET_B(net5360),
    .D(net2665),
    .Q(\soc_inst.cpu_core.csr_file.mepc[0] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _20737_ (.RESET_B(net5361),
    .D(_00059_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[1] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _20738_ (.RESET_B(net5330),
    .D(net2722),
    .Q(\soc_inst.cpu_core.csr_file.mepc[2] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _20739_ (.RESET_B(net5360),
    .D(_00061_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[3] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _20740_ (.RESET_B(net5360),
    .D(_00062_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[4] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _20741_ (.RESET_B(net5360),
    .D(_00027_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[0] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _20742_ (.RESET_B(net5360),
    .D(net2451),
    .Q(\soc_inst.cpu_core.csr_file.mcause[1] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _20743_ (.RESET_B(net5330),
    .D(_00049_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[2] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _20744_ (.RESET_B(net5330),
    .D(net2532),
    .Q(\soc_inst.cpu_core.csr_file.mcause[3] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _20745_ (.RESET_B(net5383),
    .D(_00052_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[4] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20746_ (.RESET_B(net5383),
    .D(_00053_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[5] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20747_ (.RESET_B(net5383),
    .D(_00054_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[6] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20748_ (.RESET_B(net5351),
    .D(_00055_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[7] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _20749_ (.RESET_B(net5351),
    .D(_00056_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[8] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20750_ (.RESET_B(net5352),
    .D(_00057_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[9] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20751_ (.RESET_B(net5351),
    .D(_00028_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20752_ (.RESET_B(net5351),
    .D(_00029_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[11] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _20753_ (.RESET_B(net5417),
    .D(_00030_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[12] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _20754_ (.RESET_B(net5349),
    .D(_00031_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[13] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _20755_ (.RESET_B(net5348),
    .D(_00032_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[14] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _20756_ (.RESET_B(net5341),
    .D(_00033_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[15] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _20757_ (.RESET_B(net5403),
    .D(_00034_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[16] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _20758_ (.RESET_B(net5403),
    .D(_00035_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[17] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _20759_ (.RESET_B(net5402),
    .D(_00036_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[18] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _20760_ (.RESET_B(net5338),
    .D(_00037_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[19] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _20761_ (.RESET_B(net5338),
    .D(_00039_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[20] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _20762_ (.RESET_B(net5315),
    .D(net104),
    .Q(\soc_inst.cpu_core.csr_file.mcause[21] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _20763_ (.RESET_B(net5406),
    .D(_00041_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[22] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _20764_ (.RESET_B(net5317),
    .D(net121),
    .Q(\soc_inst.cpu_core.csr_file.mcause[23] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _20765_ (.RESET_B(net5342),
    .D(_00043_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[24] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _20766_ (.RESET_B(net5340),
    .D(_00044_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[25] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _20767_ (.RESET_B(net5349),
    .D(_00045_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[26] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _20768_ (.RESET_B(net5341),
    .D(_00046_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[27] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _20769_ (.RESET_B(net5342),
    .D(_00047_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[28] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _20770_ (.RESET_B(net5339),
    .D(_00048_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[29] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _20771_ (.RESET_B(net5342),
    .D(_00050_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[30] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _20772_ (.RESET_B(net5360),
    .D(net2675),
    .Q(\soc_inst.cpu_core.csr_file.mtval[0] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _20773_ (.RESET_B(net5360),
    .D(net2479),
    .Q(\soc_inst.cpu_core.csr_file.mtval[1] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _20774_ (.RESET_B(net5330),
    .D(_00066_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[2] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _20775_ (.RESET_B(net5330),
    .D(_00067_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[3] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _20776_ (.RESET_B(net5360),
    .D(net2697),
    .Q(\soc_inst.cpu_core.csr_file.mtval[4] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _20777_ (.RESET_B(net5361),
    .D(_00558_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[0] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _20778_ (.RESET_B(net5364),
    .D(_00559_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[1] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _20779_ (.RESET_B(net5361),
    .D(_00560_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[2] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _20780_ (.RESET_B(net5331),
    .D(_00561_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[3] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _20781_ (.RESET_B(net5364),
    .D(net1534),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[4] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _20782_ (.RESET_B(net5474),
    .D(net2176),
    .Q(\soc_inst.i2c_inst.state[0] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _20783_ (.RESET_B(net5474),
    .D(net2663),
    .Q(\soc_inst.i2c_inst.state[1] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _20784_ (.RESET_B(net5474),
    .D(_00565_),
    .Q(\soc_inst.i2c_inst.state[2] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _20785_ (.RESET_B(net5474),
    .D(_00566_),
    .Q(\soc_inst.i2c_inst.state[3] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _20786_ (.RESET_B(net5392),
    .D(net1908),
    .Q(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20787_ (.RESET_B(net5387),
    .D(net2700),
    .Q(\soc_inst.mem_ctrl.spi_addr[1] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _20788_ (.RESET_B(net5386),
    .D(net2691),
    .Q(\soc_inst.mem_ctrl.spi_addr[2] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _20789_ (.RESET_B(net5392),
    .D(net2573),
    .Q(\soc_inst.mem_ctrl.spi_addr[3] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20790_ (.RESET_B(net5392),
    .D(net2504),
    .Q(\soc_inst.mem_ctrl.spi_addr[4] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _20791_ (.RESET_B(net5392),
    .D(net2336),
    .Q(\soc_inst.mem_ctrl.spi_addr[5] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20792_ (.RESET_B(net5385),
    .D(net2562),
    .Q(\soc_inst.mem_ctrl.spi_addr[6] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20793_ (.RESET_B(net5385),
    .D(net2512),
    .Q(\soc_inst.mem_ctrl.spi_addr[7] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _20794_ (.RESET_B(net5388),
    .D(net2495),
    .Q(\soc_inst.mem_ctrl.spi_addr[8] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _20795_ (.RESET_B(net5387),
    .D(net2388),
    .Q(\soc_inst.mem_ctrl.spi_addr[9] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _20796_ (.RESET_B(net5387),
    .D(net2327),
    .Q(\soc_inst.mem_ctrl.spi_addr[10] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20797_ (.RESET_B(net5387),
    .D(net2575),
    .Q(\soc_inst.mem_ctrl.spi_addr[11] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _20798_ (.RESET_B(net5392),
    .D(net2571),
    .Q(\soc_inst.mem_ctrl.spi_addr[12] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _20799_ (.RESET_B(net5392),
    .D(net2527),
    .Q(\soc_inst.mem_ctrl.spi_addr[13] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20800_ (.RESET_B(net5392),
    .D(net2422),
    .Q(\soc_inst.mem_ctrl.spi_addr[14] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _20801_ (.RESET_B(net5392),
    .D(net2508),
    .Q(\soc_inst.mem_ctrl.spi_addr[15] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20802_ (.RESET_B(net5393),
    .D(net2686),
    .Q(\soc_inst.mem_ctrl.spi_addr[16] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _20803_ (.RESET_B(net5388),
    .D(net2459),
    .Q(\soc_inst.mem_ctrl.spi_addr[17] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _20804_ (.RESET_B(net5388),
    .D(net2625),
    .Q(\soc_inst.mem_ctrl.spi_addr[18] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _20805_ (.RESET_B(net5388),
    .D(net2523),
    .Q(\soc_inst.mem_ctrl.spi_addr[19] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _20806_ (.RESET_B(net5387),
    .D(net2514),
    .Q(\soc_inst.mem_ctrl.spi_addr[20] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _20807_ (.RESET_B(net5387),
    .D(net2487),
    .Q(\soc_inst.mem_ctrl.spi_addr[21] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _20808_ (.RESET_B(net5387),
    .D(net1778),
    .Q(\soc_inst.mem_ctrl.spi_addr[22] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _20809_ (.RESET_B(net5387),
    .D(net2428),
    .Q(\soc_inst.mem_ctrl.spi_addr[23] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _20810_ (.RESET_B(net5368),
    .D(_00591_),
    .Q(\soc_inst.core_instr_data[0] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _20811_ (.RESET_B(net5367),
    .D(net544),
    .Q(\soc_inst.core_instr_data[1] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _20812_ (.RESET_B(net5285),
    .D(_00593_),
    .Q(\soc_inst.core_instr_data[2] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _20813_ (.RESET_B(net5285),
    .D(net2785),
    .Q(\soc_inst.core_instr_data[3] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _20814_ (.RESET_B(net5285),
    .D(_00595_),
    .Q(\soc_inst.core_instr_data[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _20815_ (.RESET_B(net5286),
    .D(net2891),
    .Q(\soc_inst.core_instr_data[5] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _20816_ (.RESET_B(net5305),
    .D(_00597_),
    .Q(\soc_inst.core_instr_data[6] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _20817_ (.RESET_B(net5285),
    .D(_00598_),
    .Q(\soc_inst.core_instr_data[7] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _20818_ (.RESET_B(net5301),
    .D(_00599_),
    .Q(\soc_inst.core_instr_data[8] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _20819_ (.RESET_B(net5303),
    .D(net948),
    .Q(\soc_inst.core_instr_data[9] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _20820_ (.RESET_B(net5283),
    .D(_00601_),
    .Q(\soc_inst.core_instr_data[10] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _20821_ (.RESET_B(net5303),
    .D(_00602_),
    .Q(\soc_inst.core_instr_data[11] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _20822_ (.RESET_B(net5305),
    .D(_00603_),
    .Q(\soc_inst.core_instr_data[12] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _20823_ (.RESET_B(net5303),
    .D(_00604_),
    .Q(\soc_inst.core_instr_data[13] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _20824_ (.RESET_B(net5303),
    .D(_00605_),
    .Q(\soc_inst.core_instr_data[14] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _20825_ (.RESET_B(net5305),
    .D(_00606_),
    .Q(\soc_inst.core_instr_data[15] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _20826_ (.RESET_B(net5283),
    .D(net199),
    .Q(\soc_inst.core_instr_data[16] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _20827_ (.RESET_B(net5273),
    .D(net392),
    .Q(\soc_inst.core_instr_data[17] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _20828_ (.RESET_B(net5283),
    .D(net363),
    .Q(\soc_inst.core_instr_data[18] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _20829_ (.RESET_B(net5283),
    .D(net396),
    .Q(\soc_inst.core_instr_data[19] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _20830_ (.RESET_B(net5273),
    .D(net371),
    .Q(\soc_inst.core_instr_data[20] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _20831_ (.RESET_B(net5272),
    .D(net310),
    .Q(\soc_inst.core_instr_data[21] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20832_ (.RESET_B(net5272),
    .D(net529),
    .Q(\soc_inst.core_instr_data[22] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20833_ (.RESET_B(net5272),
    .D(net192),
    .Q(\soc_inst.core_instr_data[23] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20834_ (.RESET_B(net5283),
    .D(net267),
    .Q(\soc_inst.core_instr_data[24] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _20835_ (.RESET_B(net5300),
    .D(_00616_),
    .Q(\soc_inst.core_instr_data[25] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _20836_ (.RESET_B(net5283),
    .D(net276),
    .Q(\soc_inst.core_instr_data[26] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _20837_ (.RESET_B(net5304),
    .D(_00618_),
    .Q(\soc_inst.core_instr_data[27] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _20838_ (.RESET_B(net5271),
    .D(net453),
    .Q(\soc_inst.core_instr_data[28] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _20839_ (.RESET_B(net5300),
    .D(_00620_),
    .Q(\soc_inst.core_instr_data[29] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _20840_ (.RESET_B(net5272),
    .D(net322),
    .Q(\soc_inst.core_instr_data[30] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20841_ (.RESET_B(net5272),
    .D(net320),
    .Q(\soc_inst.core_instr_data[31] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _20842_ (.RESET_B(net5443),
    .D(_00623_),
    .Q(\soc_inst.core_mem_rdata[0] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _20843_ (.RESET_B(net5384),
    .D(_00624_),
    .Q(\soc_inst.core_mem_rdata[1] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _20844_ (.RESET_B(net5380),
    .D(net290),
    .Q(\soc_inst.core_mem_rdata[2] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _20845_ (.RESET_B(net5372),
    .D(net295),
    .Q(\soc_inst.core_mem_rdata[3] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _20846_ (.RESET_B(net5442),
    .D(_00627_),
    .Q(\soc_inst.core_mem_rdata[4] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _20847_ (.RESET_B(net5381),
    .D(_00628_),
    .Q(\soc_inst.core_mem_rdata[5] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _20848_ (.RESET_B(net5384),
    .D(_00629_),
    .Q(\soc_inst.core_mem_rdata[6] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _20849_ (.RESET_B(net5381),
    .D(net763),
    .Q(\soc_inst.core_mem_rdata[7] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _20850_ (.RESET_B(net5382),
    .D(_00631_),
    .Q(\soc_inst.core_mem_rdata[8] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _20851_ (.RESET_B(net5385),
    .D(_00632_),
    .Q(\soc_inst.core_mem_rdata[9] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _20852_ (.RESET_B(net5384),
    .D(_00633_),
    .Q(\soc_inst.core_mem_rdata[10] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _20853_ (.RESET_B(net5385),
    .D(_00634_),
    .Q(\soc_inst.core_mem_rdata[11] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _20854_ (.RESET_B(net5383),
    .D(_00635_),
    .Q(\soc_inst.core_mem_rdata[12] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _20855_ (.RESET_B(net5382),
    .D(_00636_),
    .Q(\soc_inst.core_mem_rdata[13] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20856_ (.RESET_B(net5383),
    .D(_00637_),
    .Q(\soc_inst.core_mem_rdata[14] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _20857_ (.RESET_B(net5382),
    .D(_00638_),
    .Q(\soc_inst.core_mem_rdata[15] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20858_ (.RESET_B(net5416),
    .D(net1437),
    .Q(\soc_inst.core_mem_rdata[16] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20859_ (.RESET_B(net5413),
    .D(net1642),
    .Q(\soc_inst.core_mem_rdata[17] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _20860_ (.RESET_B(net5351),
    .D(net1321),
    .Q(\soc_inst.core_mem_rdata[18] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20861_ (.RESET_B(net5416),
    .D(net746),
    .Q(\soc_inst.core_mem_rdata[19] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _20862_ (.RESET_B(net5416),
    .D(net754),
    .Q(\soc_inst.core_mem_rdata[20] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20863_ (.RESET_B(net5351),
    .D(net552),
    .Q(\soc_inst.core_mem_rdata[21] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20864_ (.RESET_B(net5351),
    .D(net636),
    .Q(\soc_inst.core_mem_rdata[22] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20865_ (.RESET_B(net5351),
    .D(net903),
    .Q(\soc_inst.core_mem_rdata[23] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20866_ (.RESET_B(net5386),
    .D(_00647_),
    .Q(\soc_inst.core_mem_rdata[24] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _20867_ (.RESET_B(net5386),
    .D(net1512),
    .Q(\soc_inst.core_mem_rdata[25] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _20868_ (.RESET_B(net5386),
    .D(net1541),
    .Q(\soc_inst.core_mem_rdata[26] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20869_ (.RESET_B(net5353),
    .D(net640),
    .Q(\soc_inst.core_mem_rdata[27] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20870_ (.RESET_B(net5416),
    .D(net1467),
    .Q(\soc_inst.core_mem_rdata[28] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _20871_ (.RESET_B(net5416),
    .D(net1180),
    .Q(\soc_inst.core_mem_rdata[29] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _20872_ (.RESET_B(net5383),
    .D(net501),
    .Q(\soc_inst.core_mem_rdata[30] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20873_ (.RESET_B(net5353),
    .D(net1575),
    .Q(\soc_inst.core_mem_rdata[31] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _20874_ (.RESET_B(net5374),
    .D(net600),
    .Q(\soc_inst.mem_ctrl.spi_read_enable ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _20875_ (.RESET_B(net5374),
    .D(net676),
    .Q(\soc_inst.cpu_core.i_mem_ready ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _20876_ (.RESET_B(net5374),
    .D(net642),
    .Q(\soc_inst.mem_ctrl.instr_ready_reg ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _20877_ (.RESET_B(net5366),
    .D(net242),
    .Q(\soc_inst.mem_ctrl.next_instr_data[0] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _20878_ (.RESET_B(net5370),
    .D(net212),
    .Q(\soc_inst.mem_ctrl.next_instr_data[1] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _20879_ (.RESET_B(net5284),
    .D(net203),
    .Q(\soc_inst.mem_ctrl.next_instr_data[2] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _20880_ (.RESET_B(net5286),
    .D(net109),
    .Q(\soc_inst.mem_ctrl.next_instr_data[3] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _20881_ (.RESET_B(net5284),
    .D(net107),
    .Q(\soc_inst.mem_ctrl.next_instr_data[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _20882_ (.RESET_B(net5286),
    .D(net125),
    .Q(\soc_inst.mem_ctrl.next_instr_data[5] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _20883_ (.RESET_B(net5305),
    .D(net183),
    .Q(\soc_inst.mem_ctrl.next_instr_data[6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _20884_ (.RESET_B(net5284),
    .D(net283),
    .Q(\soc_inst.mem_ctrl.next_instr_data[7] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _20885_ (.RESET_B(net5301),
    .D(net140),
    .Q(\soc_inst.mem_ctrl.next_instr_data[8] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _20886_ (.RESET_B(net5303),
    .D(net333),
    .Q(\soc_inst.mem_ctrl.next_instr_data[9] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _20887_ (.RESET_B(net5283),
    .D(net180),
    .Q(\soc_inst.mem_ctrl.next_instr_data[10] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _20888_ (.RESET_B(net5301),
    .D(net201),
    .Q(\soc_inst.mem_ctrl.next_instr_data[11] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _20889_ (.RESET_B(net5303),
    .D(net229),
    .Q(\soc_inst.mem_ctrl.next_instr_data[12] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _20890_ (.RESET_B(net5302),
    .D(net235),
    .Q(\soc_inst.mem_ctrl.next_instr_data[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _20891_ (.RESET_B(net5302),
    .D(net288),
    .Q(\soc_inst.mem_ctrl.next_instr_data[14] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _20892_ (.RESET_B(net5284),
    .D(net256),
    .Q(\soc_inst.mem_ctrl.next_instr_data[15] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _20893_ (.RESET_B(net5282),
    .D(net205),
    .Q(\soc_inst.mem_ctrl.next_instr_data[16] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20894_ (.RESET_B(net5271),
    .D(net162),
    .Q(\soc_inst.mem_ctrl.next_instr_data[17] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _20895_ (.RESET_B(net5282),
    .D(net116),
    .Q(\soc_inst.mem_ctrl.next_instr_data[18] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _20896_ (.RESET_B(net5282),
    .D(net127),
    .Q(\soc_inst.mem_ctrl.next_instr_data[19] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _20897_ (.RESET_B(net5271),
    .D(net263),
    .Q(\soc_inst.mem_ctrl.next_instr_data[20] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _20898_ (.RESET_B(net5270),
    .D(net123),
    .Q(\soc_inst.mem_ctrl.next_instr_data[21] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20899_ (.RESET_B(net5270),
    .D(net252),
    .Q(\soc_inst.mem_ctrl.next_instr_data[22] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _20900_ (.RESET_B(net5271),
    .D(net185),
    .Q(\soc_inst.mem_ctrl.next_instr_data[23] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _20901_ (.RESET_B(net5282),
    .D(net147),
    .Q(\soc_inst.mem_ctrl.next_instr_data[24] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _20902_ (.RESET_B(net5304),
    .D(net299),
    .Q(\soc_inst.mem_ctrl.next_instr_data[25] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _20903_ (.RESET_B(net5282),
    .D(net231),
    .Q(\soc_inst.mem_ctrl.next_instr_data[26] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _20904_ (.RESET_B(net5366),
    .D(net223),
    .Q(\soc_inst.mem_ctrl.next_instr_data[27] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _20905_ (.RESET_B(net5270),
    .D(net248),
    .Q(\soc_inst.mem_ctrl.next_instr_data[28] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _20906_ (.RESET_B(net5301),
    .D(net254),
    .Q(\soc_inst.mem_ctrl.next_instr_data[29] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _20907_ (.RESET_B(net5270),
    .D(net190),
    .Q(\soc_inst.mem_ctrl.next_instr_data[30] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _20908_ (.RESET_B(net5270),
    .D(net250),
    .Q(\soc_inst.mem_ctrl.next_instr_data[31] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _20909_ (.RESET_B(net5376),
    .D(net2969),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _20910_ (.RESET_B(net5280),
    .D(_00088_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _20911_ (.RESET_B(net5222),
    .D(_00691_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _20912_ (.RESET_B(net5280),
    .D(_00692_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[1] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _20913_ (.RESET_B(net5280),
    .D(_00693_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _20914_ (.RESET_B(net5222),
    .D(_00694_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[3] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _20915_ (.RESET_B(net5222),
    .D(_00695_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _20916_ (.RESET_B(net5280),
    .D(_00696_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _20917_ (.RESET_B(net5278),
    .D(_00697_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _20918_ (.RESET_B(net5222),
    .D(_00698_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _20919_ (.RESET_B(net5214),
    .D(_00699_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _20920_ (.RESET_B(net5279),
    .D(_00700_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _20921_ (.RESET_B(net5278),
    .D(_00701_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _20922_ (.RESET_B(net5275),
    .D(_00702_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _20923_ (.RESET_B(net5214),
    .D(_00703_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[12] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _20924_ (.RESET_B(net5279),
    .D(_00704_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _20925_ (.RESET_B(net5276),
    .D(_00705_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _20926_ (.RESET_B(net5275),
    .D(_00706_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _20927_ (.RESET_B(net5222),
    .D(_00707_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _20928_ (.RESET_B(net5280),
    .D(_00708_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _20929_ (.RESET_B(net5276),
    .D(_00709_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _20930_ (.RESET_B(net5223),
    .D(_00710_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _20931_ (.RESET_B(net5222),
    .D(_00711_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _20932_ (.RESET_B(net5281),
    .D(_00712_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _20933_ (.RESET_B(net5279),
    .D(_00713_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _20934_ (.RESET_B(net5276),
    .D(_00714_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[23] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _20935_ (.RESET_B(net5222),
    .D(_00715_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _20936_ (.RESET_B(net5280),
    .D(_00716_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _20937_ (.RESET_B(net5279),
    .D(_00717_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _20938_ (.RESET_B(net5276),
    .D(_00718_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _20939_ (.RESET_B(net5222),
    .D(_00719_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[28] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _20940_ (.RESET_B(net5279),
    .D(_00720_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _20941_ (.RESET_B(net5281),
    .D(_00721_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[30] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _20942_ (.RESET_B(net5276),
    .D(_00722_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[31] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _20943_ (.RESET_B(net5218),
    .D(net98),
    .Q(\soc_inst.bus_spi_sclk ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _20944_ (.RESET_B(net5226),
    .D(net2863),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.is_write_op ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _20945_ (.RESET_B(net5224),
    .D(_00724_),
    .Q(_00262_),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _20946_ (.RESET_B(net5226),
    .D(net2736),
    .Q(\soc_inst.mem_ctrl.spi_done ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _20947_ (.RESET_B(net5218),
    .D(_00726_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _20948_ (.RESET_B(net5220),
    .D(_00727_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.write_mosi ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _20949_ (.RESET_B(net5378),
    .D(_00728_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[5] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _20950_ (.RESET_B(net5378),
    .D(_00729_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[6] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _20951_ (.RESET_B(net5344),
    .D(_00730_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[7] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _20952_ (.RESET_B(net5352),
    .D(_00731_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[8] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _20953_ (.RESET_B(net5345),
    .D(net156),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[9] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _20954_ (.RESET_B(net5382),
    .D(net143),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[10] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _20955_ (.RESET_B(net5344),
    .D(_00734_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[11] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _20956_ (.RESET_B(net5347),
    .D(_00735_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[12] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _20957_ (.RESET_B(net5328),
    .D(net221),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[13] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _20958_ (.RESET_B(net5352),
    .D(net177),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[14] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _20959_ (.RESET_B(net5347),
    .D(net134),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _20960_ (.RESET_B(net5338),
    .D(net208),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[16] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _20961_ (.RESET_B(net5338),
    .D(net261),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[17] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _20962_ (.RESET_B(net5334),
    .D(net195),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[18] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _20963_ (.RESET_B(net5334),
    .D(net174),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[19] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _20964_ (.RESET_B(net5335),
    .D(net286),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[20] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _20965_ (.RESET_B(net5315),
    .D(net131),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[21] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _20966_ (.RESET_B(net5334),
    .D(net293),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[22] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _20967_ (.RESET_B(net5317),
    .D(net153),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[23] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _20968_ (.RESET_B(net5348),
    .D(net1345),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[24] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _20969_ (.RESET_B(net5339),
    .D(_00748_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[25] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _20970_ (.RESET_B(net5348),
    .D(net1469),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[26] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _20971_ (.RESET_B(net5341),
    .D(net1706),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[27] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _20972_ (.RESET_B(net5342),
    .D(net1573),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[28] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _20973_ (.RESET_B(net5339),
    .D(_00752_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[29] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _20974_ (.RESET_B(net5342),
    .D(net1259),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[30] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _20975_ (.RESET_B(net5348),
    .D(net1333),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[31] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _20976_ (.RESET_B(net5218),
    .D(net2860),
    .Q(uio_oe[5]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _20977_ (.RESET_B(net5396),
    .D(_00756_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _20978_ (.RESET_B(net5394),
    .D(net1906),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20979_ (.RESET_B(net5394),
    .D(net1629),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _20980_ (.RESET_B(net5394),
    .D(net1526),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _20981_ (.RESET_B(net5396),
    .D(net1775),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _20982_ (.RESET_B(net5394),
    .D(net1792),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _20983_ (.RESET_B(net5394),
    .D(net1770),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _20984_ (.RESET_B(net5394),
    .D(net1951),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20985_ (.RESET_B(net5394),
    .D(net554),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _20986_ (.RESET_B(net5397),
    .D(net862),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _20987_ (.RESET_B(net5393),
    .D(net590),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _20988_ (.RESET_B(net5393),
    .D(net807),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _20989_ (.RESET_B(net5393),
    .D(net1396),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _20990_ (.RESET_B(net5393),
    .D(net1032),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _20991_ (.RESET_B(net5395),
    .D(net915),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _20992_ (.RESET_B(net5395),
    .D(net705),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _20993_ (.RESET_B(net5395),
    .D(net629),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _20994_ (.RESET_B(net5395),
    .D(net853),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _20995_ (.RESET_B(net5395),
    .D(net550),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[18] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _20996_ (.RESET_B(net5390),
    .D(net956),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _20997_ (.RESET_B(net5390),
    .D(net596),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _20998_ (.RESET_B(net5395),
    .D(net516),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _20999_ (.RESET_B(net5395),
    .D(net1813),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _21000_ (.RESET_B(net5390),
    .D(net741),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _21001_ (.RESET_B(net5389),
    .D(net1881),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _21002_ (.RESET_B(net5390),
    .D(net1561),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[25] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _21003_ (.RESET_B(net5390),
    .D(net1679),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _21004_ (.RESET_B(net5389),
    .D(net1780),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _21005_ (.RESET_B(net5391),
    .D(_00784_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _21006_ (.RESET_B(net5391),
    .D(_00785_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _21007_ (.RESET_B(net5391),
    .D(_00786_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _21008_ (.RESET_B(net5376),
    .D(_00787_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _21009_ (.RESET_B(net5225),
    .D(_00788_),
    .Q(uio_out[1]),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _21010_ (.RESET_B(net5226),
    .D(_00789_),
    .Q(uio_out[2]),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _21011_ (.RESET_B(net5221),
    .D(_00790_),
    .Q(uio_out[4]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _21012_ (.RESET_B(net5225),
    .D(net2780),
    .Q(uio_out[5]),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _21013_ (.RESET_B(net5217),
    .D(_00792_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.initialized ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _21014_ (.RESET_B(net5374),
    .D(_00793_),
    .Q(\soc_inst.mem_ctrl.spi_is_instr ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _21015_ (.RESET_B(net5224),
    .D(net2205),
    .Q(_00263_),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _21016_ (.RESET_B(net5221),
    .D(net2579),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _21017_ (.RESET_B(net5223),
    .D(net411),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _21018_ (.RESET_B(net5224),
    .D(_00001_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _21019_ (.RESET_B(net5223),
    .D(_00013_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _21020_ (.RESET_B(net5220),
    .D(net1035),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _21021_ (.RESET_B(net5226),
    .D(net2947),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _21022_ (.RESET_B(net5220),
    .D(_00016_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _21023_ (.RESET_B(net5220),
    .D(_00017_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _21024_ (.RESET_B(net5220),
    .D(_00018_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _21025_ (.RESET_B(net5226),
    .D(net2954),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _21026_ (.RESET_B(net5224),
    .D(net92),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _21027_ (.RESET_B(net5223),
    .D(_00011_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _21028_ (.RESET_B(net5217),
    .D(net475),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _21029_ (.RESET_B(net5225),
    .D(net2510),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _21030_ (.RESET_B(net5224),
    .D(_00005_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _21031_ (.RESET_B(net5364),
    .D(net2174),
    .Q(\soc_inst.core_instr_addr[0] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21032_ (.RESET_B(net5362),
    .D(net2534),
    .Q(\soc_inst.core_instr_addr[1] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _21033_ (.RESET_B(net5380),
    .D(_00796_),
    .Q(\soc_inst.core_instr_addr[2] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21034_ (.RESET_B(net5364),
    .D(net2497),
    .Q(\soc_inst.core_instr_addr[3] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21035_ (.RESET_B(net5380),
    .D(net2538),
    .Q(\soc_inst.core_instr_addr[4] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _21036_ (.RESET_B(net5380),
    .D(_00799_),
    .Q(\soc_inst.core_instr_addr[5] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21037_ (.RESET_B(net5380),
    .D(_00800_),
    .Q(\soc_inst.core_instr_addr[6] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _21038_ (.RESET_B(net5380),
    .D(_00801_),
    .Q(\soc_inst.core_instr_addr[7] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21039_ (.RESET_B(net5379),
    .D(_00802_),
    .Q(\soc_inst.core_instr_addr[8] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _21040_ (.RESET_B(net5346),
    .D(_00803_),
    .Q(\soc_inst.core_instr_addr[9] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _21041_ (.RESET_B(net5379),
    .D(_00804_),
    .Q(\soc_inst.core_instr_addr[10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _21042_ (.RESET_B(net5331),
    .D(_00805_),
    .Q(\soc_inst.core_instr_addr[11] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _21043_ (.RESET_B(net5344),
    .D(_00806_),
    .Q(\soc_inst.core_instr_addr[12] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _21044_ (.RESET_B(net5328),
    .D(_00807_),
    .Q(\soc_inst.core_instr_addr[13] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _21045_ (.RESET_B(net5352),
    .D(_00808_),
    .Q(\soc_inst.core_instr_addr[14] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _21046_ (.RESET_B(net5329),
    .D(_00809_),
    .Q(\soc_inst.core_instr_addr[15] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _21047_ (.RESET_B(net5337),
    .D(_00810_),
    .Q(\soc_inst.core_instr_addr[16] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _21048_ (.RESET_B(net5337),
    .D(_00811_),
    .Q(\soc_inst.core_instr_addr[17] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _21049_ (.RESET_B(net5319),
    .D(_00812_),
    .Q(\soc_inst.core_instr_addr[18] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _21050_ (.RESET_B(net5320),
    .D(_00813_),
    .Q(\soc_inst.core_instr_addr[19] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _21051_ (.RESET_B(net5336),
    .D(_00814_),
    .Q(\soc_inst.core_instr_addr[20] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _21052_ (.RESET_B(net5319),
    .D(_00815_),
    .Q(\soc_inst.core_instr_addr[21] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _21053_ (.RESET_B(net5336),
    .D(_00816_),
    .Q(\soc_inst.core_instr_addr[22] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _21054_ (.RESET_B(net5320),
    .D(_00817_),
    .Q(\soc_inst.core_instr_addr[23] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _21055_ (.RESET_B(net5361),
    .D(_00818_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[0] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _21056_ (.RESET_B(net5361),
    .D(_00819_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[1] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _21057_ (.RESET_B(net5331),
    .D(_00820_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[2] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _21058_ (.RESET_B(net5379),
    .D(_00821_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[4] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _21059_ (.RESET_B(net68),
    .D(_00822_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _21060_ (.RESET_B(net67),
    .D(_00823_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _21061_ (.RESET_B(net5361),
    .D(_00824_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[0] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _21062_ (.RESET_B(net5364),
    .D(_00825_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[1] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _21063_ (.RESET_B(net5331),
    .D(_00826_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[2] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _21064_ (.RESET_B(net5330),
    .D(_00827_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[3] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _21065_ (.RESET_B(net5364),
    .D(net760),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[4] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _21066_ (.RESET_B(net5220),
    .D(net2900),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _21067_ (.RESET_B(net5225),
    .D(net2869),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _21068_ (.RESET_B(net5225),
    .D(net2949),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _21069_ (.RESET_B(net5225),
    .D(net2374),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _21070_ (.RESET_B(net5201),
    .D(net461),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _21071_ (.RESET_B(net5202),
    .D(_00834_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _21072_ (.RESET_B(net5202),
    .D(net402),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _21073_ (.RESET_B(net5202),
    .D(net398),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[3] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _21074_ (.RESET_B(net5196),
    .D(net218),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[4] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _21075_ (.RESET_B(net5195),
    .D(net246),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[5] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21076_ (.RESET_B(net5195),
    .D(_00839_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _21077_ (.RESET_B(net5195),
    .D(net419),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21078_ (.RESET_B(net5197),
    .D(net369),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _21079_ (.RESET_B(net5197),
    .D(net304),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21080_ (.RESET_B(net5197),
    .D(_00843_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21081_ (.RESET_B(net5197),
    .D(net145),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[11] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21082_ (.RESET_B(net5226),
    .D(net335),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.flash_in_cont_mode ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _21083_ (.RESET_B(net5214),
    .D(_00846_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _21084_ (.RESET_B(net5284),
    .D(_00847_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _21085_ (.RESET_B(net5277),
    .D(_00848_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _21086_ (.RESET_B(net5275),
    .D(_00849_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21087_ (.RESET_B(net5264),
    .D(_00850_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21088_ (.RESET_B(net5277),
    .D(_00851_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _21089_ (.RESET_B(net5277),
    .D(net2821),
    .Q(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _21090_ (.RESET_B(net5264),
    .D(net2715),
    .Q(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21091_ (.RESET_B(net5275),
    .D(_00854_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21092_ (.RESET_B(net5277),
    .D(_00855_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _21093_ (.RESET_B(net5277),
    .D(net2670),
    .Q(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _21094_ (.RESET_B(net5275),
    .D(net2657),
    .Q(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _21095_ (.RESET_B(net5214),
    .D(_00858_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _21096_ (.RESET_B(net5284),
    .D(_00859_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _21097_ (.RESET_B(net5264),
    .D(net2812),
    .Q(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21098_ (.RESET_B(net5264),
    .D(net2694),
    .Q(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21099_ (.RESET_B(net5275),
    .D(net2678),
    .Q(\soc_inst.mem_ctrl.spi_data_out[16] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21100_ (.RESET_B(net5285),
    .D(_00863_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[17] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _21101_ (.RESET_B(net5278),
    .D(_00864_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _21102_ (.RESET_B(net5282),
    .D(net2882),
    .Q(\soc_inst.mem_ctrl.spi_data_out[19] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _21103_ (.RESET_B(net5282),
    .D(net2849),
    .Q(\soc_inst.mem_ctrl.spi_data_out[20] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _21104_ (.RESET_B(net5285),
    .D(_00867_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[21] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _21105_ (.RESET_B(net5284),
    .D(_00868_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[22] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _21106_ (.RESET_B(net5275),
    .D(net2667),
    .Q(\soc_inst.mem_ctrl.spi_data_out[23] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _21107_ (.RESET_B(net5282),
    .D(_00870_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[24] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _21108_ (.RESET_B(net5284),
    .D(net2642),
    .Q(\soc_inst.mem_ctrl.spi_data_out[25] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _21109_ (.RESET_B(net5279),
    .D(net2073),
    .Q(\soc_inst.mem_ctrl.spi_data_out[26] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _21110_ (.RESET_B(net5278),
    .D(net2842),
    .Q(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _21111_ (.RESET_B(net5277),
    .D(net2616),
    .Q(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _21112_ (.RESET_B(net5279),
    .D(net2464),
    .Q(\soc_inst.mem_ctrl.spi_data_out[29] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _21113_ (.RESET_B(net5285),
    .D(net2001),
    .Q(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _21114_ (.RESET_B(net5279),
    .D(net2098),
    .Q(\soc_inst.mem_ctrl.spi_data_out[31] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _21115_ (.RESET_B(net5474),
    .D(net79),
    .Q(\soc_inst.cpu_core.csr_file.mip_eip ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _21116_ (.RESET_B(net5322),
    .D(_00878_),
    .Q(\soc_inst.cpu_core.id_int_is_interrupt ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _21117_ (.RESET_B(net5357),
    .D(net617),
    .Q(\soc_inst.cpu_core.ex_reg_we ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _21118_ (.RESET_B(net5322),
    .D(_00880_),
    .Q(\soc_inst.cpu_core.csr_file.mret_trigger ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _21119_ (.RESET_B(net5323),
    .D(_00881_),
    .Q(\soc_inst.cpu_core.ex_is_ebreak ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _21120_ (.RESET_B(net5369),
    .D(_00882_),
    .Q(\soc_inst.core_mem_wdata[0] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _21121_ (.RESET_B(net5305),
    .D(net897),
    .Q(\soc_inst.core_mem_wdata[1] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _21122_ (.RESET_B(net5371),
    .D(net1266),
    .Q(\soc_inst.core_mem_wdata[2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _21123_ (.RESET_B(net5369),
    .D(net784),
    .Q(\soc_inst.core_mem_wdata[3] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _21124_ (.RESET_B(net5369),
    .D(_00886_),
    .Q(\soc_inst.core_mem_wdata[4] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _21125_ (.RESET_B(net5301),
    .D(_00887_),
    .Q(\soc_inst.core_mem_wdata[5] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _21126_ (.RESET_B(net5370),
    .D(net1148),
    .Q(\soc_inst.core_mem_wdata[6] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _21127_ (.RESET_B(net5367),
    .D(_00889_),
    .Q(\soc_inst.core_mem_wdata[7] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _21128_ (.RESET_B(net5389),
    .D(_00890_),
    .Q(\soc_inst.core_mem_wdata[8] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _21129_ (.RESET_B(net5370),
    .D(_00891_),
    .Q(\soc_inst.core_mem_wdata[9] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _21130_ (.RESET_B(net5389),
    .D(_00892_),
    .Q(\soc_inst.core_mem_wdata[10] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _21131_ (.RESET_B(net5370),
    .D(_00893_),
    .Q(\soc_inst.core_mem_wdata[11] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _21132_ (.RESET_B(net5370),
    .D(net1103),
    .Q(\soc_inst.core_mem_wdata[12] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _21133_ (.RESET_B(net5313),
    .D(net2163),
    .Q(\soc_inst.core_mem_wdata[13] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _21134_ (.RESET_B(net5325),
    .D(net1294),
    .Q(\soc_inst.core_mem_wdata[14] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _21135_ (.RESET_B(net5369),
    .D(_00897_),
    .Q(\soc_inst.core_mem_wdata[15] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _21136_ (.RESET_B(net5402),
    .D(net1067),
    .Q(\soc_inst.core_mem_wdata[16] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _21137_ (.RESET_B(net5403),
    .D(net2871),
    .Q(\soc_inst.core_mem_wdata[17] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _21138_ (.RESET_B(net5404),
    .D(_00900_),
    .Q(\soc_inst.core_mem_wdata[18] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _21139_ (.RESET_B(net5442),
    .D(_00901_),
    .Q(\soc_inst.core_mem_wdata[19] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _21140_ (.RESET_B(net5403),
    .D(net2852),
    .Q(\soc_inst.core_mem_wdata[20] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _21141_ (.RESET_B(net5402),
    .D(net1175),
    .Q(\soc_inst.core_mem_wdata[21] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _21142_ (.RESET_B(net5442),
    .D(net2755),
    .Q(\soc_inst.core_mem_wdata[22] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _21143_ (.RESET_B(net5403),
    .D(_00905_),
    .Q(\soc_inst.core_mem_wdata[23] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _21144_ (.RESET_B(net5370),
    .D(_00906_),
    .Q(\soc_inst.core_mem_wdata[24] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _21145_ (.RESET_B(net5372),
    .D(net1173),
    .Q(\soc_inst.core_mem_wdata[25] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _21146_ (.RESET_B(net5442),
    .D(_00908_),
    .Q(\soc_inst.core_mem_wdata[26] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _21147_ (.RESET_B(net5386),
    .D(_00909_),
    .Q(\soc_inst.core_mem_wdata[27] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _21148_ (.RESET_B(net5450),
    .D(_00910_),
    .Q(\soc_inst.core_mem_wdata[28] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _21149_ (.RESET_B(net5357),
    .D(net714),
    .Q(\soc_inst.core_mem_wdata[29] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _21150_ (.RESET_B(net5384),
    .D(_00912_),
    .Q(\soc_inst.core_mem_wdata[30] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _21151_ (.RESET_B(net5442),
    .D(_00913_),
    .Q(\soc_inst.core_mem_wdata[31] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _21152_ (.RESET_B(net5322),
    .D(net575),
    .Q(\soc_inst.cpu_core.ex_is_ecall ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _21153_ (.RESET_B(net5280),
    .D(_00915_),
    .Q(\soc_inst.cpu_core.error_flag_reg ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21154_ (.RESET_B(net5300),
    .D(_00916_),
    .Q(_00264_),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _21155_ (.RESET_B(net5300),
    .D(_00917_),
    .Q(_00265_),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _21156_ (.RESET_B(net5293),
    .D(_00918_),
    .Q(\soc_inst.cpu_core.if_instr[2] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _21157_ (.RESET_B(net5293),
    .D(_00919_),
    .Q(\soc_inst.cpu_core.if_instr[3] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21158_ (.RESET_B(net5293),
    .D(_00920_),
    .Q(_00266_),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21159_ (.RESET_B(net5292),
    .D(_00921_),
    .Q(\soc_inst.cpu_core.if_instr[5] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21160_ (.RESET_B(net5293),
    .D(_00922_),
    .Q(\soc_inst.cpu_core.if_instr[6] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21161_ (.RESET_B(net5288),
    .D(_00923_),
    .Q(\soc_inst.cpu_core.if_instr[7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _21162_ (.RESET_B(net5292),
    .D(_00924_),
    .Q(\soc_inst.cpu_core.if_instr[8] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _21163_ (.RESET_B(net5292),
    .D(_00925_),
    .Q(\soc_inst.cpu_core.if_instr[9] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21164_ (.RESET_B(net5292),
    .D(net668),
    .Q(\soc_inst.cpu_core.if_instr[10] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _21165_ (.RESET_B(net5293),
    .D(_00927_),
    .Q(\soc_inst.cpu_core.if_instr[11] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21166_ (.RESET_B(net5256),
    .D(_00928_),
    .Q(\soc_inst.cpu_core.if_funct3[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21167_ (.RESET_B(net5288),
    .D(_00929_),
    .Q(\soc_inst.cpu_core.if_funct3[1] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21168_ (.RESET_B(net5256),
    .D(_00930_),
    .Q(\soc_inst.cpu_core.if_funct3[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21169_ (.RESET_B(net5255),
    .D(_00931_),
    .Q(\soc_inst.cpu_core.if_instr[15] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _21170_ (.RESET_B(net5268),
    .D(_00932_),
    .Q(\soc_inst.cpu_core.if_instr[16] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _21171_ (.RESET_B(net5273),
    .D(_00933_),
    .Q(\soc_inst.cpu_core.if_instr[17] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _21172_ (.RESET_B(net5292),
    .D(_00934_),
    .Q(\soc_inst.cpu_core.if_instr[18] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21173_ (.RESET_B(net5289),
    .D(_00935_),
    .Q(\soc_inst.cpu_core.if_instr[19] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21174_ (.RESET_B(net5293),
    .D(_00936_),
    .Q(\soc_inst.cpu_core.if_imm12[0] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _21175_ (.RESET_B(net5268),
    .D(_00937_),
    .Q(\soc_inst.cpu_core.if_imm12[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _21176_ (.RESET_B(net5268),
    .D(_00938_),
    .Q(\soc_inst.cpu_core.if_imm12[2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21177_ (.RESET_B(net5290),
    .D(_00939_),
    .Q(\soc_inst.cpu_core.if_imm12[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21178_ (.RESET_B(net5272),
    .D(_00940_),
    .Q(\soc_inst.cpu_core.if_imm12[4] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _21179_ (.RESET_B(net5289),
    .D(_00941_),
    .Q(\soc_inst.cpu_core.if_funct7[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21180_ (.RESET_B(net5273),
    .D(_00942_),
    .Q(\soc_inst.cpu_core.if_funct7[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21181_ (.RESET_B(net5288),
    .D(_00943_),
    .Q(\soc_inst.cpu_core.if_funct7[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21182_ (.RESET_B(net5272),
    .D(_00944_),
    .Q(\soc_inst.cpu_core.if_funct7[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _21183_ (.RESET_B(net5300),
    .D(_00945_),
    .Q(\soc_inst.cpu_core.if_funct7[4] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _21184_ (.RESET_B(net5272),
    .D(_00946_),
    .Q(\soc_inst.cpu_core.if_funct7[5] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _21185_ (.RESET_B(net5268),
    .D(_00947_),
    .Q(\soc_inst.cpu_core.if_funct7[6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _21186_ (.RESET_B(net5373),
    .D(_00948_),
    .Q(\soc_inst.cpu_core.if_pc[0] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _21187_ (.RESET_B(net5372),
    .D(net2136),
    .Q(\soc_inst.cpu_core.if_pc[1] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _21188_ (.RESET_B(net5372),
    .D(net979),
    .Q(\soc_inst.cpu_core.if_pc[2] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _21189_ (.RESET_B(net5372),
    .D(net2035),
    .Q(\soc_inst.cpu_core.if_pc[3] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _21190_ (.RESET_B(net5362),
    .D(net2403),
    .Q(\soc_inst.cpu_core.if_pc[4] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _21191_ (.RESET_B(net5362),
    .D(net2288),
    .Q(\soc_inst.cpu_core.if_pc[5] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _21192_ (.RESET_B(net5362),
    .D(net2316),
    .Q(\soc_inst.cpu_core.if_pc[6] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _21193_ (.RESET_B(net5363),
    .D(net2230),
    .Q(\soc_inst.cpu_core.if_pc[7] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _21194_ (.RESET_B(net5326),
    .D(net2031),
    .Q(\soc_inst.cpu_core.if_pc[8] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21195_ (.RESET_B(net5327),
    .D(net2286),
    .Q(\soc_inst.cpu_core.if_pc[9] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _21196_ (.RESET_B(net5327),
    .D(net2033),
    .Q(\soc_inst.cpu_core.if_pc[10] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21197_ (.RESET_B(net5326),
    .D(net1899),
    .Q(\soc_inst.cpu_core.if_pc[11] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21198_ (.RESET_B(net5326),
    .D(net1989),
    .Q(\soc_inst.cpu_core.if_pc[12] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _21199_ (.RESET_B(net5322),
    .D(net1817),
    .Q(\soc_inst.cpu_core.if_pc[13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _21200_ (.RESET_B(net5324),
    .D(net1976),
    .Q(\soc_inst.cpu_core.if_pc[14] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _21201_ (.RESET_B(net5324),
    .D(net1947),
    .Q(\soc_inst.cpu_core.if_pc[15] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _21202_ (.RESET_B(net5309),
    .D(net1722),
    .Q(\soc_inst.cpu_core.if_pc[16] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _21203_ (.RESET_B(net5311),
    .D(net2369),
    .Q(\soc_inst.cpu_core.if_pc[17] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _21204_ (.RESET_B(net5247),
    .D(net2344),
    .Q(\soc_inst.cpu_core.if_pc[18] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _21205_ (.RESET_B(net5247),
    .D(net2027),
    .Q(\soc_inst.cpu_core.if_pc[19] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _21206_ (.RESET_B(net5311),
    .D(net1872),
    .Q(\soc_inst.cpu_core.if_pc[20] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _21207_ (.RESET_B(net5309),
    .D(net1742),
    .Q(\soc_inst.cpu_core.if_pc[21] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _21208_ (.RESET_B(net5309),
    .D(net2007),
    .Q(\soc_inst.cpu_core.if_pc[22] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _21209_ (.RESET_B(net5309),
    .D(net2165),
    .Q(\soc_inst.cpu_core.if_pc[23] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _21210_ (.RESET_B(net5374),
    .D(_00026_),
    .Q(\soc_inst.cpu_core.mem_stall ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _21211_ (.RESET_B(net5292),
    .D(_00972_),
    .Q(\soc_inst.cpu_core.if_is_compressed ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _21212_ (.RESET_B(net5370),
    .D(_00973_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[0] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _21213_ (.RESET_B(net5256),
    .D(net809),
    .Q(\soc_inst.cpu_core.mem_rs1_data[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _21214_ (.RESET_B(net5367),
    .D(_00975_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[2] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _21215_ (.RESET_B(net5372),
    .D(net775),
    .Q(\soc_inst.cpu_core.mem_rs1_data[3] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _21216_ (.RESET_B(net5357),
    .D(_00977_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[4] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _21217_ (.RESET_B(net5299),
    .D(_00978_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _21218_ (.RESET_B(net5300),
    .D(_00979_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _21219_ (.RESET_B(net5299),
    .D(_00980_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _21220_ (.RESET_B(net5295),
    .D(_00981_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21221_ (.RESET_B(net5346),
    .D(_00982_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _21222_ (.RESET_B(net5378),
    .D(net2457),
    .Q(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _21223_ (.RESET_B(net5325),
    .D(net638),
    .Q(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _21224_ (.RESET_B(net5323),
    .D(_00985_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _21225_ (.RESET_B(net5258),
    .D(_00986_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _21226_ (.RESET_B(net5322),
    .D(_00987_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _21227_ (.RESET_B(net5323),
    .D(_00988_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _21228_ (.RESET_B(net5310),
    .D(net1138),
    .Q(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _21229_ (.RESET_B(net5309),
    .D(net2224),
    .Q(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _21230_ (.RESET_B(net5315),
    .D(_00991_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _21231_ (.RESET_B(net5317),
    .D(_00992_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _21232_ (.RESET_B(net5310),
    .D(_00993_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _21233_ (.RESET_B(net5317),
    .D(_00994_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _21234_ (.RESET_B(net5317),
    .D(_00995_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _21235_ (.RESET_B(net5315),
    .D(_00996_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _21236_ (.RESET_B(net5348),
    .D(net1257),
    .Q(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _21237_ (.RESET_B(net5403),
    .D(_00998_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[25] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _21238_ (.RESET_B(net5350),
    .D(_00999_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _21239_ (.RESET_B(net5342),
    .D(net935),
    .Q(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _21240_ (.RESET_B(net5402),
    .D(net917),
    .Q(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _21241_ (.RESET_B(net5406),
    .D(_01002_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[29] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _21242_ (.RESET_B(net5341),
    .D(_01003_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _21243_ (.RESET_B(net5350),
    .D(_01004_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _21244_ (.RESET_B(net5366),
    .D(_01005_),
    .Q(_00267_),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _21245_ (.RESET_B(net5366),
    .D(_01006_),
    .Q(_00268_),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _21246_ (.RESET_B(net5296),
    .D(_01007_),
    .Q(\soc_inst.cpu_core.id_instr[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21247_ (.RESET_B(net5299),
    .D(_01008_),
    .Q(\soc_inst.cpu_core.id_instr[3] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _21248_ (.RESET_B(net5299),
    .D(_01009_),
    .Q(_00269_),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _21249_ (.RESET_B(net5297),
    .D(_01010_),
    .Q(\soc_inst.cpu_core.id_instr[5] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _21250_ (.RESET_B(net5297),
    .D(_01011_),
    .Q(\soc_inst.cpu_core.id_instr[6] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _21251_ (.RESET_B(net5268),
    .D(_01012_),
    .Q(\soc_inst.cpu_core.id_instr[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _21252_ (.RESET_B(net5289),
    .D(_01013_),
    .Q(\soc_inst.cpu_core.id_instr[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _21253_ (.RESET_B(net5289),
    .D(_01014_),
    .Q(\soc_inst.cpu_core.id_instr[9] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _21254_ (.RESET_B(net5289),
    .D(_01015_),
    .Q(\soc_inst.cpu_core.id_instr[10] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21255_ (.RESET_B(net5290),
    .D(_01016_),
    .Q(\soc_inst.cpu_core.id_instr[11] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21256_ (.RESET_B(net5256),
    .D(_01017_),
    .Q(\soc_inst.cpu_core.id_funct3[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _21257_ (.RESET_B(net5255),
    .D(_01018_),
    .Q(\soc_inst.cpu_core.id_funct3[1] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _21258_ (.RESET_B(net5256),
    .D(_01019_),
    .Q(\soc_inst.cpu_core.id_funct3[2] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _21259_ (.RESET_B(net5296),
    .D(_01020_),
    .Q(\soc_inst.cpu_core.id_instr[15] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21260_ (.RESET_B(net5233),
    .D(_01021_),
    .Q(\soc_inst.cpu_core.id_instr[16] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _21261_ (.RESET_B(net5244),
    .D(_01022_),
    .Q(\soc_inst.cpu_core.id_instr[17] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _21262_ (.RESET_B(net5246),
    .D(_01023_),
    .Q(\soc_inst.cpu_core.id_instr[18] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _21263_ (.RESET_B(net5245),
    .D(_01024_),
    .Q(\soc_inst.cpu_core.id_instr[19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _21264_ (.RESET_B(net5244),
    .D(_01025_),
    .Q(\soc_inst.cpu_core.id_imm12[0] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21265_ (.RESET_B(net5245),
    .D(_01026_),
    .Q(\soc_inst.cpu_core.id_imm12[1] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _21266_ (.RESET_B(net5251),
    .D(_01027_),
    .Q(\soc_inst.cpu_core.id_imm12[2] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _21267_ (.RESET_B(net5245),
    .D(_01028_),
    .Q(\soc_inst.cpu_core.id_imm12[3] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _21268_ (.RESET_B(net5254),
    .D(_01029_),
    .Q(\soc_inst.cpu_core.id_imm12[4] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _21269_ (.RESET_B(net5257),
    .D(_01030_),
    .Q(\soc_inst.cpu_core.id_imm12[5] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _21270_ (.RESET_B(net5253),
    .D(_01031_),
    .Q(\soc_inst.cpu_core.id_imm12[6] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21271_ (.RESET_B(net5254),
    .D(_01032_),
    .Q(\soc_inst.cpu_core.id_imm12[7] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21272_ (.RESET_B(net5253),
    .D(_01033_),
    .Q(\soc_inst.cpu_core.id_imm12[8] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21273_ (.RESET_B(net5250),
    .D(_01034_),
    .Q(\soc_inst.cpu_core.id_imm12[9] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _21274_ (.RESET_B(net5323),
    .D(_01035_),
    .Q(\soc_inst.cpu_core.id_imm12[10] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _21275_ (.RESET_B(net5259),
    .D(_01036_),
    .Q(\soc_inst.cpu_core.id_imm12[11] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _21276_ (.RESET_B(net5421),
    .D(_00169_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _21277_ (.RESET_B(net5421),
    .D(_00180_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _21278_ (.RESET_B(net5421),
    .D(_00191_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _21279_ (.RESET_B(net5421),
    .D(net968),
    .Q(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _21280_ (.RESET_B(net5445),
    .D(net1661),
    .Q(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _21281_ (.RESET_B(net5445),
    .D(_00212_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _21282_ (.RESET_B(net5445),
    .D(net827),
    .Q(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _21283_ (.RESET_B(net5422),
    .D(net1263),
    .Q(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _21284_ (.RESET_B(net5414),
    .D(net885),
    .Q(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _21285_ (.RESET_B(net5414),
    .D(net2887),
    .Q(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _21286_ (.RESET_B(net5413),
    .D(net646),
    .Q(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _21287_ (.RESET_B(net5406),
    .D(net1169),
    .Q(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _21288_ (.RESET_B(net5404),
    .D(_00172_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _21289_ (.RESET_B(net5409),
    .D(net1612),
    .Q(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _21290_ (.RESET_B(net5409),
    .D(_00174_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _21291_ (.RESET_B(net5409),
    .D(_00175_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _21292_ (.RESET_B(net5402),
    .D(net2425),
    .Q(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _21293_ (.RESET_B(net5402),
    .D(net2439),
    .Q(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _21294_ (.RESET_B(net5401),
    .D(net2127),
    .Q(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _21295_ (.RESET_B(net5401),
    .D(_00179_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _21296_ (.RESET_B(net5401),
    .D(net2420),
    .Q(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _21297_ (.RESET_B(net5401),
    .D(_00182_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _21298_ (.RESET_B(net5401),
    .D(net1528),
    .Q(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _21299_ (.RESET_B(net5401),
    .D(net2542),
    .Q(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _21300_ (.RESET_B(net5403),
    .D(net2228),
    .Q(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _21301_ (.RESET_B(net5405),
    .D(net2220),
    .Q(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _21302_ (.RESET_B(net5413),
    .D(net1657),
    .Q(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _21303_ (.RESET_B(net5405),
    .D(_00188_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _21304_ (.RESET_B(net5413),
    .D(net1773),
    .Q(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _21305_ (.RESET_B(net5416),
    .D(_00190_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _21306_ (.RESET_B(net5416),
    .D(net2050),
    .Q(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _21307_ (.RESET_B(net5413),
    .D(net1901),
    .Q(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _21308_ (.RESET_B(net5420),
    .D(_00194_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _21309_ (.RESET_B(net5420),
    .D(net1894),
    .Q(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _21310_ (.RESET_B(net5420),
    .D(net2588),
    .Q(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _21311_ (.RESET_B(net5420),
    .D(net1245),
    .Q(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _21312_ (.RESET_B(net5422),
    .D(net1716),
    .Q(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _21313_ (.RESET_B(net5422),
    .D(_00199_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _21314_ (.RESET_B(net5422),
    .D(net794),
    .Q(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _21315_ (.RESET_B(net5418),
    .D(net1654),
    .Q(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _21316_ (.RESET_B(net5418),
    .D(_00203_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _21317_ (.RESET_B(net5418),
    .D(_00204_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _21318_ (.RESET_B(net5418),
    .D(net725),
    .Q(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _21319_ (.RESET_B(net5410),
    .D(_00206_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _21320_ (.RESET_B(net5410),
    .D(net1094),
    .Q(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _21321_ (.RESET_B(net5410),
    .D(_00208_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _21322_ (.RESET_B(net5410),
    .D(_00209_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _21323_ (.RESET_B(net5410),
    .D(net695),
    .Q(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _21324_ (.RESET_B(net5264),
    .D(_01037_),
    .Q(\soc_inst.cpu_core.id_rs1_data[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21325_ (.RESET_B(net5264),
    .D(_01038_),
    .Q(\soc_inst.cpu_core.id_rs1_data[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21326_ (.RESET_B(net5270),
    .D(_01039_),
    .Q(\soc_inst.cpu_core.id_rs1_data[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21327_ (.RESET_B(net5265),
    .D(_01040_),
    .Q(\soc_inst.cpu_core.id_rs1_data[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21328_ (.RESET_B(net5265),
    .D(_01041_),
    .Q(\soc_inst.cpu_core.id_rs1_data[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21329_ (.RESET_B(net5264),
    .D(_01042_),
    .Q(\soc_inst.cpu_core.id_rs1_data[5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _21330_ (.RESET_B(net5270),
    .D(_01043_),
    .Q(\soc_inst.cpu_core.id_rs1_data[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21331_ (.RESET_B(net5264),
    .D(_01044_),
    .Q(\soc_inst.cpu_core.id_rs1_data[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _21332_ (.RESET_B(net5267),
    .D(_01045_),
    .Q(\soc_inst.cpu_core.id_rs1_data[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21333_ (.RESET_B(net5267),
    .D(_01046_),
    .Q(\soc_inst.cpu_core.id_rs1_data[9] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21334_ (.RESET_B(net5267),
    .D(_01047_),
    .Q(\soc_inst.cpu_core.id_rs1_data[10] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _21335_ (.RESET_B(net5267),
    .D(_01048_),
    .Q(\soc_inst.cpu_core.id_rs1_data[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21336_ (.RESET_B(net5265),
    .D(_01049_),
    .Q(\soc_inst.cpu_core.id_rs1_data[12] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21337_ (.RESET_B(net5172),
    .D(_01050_),
    .Q(\soc_inst.cpu_core.id_rs1_data[13] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _21338_ (.RESET_B(net5255),
    .D(_01051_),
    .Q(\soc_inst.cpu_core.id_rs1_data[14] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21339_ (.RESET_B(net5253),
    .D(_01052_),
    .Q(\soc_inst.cpu_core.id_rs1_data[15] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21340_ (.RESET_B(net5231),
    .D(_01053_),
    .Q(\soc_inst.cpu_core.id_rs1_data[16] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21341_ (.RESET_B(net5243),
    .D(_01054_),
    .Q(\soc_inst.cpu_core.id_rs1_data[17] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21342_ (.RESET_B(net5165),
    .D(_01055_),
    .Q(\soc_inst.cpu_core.id_rs1_data[18] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _21343_ (.RESET_B(net5231),
    .D(_01056_),
    .Q(\soc_inst.cpu_core.id_rs1_data[19] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21344_ (.RESET_B(net5230),
    .D(_01057_),
    .Q(\soc_inst.cpu_core.id_rs1_data[20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21345_ (.RESET_B(net5241),
    .D(_01058_),
    .Q(\soc_inst.cpu_core.id_rs1_data[21] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21346_ (.RESET_B(net5165),
    .D(_01059_),
    .Q(\soc_inst.cpu_core.id_rs1_data[22] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _21347_ (.RESET_B(net5229),
    .D(_01060_),
    .Q(\soc_inst.cpu_core.id_rs1_data[23] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21348_ (.RESET_B(net5237),
    .D(_01061_),
    .Q(\soc_inst.cpu_core.id_rs1_data[24] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21349_ (.RESET_B(net5269),
    .D(_01062_),
    .Q(\soc_inst.cpu_core.id_rs1_data[25] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21350_ (.RESET_B(net5262),
    .D(_01063_),
    .Q(\soc_inst.cpu_core.id_rs1_data[26] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _21351_ (.RESET_B(net5172),
    .D(_01064_),
    .Q(\soc_inst.cpu_core.id_rs1_data[27] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _21352_ (.RESET_B(net5230),
    .D(_01065_),
    .Q(\soc_inst.cpu_core.id_rs1_data[28] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21353_ (.RESET_B(net5240),
    .D(_01066_),
    .Q(\soc_inst.cpu_core.id_rs1_data[29] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21354_ (.RESET_B(net5267),
    .D(_01067_),
    .Q(\soc_inst.cpu_core.id_rs1_data[30] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21355_ (.RESET_B(net5267),
    .D(_01068_),
    .Q(\soc_inst.cpu_core.id_rs1_data[31] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _21356_ (.RESET_B(net5362),
    .D(net850),
    .Q(_00270_),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _21357_ (.RESET_B(net5358),
    .D(net1286),
    .Q(_00271_),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _21358_ (.RESET_B(net5362),
    .D(net197),
    .Q(\soc_inst.cpu_core.mem_instr[2] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _21359_ (.RESET_B(net5358),
    .D(net822),
    .Q(\soc_inst.cpu_core.mem_instr[3] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _21360_ (.RESET_B(net5373),
    .D(net604),
    .Q(_00272_),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _21361_ (.RESET_B(net5365),
    .D(net587),
    .Q(\soc_inst.cpu_core.mem_instr[5] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21362_ (.RESET_B(net5373),
    .D(net2188),
    .Q(\soc_inst.cpu_core.mem_instr[6] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _21363_ (.RESET_B(net5288),
    .D(_01076_),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _21364_ (.RESET_B(net5331),
    .D(_01077_),
    .Q(\soc_inst.core_mem_flag[0] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _21365_ (.RESET_B(net5329),
    .D(_01078_),
    .Q(\soc_inst.core_mem_flag[1] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _21366_ (.RESET_B(net5330),
    .D(_01079_),
    .Q(\soc_inst.core_mem_flag[2] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _21367_ (.RESET_B(net5363),
    .D(net811),
    .Q(\soc_inst.cpu_core.mem_instr[15] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _21368_ (.RESET_B(net5312),
    .D(net2131),
    .Q(\soc_inst.cpu_core.mem_instr[16] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _21369_ (.RESET_B(net5319),
    .D(net1883),
    .Q(\soc_inst.cpu_core.mem_instr[17] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _21370_ (.RESET_B(net5319),
    .D(_01083_),
    .Q(\soc_inst.cpu_core.mem_instr[18] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _21371_ (.RESET_B(net5358),
    .D(net1075),
    .Q(\soc_inst.cpu_core.mem_instr[19] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _21372_ (.RESET_B(net5336),
    .D(_01085_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _21373_ (.RESET_B(net5336),
    .D(_01086_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _21374_ (.RESET_B(net5343),
    .D(net1810),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _21375_ (.RESET_B(net5319),
    .D(net856),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _21376_ (.RESET_B(net5337),
    .D(_01089_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _21377_ (.RESET_B(net5312),
    .D(net743),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _21378_ (.RESET_B(net5323),
    .D(net2068),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _21379_ (.RESET_B(net5250),
    .D(_01092_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _21380_ (.RESET_B(net5320),
    .D(_01093_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _21381_ (.RESET_B(net5319),
    .D(net425),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _21382_ (.RESET_B(net5328),
    .D(net449),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _21383_ (.RESET_B(net5328),
    .D(net2046),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _21384_ (.RESET_B(net5292),
    .D(_01097_),
    .Q(\soc_inst.cpu_core.id_rs2_data[0] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _21385_ (.RESET_B(net5265),
    .D(_01098_),
    .Q(\soc_inst.cpu_core.id_rs2_data[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21386_ (.RESET_B(net5292),
    .D(_01099_),
    .Q(\soc_inst.cpu_core.id_rs2_data[2] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _21387_ (.RESET_B(net5277),
    .D(_01100_),
    .Q(\soc_inst.cpu_core.id_rs2_data[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21388_ (.RESET_B(net5300),
    .D(_01101_),
    .Q(\soc_inst.cpu_core.id_rs2_data[4] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _21389_ (.RESET_B(net5296),
    .D(_01102_),
    .Q(\soc_inst.cpu_core.id_rs2_data[5] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _21390_ (.RESET_B(net5275),
    .D(_01103_),
    .Q(\soc_inst.cpu_core.id_rs2_data[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21391_ (.RESET_B(net5277),
    .D(_01104_),
    .Q(\soc_inst.cpu_core.id_rs2_data[7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _21392_ (.RESET_B(net5255),
    .D(_01105_),
    .Q(\soc_inst.cpu_core.id_rs2_data[8] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _21393_ (.RESET_B(net5270),
    .D(_01106_),
    .Q(\soc_inst.cpu_core.id_rs2_data[9] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _21394_ (.RESET_B(net5269),
    .D(_01107_),
    .Q(\soc_inst.cpu_core.id_rs2_data[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21395_ (.RESET_B(net5267),
    .D(_01108_),
    .Q(\soc_inst.cpu_core.id_rs2_data[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21396_ (.RESET_B(net5269),
    .D(_01109_),
    .Q(\soc_inst.cpu_core.id_rs2_data[12] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _21397_ (.RESET_B(net5254),
    .D(_01110_),
    .Q(\soc_inst.cpu_core.id_rs2_data[13] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21398_ (.RESET_B(net5263),
    .D(_01111_),
    .Q(\soc_inst.cpu_core.id_rs2_data[14] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21399_ (.RESET_B(net5240),
    .D(net2637),
    .Q(\soc_inst.cpu_core.id_rs2_data[15] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _21400_ (.RESET_B(net5242),
    .D(_01113_),
    .Q(\soc_inst.cpu_core.id_rs2_data[16] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21401_ (.RESET_B(net5242),
    .D(_01114_),
    .Q(\soc_inst.cpu_core.id_rs2_data[17] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21402_ (.RESET_B(net5243),
    .D(_01115_),
    .Q(\soc_inst.cpu_core.id_rs2_data[18] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21403_ (.RESET_B(net5230),
    .D(_01116_),
    .Q(\soc_inst.cpu_core.id_rs2_data[19] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _21404_ (.RESET_B(net5242),
    .D(_01117_),
    .Q(\soc_inst.cpu_core.id_rs2_data[20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21405_ (.RESET_B(net5243),
    .D(_01118_),
    .Q(\soc_inst.cpu_core.id_rs2_data[21] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21406_ (.RESET_B(net5242),
    .D(_01119_),
    .Q(\soc_inst.cpu_core.id_rs2_data[22] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _21407_ (.RESET_B(net5242),
    .D(_01120_),
    .Q(\soc_inst.cpu_core.id_rs2_data[23] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _21408_ (.RESET_B(net5254),
    .D(_01121_),
    .Q(\soc_inst.cpu_core.id_rs2_data[24] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21409_ (.RESET_B(net5237),
    .D(_01122_),
    .Q(\soc_inst.cpu_core.id_rs2_data[25] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21410_ (.RESET_B(net5237),
    .D(_01123_),
    .Q(\soc_inst.cpu_core.id_rs2_data[26] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21411_ (.RESET_B(net5236),
    .D(_01124_),
    .Q(\soc_inst.cpu_core.id_rs2_data[27] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21412_ (.RESET_B(net5233),
    .D(_01125_),
    .Q(\soc_inst.cpu_core.id_rs2_data[28] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _21413_ (.RESET_B(net5253),
    .D(_01126_),
    .Q(\soc_inst.cpu_core.id_rs2_data[29] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _21414_ (.RESET_B(net5239),
    .D(_01127_),
    .Q(\soc_inst.cpu_core.id_rs2_data[30] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _21415_ (.RESET_B(net5255),
    .D(_01128_),
    .Q(\soc_inst.cpu_core.id_rs2_data[31] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21416_ (.RESET_B(net5290),
    .D(_01129_),
    .Q(\soc_inst.cpu_core.id_imm[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _21417_ (.RESET_B(net5290),
    .D(net1916),
    .Q(\soc_inst.cpu_core.id_imm[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21418_ (.RESET_B(net5290),
    .D(_01131_),
    .Q(\soc_inst.cpu_core.id_imm[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21419_ (.RESET_B(net5294),
    .D(_01132_),
    .Q(\soc_inst.cpu_core.id_imm[3] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21420_ (.RESET_B(net5294),
    .D(net2020),
    .Q(\soc_inst.cpu_core.id_imm[4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21421_ (.RESET_B(net5295),
    .D(net2239),
    .Q(\soc_inst.cpu_core.id_imm[5] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _21422_ (.RESET_B(net5294),
    .D(_01135_),
    .Q(\soc_inst.cpu_core.id_imm[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21423_ (.RESET_B(net5291),
    .D(net2037),
    .Q(\soc_inst.cpu_core.id_imm[7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _21424_ (.RESET_B(net5290),
    .D(net1491),
    .Q(\soc_inst.cpu_core.id_imm[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _21425_ (.RESET_B(net5290),
    .D(net1582),
    .Q(\soc_inst.cpu_core.id_imm[9] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _21426_ (.RESET_B(net5256),
    .D(_01139_),
    .Q(\soc_inst.cpu_core.id_imm[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _21427_ (.RESET_B(net5268),
    .D(net1063),
    .Q(\soc_inst.cpu_core.id_imm[11] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21428_ (.RESET_B(net5256),
    .D(net1804),
    .Q(\soc_inst.cpu_core.id_imm[12] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _21429_ (.RESET_B(net5253),
    .D(_01142_),
    .Q(\soc_inst.cpu_core.id_imm[13] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21430_ (.RESET_B(net5237),
    .D(_01143_),
    .Q(\soc_inst.cpu_core.id_imm[14] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _21431_ (.RESET_B(net5253),
    .D(_01144_),
    .Q(\soc_inst.cpu_core.id_imm[15] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21432_ (.RESET_B(net5244),
    .D(net2190),
    .Q(\soc_inst.cpu_core.id_imm[16] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _21433_ (.RESET_B(net5242),
    .D(_01146_),
    .Q(\soc_inst.cpu_core.id_imm[17] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21434_ (.RESET_B(net5244),
    .D(net2090),
    .Q(\soc_inst.cpu_core.id_imm[18] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _21435_ (.RESET_B(net5242),
    .D(net1252),
    .Q(\soc_inst.cpu_core.id_imm[19] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21436_ (.RESET_B(net5230),
    .D(_01149_),
    .Q(\soc_inst.cpu_core.id_imm[20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21437_ (.RESET_B(net5230),
    .D(_01150_),
    .Q(\soc_inst.cpu_core.id_imm[21] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21438_ (.RESET_B(net5230),
    .D(_01151_),
    .Q(\soc_inst.cpu_core.id_imm[22] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21439_ (.RESET_B(net5230),
    .D(_01152_),
    .Q(\soc_inst.cpu_core.id_imm[23] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21440_ (.RESET_B(net5232),
    .D(_01153_),
    .Q(\soc_inst.cpu_core.id_imm[24] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21441_ (.RESET_B(net5233),
    .D(_01154_),
    .Q(\soc_inst.cpu_core.id_imm[25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21442_ (.RESET_B(net5236),
    .D(_01155_),
    .Q(\soc_inst.cpu_core.id_imm[26] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21443_ (.RESET_B(net5236),
    .D(_01156_),
    .Q(\soc_inst.cpu_core.id_imm[27] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21444_ (.RESET_B(net5233),
    .D(_01157_),
    .Q(\soc_inst.cpu_core.id_imm[28] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _21445_ (.RESET_B(net5236),
    .D(_01158_),
    .Q(\soc_inst.cpu_core.id_imm[29] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21446_ (.RESET_B(net5253),
    .D(_01159_),
    .Q(\soc_inst.cpu_core.id_imm[30] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21447_ (.RESET_B(net5255),
    .D(net994),
    .Q(\soc_inst.cpu_core.id_imm[31] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _21448_ (.RESET_B(net5355),
    .D(_01161_),
    .Q(\soc_inst.cpu_core.mem_reg_we ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _21449_ (.RESET_B(net5235),
    .D(_01162_),
    .Q(\soc_inst.cpu_core.alu.op[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _21450_ (.RESET_B(net5237),
    .D(_01163_),
    .Q(\soc_inst.cpu_core.alu.op[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21451_ (.RESET_B(net5237),
    .D(_01164_),
    .Q(\soc_inst.cpu_core.alu.op[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21452_ (.RESET_B(net5235),
    .D(_01165_),
    .Q(\soc_inst.cpu_core.alu.op[3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21453_ (.RESET_B(net5212),
    .D(_01166_),
    .Q(\soc_inst.cpu_core.alu.a[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21454_ (.RESET_B(net5262),
    .D(_01167_),
    .Q(\soc_inst.cpu_core.alu.a[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _21455_ (.RESET_B(net5269),
    .D(_01168_),
    .Q(\soc_inst.cpu_core.alu.a[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _21456_ (.RESET_B(net5265),
    .D(_01169_),
    .Q(\soc_inst.cpu_core.alu.a[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21457_ (.RESET_B(net5212),
    .D(_01170_),
    .Q(\soc_inst.cpu_core.alu.a[4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21458_ (.RESET_B(net5212),
    .D(_01171_),
    .Q(\soc_inst.cpu_core.alu.a[5] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _21459_ (.RESET_B(net5212),
    .D(net1923),
    .Q(\soc_inst.cpu_core.alu.a[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _21460_ (.RESET_B(net5214),
    .D(net1689),
    .Q(\soc_inst.cpu_core.alu.a[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _21461_ (.RESET_B(net5262),
    .D(_01174_),
    .Q(\soc_inst.cpu_core.alu.a[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _21462_ (.RESET_B(net5262),
    .D(_01175_),
    .Q(\soc_inst.cpu_core.alu.a[9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _21463_ (.RESET_B(net5240),
    .D(_01176_),
    .Q(\soc_inst.cpu_core.alu.a[10] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21464_ (.RESET_B(net5263),
    .D(_01177_),
    .Q(\soc_inst.cpu_core.alu.a[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21465_ (.RESET_B(net5238),
    .D(_01178_),
    .Q(\soc_inst.cpu_core.alu.a[12] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _21466_ (.RESET_B(net5172),
    .D(_01179_),
    .Q(\soc_inst.cpu_core.alu.a[13] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _21467_ (.RESET_B(net5232),
    .D(_01180_),
    .Q(\soc_inst.cpu_core.alu.a[14] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _21468_ (.RESET_B(net5232),
    .D(_01181_),
    .Q(\soc_inst.cpu_core.alu.a[15] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _21469_ (.RESET_B(net5229),
    .D(_01182_),
    .Q(\soc_inst.cpu_core.alu.a[16] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21470_ (.RESET_B(net5231),
    .D(_01183_),
    .Q(\soc_inst.cpu_core.alu.a[17] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21471_ (.RESET_B(net5165),
    .D(_01184_),
    .Q(\soc_inst.cpu_core.alu.a[18] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _21472_ (.RESET_B(net5229),
    .D(_01185_),
    .Q(\soc_inst.cpu_core.alu.a[19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _21473_ (.RESET_B(net5229),
    .D(_01186_),
    .Q(\soc_inst.cpu_core.alu.a[20] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _21474_ (.RESET_B(net5229),
    .D(_01187_),
    .Q(\soc_inst.cpu_core.alu.a[21] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_2 _21475_ (.RESET_B(net5165),
    .D(_01188_),
    .Q(\soc_inst.cpu_core.alu.a[22] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _21476_ (.RESET_B(net5229),
    .D(net1131),
    .Q(\soc_inst.cpu_core.alu.a[23] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _21477_ (.RESET_B(net5211),
    .D(_01190_),
    .Q(\soc_inst.cpu_core.alu.a[24] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _21478_ (.RESET_B(net5211),
    .D(_01191_),
    .Q(\soc_inst.cpu_core.alu.a[25] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _21479_ (.RESET_B(net5211),
    .D(_01192_),
    .Q(\soc_inst.cpu_core.alu.a[26] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _21480_ (.RESET_B(net5173),
    .D(_01193_),
    .Q(\soc_inst.cpu_core.alu.a[27] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _21481_ (.RESET_B(net5165),
    .D(_01194_),
    .Q(\soc_inst.cpu_core.alu.a[28] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _21482_ (.RESET_B(net5172),
    .D(_01195_),
    .Q(\soc_inst.cpu_core.alu.a[29] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _21483_ (.RESET_B(net5212),
    .D(_01196_),
    .Q(\soc_inst.cpu_core.alu.a[30] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _21484_ (.RESET_B(net5263),
    .D(_01197_),
    .Q(\soc_inst.cpu_core.alu.a[31] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _21485_ (.RESET_B(net5263),
    .D(_01198_),
    .Q(\soc_inst.cpu_core.alu.b[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _21486_ (.RESET_B(net5214),
    .D(_01199_),
    .Q(\soc_inst.cpu_core.alu.b[1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _21487_ (.RESET_B(net5268),
    .D(_01200_),
    .Q(\soc_inst.cpu_core.alu.b[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _21488_ (.RESET_B(net5238),
    .D(_01201_),
    .Q(\soc_inst.cpu_core.alu.b[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _21489_ (.RESET_B(net5263),
    .D(_01202_),
    .Q(\soc_inst.cpu_core.alu.b[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _21490_ (.RESET_B(net5262),
    .D(net1160),
    .Q(\soc_inst.cpu_core.alu.b[5] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _21491_ (.RESET_B(net5212),
    .D(net1387),
    .Q(\soc_inst.cpu_core.alu.b[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _21492_ (.RESET_B(net5212),
    .D(net1412),
    .Q(\soc_inst.cpu_core.alu.b[7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _21493_ (.RESET_B(net5240),
    .D(_01206_),
    .Q(\soc_inst.cpu_core.alu.b[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21494_ (.RESET_B(net5262),
    .D(_01207_),
    .Q(\soc_inst.cpu_core.alu.b[9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _21495_ (.RESET_B(net5240),
    .D(net1961),
    .Q(\soc_inst.cpu_core.alu.b[10] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21496_ (.RESET_B(net5267),
    .D(_01209_),
    .Q(\soc_inst.cpu_core.alu.b[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _21497_ (.RESET_B(net5235),
    .D(_01210_),
    .Q(\soc_inst.cpu_core.alu.b[12] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21498_ (.RESET_B(net5232),
    .D(_01211_),
    .Q(\soc_inst.cpu_core.alu.b[13] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _21499_ (.RESET_B(net5238),
    .D(_01212_),
    .Q(\soc_inst.cpu_core.alu.b[14] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _21500_ (.RESET_B(net5232),
    .D(_01213_),
    .Q(\soc_inst.cpu_core.alu.b[15] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _21501_ (.RESET_B(net5229),
    .D(_01214_),
    .Q(\soc_inst.cpu_core.alu.b[16] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _21502_ (.RESET_B(net5231),
    .D(_01215_),
    .Q(\soc_inst.cpu_core.alu.b[17] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21503_ (.RESET_B(net5230),
    .D(_01216_),
    .Q(\soc_inst.cpu_core.alu.b[18] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _21504_ (.RESET_B(net5231),
    .D(net2618),
    .Q(\soc_inst.cpu_core.alu.b[19] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21505_ (.RESET_B(net5231),
    .D(_01218_),
    .Q(\soc_inst.cpu_core.alu.b[20] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21506_ (.RESET_B(net5231),
    .D(_01219_),
    .Q(\soc_inst.cpu_core.alu.b[21] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21507_ (.RESET_B(net5234),
    .D(_01220_),
    .Q(\soc_inst.cpu_core.alu.b[22] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _21508_ (.RESET_B(net5231),
    .D(_01221_),
    .Q(\soc_inst.cpu_core.alu.b[23] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _21509_ (.RESET_B(net5172),
    .D(_01222_),
    .Q(\soc_inst.cpu_core.alu.b[24] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _21510_ (.RESET_B(net5172),
    .D(_01223_),
    .Q(\soc_inst.cpu_core.alu.b[25] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _21511_ (.RESET_B(net5238),
    .D(_01224_),
    .Q(\soc_inst.cpu_core.alu.b[26] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _21512_ (.RESET_B(net5172),
    .D(_01225_),
    .Q(\soc_inst.cpu_core.alu.b[27] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _21513_ (.RESET_B(net5229),
    .D(_01226_),
    .Q(\soc_inst.cpu_core.alu.b[28] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _21514_ (.RESET_B(net5172),
    .D(net2912),
    .Q(\soc_inst.cpu_core.alu.b[29] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _21515_ (.RESET_B(net5235),
    .D(_01228_),
    .Q(\soc_inst.cpu_core.alu.b[30] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21516_ (.RESET_B(net5236),
    .D(net2284),
    .Q(\soc_inst.cpu_core.alu.b[31] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21517_ (.RESET_B(net5262),
    .D(net2106),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _21518_ (.RESET_B(net5268),
    .D(net2681),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _21519_ (.RESET_B(net5288),
    .D(net2558),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _21520_ (.RESET_B(net5290),
    .D(_01233_),
    .Q(\soc_inst.cpu_core.id_is_compressed ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21521_ (.RESET_B(net5367),
    .D(net2290),
    .Q(_00273_),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _21522_ (.RESET_B(net5366),
    .D(net2282),
    .Q(_00274_),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _21523_ (.RESET_B(net5358),
    .D(net2015),
    .Q(\soc_inst.cpu_core.ex_instr[2] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _21524_ (.RESET_B(net5357),
    .D(net2443),
    .Q(\soc_inst.cpu_core.ex_instr[3] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _21525_ (.RESET_B(net5367),
    .D(net2342),
    .Q(_00275_),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _21526_ (.RESET_B(net5358),
    .D(_01239_),
    .Q(\soc_inst.cpu_core.ex_instr[5] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _21527_ (.RESET_B(net5357),
    .D(net2710),
    .Q(\soc_inst.cpu_core.ex_instr[6] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _21528_ (.RESET_B(net5237),
    .D(net961),
    .Q(\soc_inst.cpu_core.ex_instr[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _21529_ (.RESET_B(net5288),
    .D(net2184),
    .Q(\soc_inst.cpu_core.ex_instr[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _21530_ (.RESET_B(net5288),
    .D(net1982),
    .Q(\soc_inst.cpu_core.ex_instr[9] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _21531_ (.RESET_B(net5288),
    .D(_01244_),
    .Q(\soc_inst.cpu_core.ex_instr[10] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _21532_ (.RESET_B(net5298),
    .D(_01245_),
    .Q(\soc_inst.cpu_core.ex_instr[11] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _21533_ (.RESET_B(net5325),
    .D(net2610),
    .Q(\soc_inst.cpu_core.ex_funct3[0] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _21534_ (.RESET_B(net5325),
    .D(_01247_),
    .Q(\soc_inst.cpu_core.ex_funct3[1] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _21535_ (.RESET_B(net5260),
    .D(_01248_),
    .Q(\soc_inst.cpu_core.ex_funct3[2] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _21536_ (.RESET_B(net5297),
    .D(net1049),
    .Q(\soc_inst.cpu_core.ex_instr[15] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _21537_ (.RESET_B(net5313),
    .D(net2152),
    .Q(\soc_inst.cpu_core.ex_instr[16] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _21538_ (.RESET_B(net5244),
    .D(net1004),
    .Q(\soc_inst.cpu_core.ex_instr[17] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _21539_ (.RESET_B(net5245),
    .D(_01252_),
    .Q(\soc_inst.cpu_core.ex_instr[18] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _21540_ (.RESET_B(net5251),
    .D(net1243),
    .Q(\soc_inst.cpu_core.ex_instr[19] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _21541_ (.RESET_B(net5312),
    .D(net2042),
    .Q(\soc_inst.cpu_core.ex_instr[20] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _21542_ (.RESET_B(net5250),
    .D(net2536),
    .Q(\soc_inst.cpu_core.ex_instr[21] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _21543_ (.RESET_B(net5312),
    .D(net2331),
    .Q(\soc_inst.cpu_core.ex_instr[22] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _21544_ (.RESET_B(net5312),
    .D(net1785),
    .Q(\soc_inst.cpu_core.ex_instr[23] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _21545_ (.RESET_B(net5258),
    .D(_01258_),
    .Q(\soc_inst.cpu_core.ex_instr[24] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _21546_ (.RESET_B(net5251),
    .D(net721),
    .Q(\soc_inst.cpu_core.ex_funct7[0] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _21547_ (.RESET_B(net5258),
    .D(_01260_),
    .Q(\soc_inst.cpu_core.ex_funct7[1] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _21548_ (.RESET_B(net5258),
    .D(net2079),
    .Q(\soc_inst.cpu_core.ex_funct7[2] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _21549_ (.RESET_B(net5250),
    .D(net2083),
    .Q(\soc_inst.cpu_core.ex_funct7[3] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _21550_ (.RESET_B(net5313),
    .D(_01263_),
    .Q(\soc_inst.cpu_core.ex_funct7[4] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _21551_ (.RESET_B(net5323),
    .D(_01264_),
    .Q(\soc_inst.cpu_core.ex_funct7[5] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _21552_ (.RESET_B(net5323),
    .D(net2270),
    .Q(\soc_inst.cpu_core.ex_funct7[6] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _21553_ (.RESET_B(net5325),
    .D(net1297),
    .Q(\soc_inst.cpu_core.ex_exception_pc[0] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _21554_ (.RESET_B(net5355),
    .D(net2186),
    .Q(\soc_inst.cpu_core.ex_exception_pc[1] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _21555_ (.RESET_B(net5356),
    .D(net1071),
    .Q(\soc_inst.cpu_core.ex_exception_pc[2] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _21556_ (.RESET_B(net5355),
    .D(net2246),
    .Q(\soc_inst.cpu_core.ex_exception_pc[3] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _21557_ (.RESET_B(net5356),
    .D(net1351),
    .Q(\soc_inst.cpu_core.ex_exception_pc[4] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _21558_ (.RESET_B(net5355),
    .D(net1749),
    .Q(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _21559_ (.RESET_B(net5355),
    .D(net1738),
    .Q(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _21560_ (.RESET_B(net5326),
    .D(net944),
    .Q(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21561_ (.RESET_B(net5326),
    .D(net1207),
    .Q(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21562_ (.RESET_B(net5326),
    .D(net860),
    .Q(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21563_ (.RESET_B(net5325),
    .D(net2052),
    .Q(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _21564_ (.RESET_B(net5325),
    .D(net919),
    .Q(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _21565_ (.RESET_B(net5322),
    .D(net1196),
    .Q(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _21566_ (.RESET_B(net5322),
    .D(net888),
    .Q(\soc_inst.cpu_core.ex_exception_pc[13] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _21567_ (.RESET_B(net5324),
    .D(net1167),
    .Q(\soc_inst.cpu_core.ex_exception_pc[14] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _21568_ (.RESET_B(net5312),
    .D(net1162),
    .Q(\soc_inst.cpu_core.ex_exception_pc[15] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _21569_ (.RESET_B(net5310),
    .D(net1958),
    .Q(\soc_inst.cpu_core.ex_exception_pc[16] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _21570_ (.RESET_B(net5310),
    .D(net1659),
    .Q(\soc_inst.cpu_core.ex_exception_pc[17] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _21571_ (.RESET_B(net5310),
    .D(net1247),
    .Q(\soc_inst.cpu_core.ex_exception_pc[18] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _21572_ (.RESET_B(net5313),
    .D(net1420),
    .Q(\soc_inst.cpu_core.ex_exception_pc[19] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _21573_ (.RESET_B(net5311),
    .D(net1510),
    .Q(\soc_inst.cpu_core.ex_exception_pc[20] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _21574_ (.RESET_B(net5313),
    .D(net1570),
    .Q(\soc_inst.cpu_core.ex_exception_pc[21] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _21575_ (.RESET_B(net5310),
    .D(net1647),
    .Q(\soc_inst.cpu_core.ex_exception_pc[22] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _21576_ (.RESET_B(net5311),
    .D(net1440),
    .Q(\soc_inst.cpu_core.ex_exception_pc[23] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _21577_ (.RESET_B(net5372),
    .D(net527),
    .Q(\soc_inst.core_mem_re ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _21578_ (.RESET_B(net5371),
    .D(net1214),
    .Q(\soc_inst.cpu_core.ex_rs1_data[0] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _21579_ (.RESET_B(net5255),
    .D(_01291_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _21580_ (.RESET_B(net5359),
    .D(net802),
    .Q(\soc_inst.cpu_core.ex_rs1_data[2] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _21581_ (.RESET_B(net5367),
    .D(net858),
    .Q(\soc_inst.cpu_core.ex_rs1_data[3] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _21582_ (.RESET_B(net5297),
    .D(net258),
    .Q(\soc_inst.cpu_core.ex_rs1_data[4] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _21583_ (.RESET_B(net5299),
    .D(net306),
    .Q(\soc_inst.cpu_core.ex_rs1_data[5] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _21584_ (.RESET_B(net5300),
    .D(net353),
    .Q(\soc_inst.cpu_core.ex_rs1_data[6] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _21585_ (.RESET_B(net5299),
    .D(net272),
    .Q(\soc_inst.cpu_core.ex_rs1_data[7] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _21586_ (.RESET_B(net5295),
    .D(net1145),
    .Q(\soc_inst.cpu_core.ex_rs1_data[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _21587_ (.RESET_B(net5260),
    .D(net2590),
    .Q(\soc_inst.cpu_core.ex_rs1_data[9] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _21588_ (.RESET_B(net5355),
    .D(_01300_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[10] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _21589_ (.RESET_B(net5260),
    .D(_01301_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[11] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _21590_ (.RESET_B(net5257),
    .D(net2108),
    .Q(\soc_inst.cpu_core.ex_rs1_data[12] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _21591_ (.RESET_B(net5257),
    .D(net781),
    .Q(\soc_inst.cpu_core.ex_rs1_data[13] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _21592_ (.RESET_B(net5254),
    .D(net836),
    .Q(\soc_inst.cpu_core.ex_rs1_data[14] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _21593_ (.RESET_B(net5258),
    .D(net445),
    .Q(\soc_inst.cpu_core.ex_rs1_data[15] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _21594_ (.RESET_B(net5310),
    .D(_01306_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[16] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _21595_ (.RESET_B(net5249),
    .D(_01307_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[17] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _21596_ (.RESET_B(net5247),
    .D(net874),
    .Q(\soc_inst.cpu_core.ex_rs1_data[18] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _21597_ (.RESET_B(net5247),
    .D(net738),
    .Q(\soc_inst.cpu_core.ex_rs1_data[19] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _21598_ (.RESET_B(net5309),
    .D(net1315),
    .Q(\soc_inst.cpu_core.ex_rs1_data[20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _21599_ (.RESET_B(net5247),
    .D(net731),
    .Q(\soc_inst.cpu_core.ex_rs1_data[21] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _21600_ (.RESET_B(net5247),
    .D(net648),
    .Q(\soc_inst.cpu_core.ex_rs1_data[22] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _21601_ (.RESET_B(net5309),
    .D(net756),
    .Q(\soc_inst.cpu_core.ex_rs1_data[23] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _21602_ (.RESET_B(net5348),
    .D(_01314_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[24] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _21603_ (.RESET_B(net5339),
    .D(net878),
    .Q(\soc_inst.cpu_core.ex_rs1_data[25] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _21604_ (.RESET_B(net5259),
    .D(net2265),
    .Q(\soc_inst.cpu_core.ex_rs1_data[26] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _21605_ (.RESET_B(net5343),
    .D(_01317_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[27] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _21606_ (.RESET_B(net5401),
    .D(_01318_),
    .Q(\soc_inst.cpu_core.ex_rs1_data[28] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _21607_ (.RESET_B(net5404),
    .D(net848),
    .Q(\soc_inst.cpu_core.ex_rs1_data[29] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _21608_ (.RESET_B(net5251),
    .D(net2093),
    .Q(\soc_inst.cpu_core.ex_rs1_data[30] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _21609_ (.RESET_B(net5259),
    .D(net2634),
    .Q(\soc_inst.cpu_core.ex_rs1_data[31] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _21610_ (.RESET_B(net5380),
    .D(net2761),
    .Q(\soc_inst.core_mem_addr[0] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _21611_ (.RESET_B(net5380),
    .D(_01323_),
    .Q(\soc_inst.core_mem_addr[1] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _21612_ (.RESET_B(net5382),
    .D(net2752),
    .Q(\soc_inst.core_mem_addr[2] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _21613_ (.RESET_B(net5382),
    .D(net2778),
    .Q(\soc_inst.core_mem_addr[3] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _21614_ (.RESET_B(net5384),
    .D(net2744),
    .Q(\soc_inst.pwm_inst.channel_idx [0]),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _21615_ (.RESET_B(net5385),
    .D(net2018),
    .Q(\soc_inst.core_mem_addr[5] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _21616_ (.RESET_B(net5385),
    .D(net1903),
    .Q(\soc_inst.core_mem_addr[6] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _21617_ (.RESET_B(net5385),
    .D(net1799),
    .Q(\soc_inst.core_mem_addr[7] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _21618_ (.RESET_B(net5379),
    .D(net2584),
    .Q(\soc_inst.core_mem_addr[8] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _21619_ (.RESET_B(net5364),
    .D(net2372),
    .Q(\soc_inst.core_mem_addr[9] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _21620_ (.RESET_B(net5362),
    .D(net2196),
    .Q(\soc_inst.core_mem_addr[10] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _21621_ (.RESET_B(net5373),
    .D(net1808),
    .Q(\soc_inst.core_mem_addr[11] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _21622_ (.RESET_B(net5383),
    .D(_01334_),
    .Q(\soc_inst.core_mem_addr[12] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _21623_ (.RESET_B(net5350),
    .D(_01335_),
    .Q(\soc_inst.core_mem_addr[13] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _21624_ (.RESET_B(net5384),
    .D(net2490),
    .Q(\soc_inst.core_mem_addr[14] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _21625_ (.RESET_B(net5384),
    .D(_01337_),
    .Q(\soc_inst.core_mem_addr[15] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _21626_ (.RESET_B(net5341),
    .D(_01338_),
    .Q(\soc_inst.core_mem_addr[16] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _21627_ (.RESET_B(net5340),
    .D(_01339_),
    .Q(\soc_inst.core_mem_addr[17] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _21628_ (.RESET_B(net5335),
    .D(_01340_),
    .Q(\soc_inst.core_mem_addr[18] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _21629_ (.RESET_B(net5337),
    .D(_01341_),
    .Q(\soc_inst.core_mem_addr[19] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _21630_ (.RESET_B(net5336),
    .D(_01342_),
    .Q(\soc_inst.core_mem_addr[20] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _21631_ (.RESET_B(net5320),
    .D(_01343_),
    .Q(\soc_inst.core_mem_addr[21] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _21632_ (.RESET_B(net5320),
    .D(_01344_),
    .Q(\soc_inst.core_mem_addr[22] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _21633_ (.RESET_B(net5320),
    .D(_01345_),
    .Q(\soc_inst.core_mem_addr[23] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _21634_ (.RESET_B(net5359),
    .D(net2268),
    .Q(\soc_inst.core_mem_addr[24] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _21635_ (.RESET_B(net5359),
    .D(net2347),
    .Q(\soc_inst.core_mem_addr[25] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _21636_ (.RESET_B(net5366),
    .D(net2154),
    .Q(\soc_inst.core_mem_addr[26] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _21637_ (.RESET_B(net5366),
    .D(net2413),
    .Q(\soc_inst.core_mem_addr[27] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _21638_ (.RESET_B(net5312),
    .D(net2260),
    .Q(\soc_inst.core_mem_addr[28] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _21639_ (.RESET_B(net5314),
    .D(net634),
    .Q(\soc_inst.core_mem_addr[29] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _21640_ (.RESET_B(net5362),
    .D(net1879),
    .Q(\soc_inst.core_mem_addr[30] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _21641_ (.RESET_B(net5322),
    .D(net2255),
    .Q(\soc_inst.core_mem_addr[31] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _21642_ (.RESET_B(net5368),
    .D(net337),
    .Q(\soc_inst.cpu_core.ex_rs2_data[0] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _21643_ (.RESET_B(net5283),
    .D(_01355_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[1] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _21644_ (.RESET_B(net5369),
    .D(_01356_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _21645_ (.RESET_B(net5302),
    .D(_01357_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[3] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _21646_ (.RESET_B(net5301),
    .D(net400),
    .Q(\soc_inst.cpu_core.ex_rs2_data[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _21647_ (.RESET_B(net5301),
    .D(net365),
    .Q(\soc_inst.cpu_core.ex_rs2_data[5] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _21648_ (.RESET_B(net5369),
    .D(_01360_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[6] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _21649_ (.RESET_B(net5299),
    .D(_01361_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[7] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _21650_ (.RESET_B(net5366),
    .D(net708),
    .Q(\soc_inst.cpu_core.ex_rs2_data[8] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _21651_ (.RESET_B(net5371),
    .D(net941),
    .Q(\soc_inst.cpu_core.ex_rs2_data[9] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _21652_ (.RESET_B(net5369),
    .D(net718),
    .Q(\soc_inst.cpu_core.ex_rs2_data[10] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _21653_ (.RESET_B(net5370),
    .D(net1477),
    .Q(\soc_inst.cpu_core.ex_rs2_data[11] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _21654_ (.RESET_B(net5369),
    .D(_01366_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[12] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _21655_ (.RESET_B(net5257),
    .D(_01367_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[13] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _21656_ (.RESET_B(net5325),
    .D(_01368_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[14] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _21657_ (.RESET_B(net5301),
    .D(net373),
    .Q(\soc_inst.cpu_core.ex_rs2_data[15] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _21658_ (.RESET_B(net5409),
    .D(_01370_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[16] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _21659_ (.RESET_B(net5247),
    .D(net2445),
    .Q(\soc_inst.cpu_core.ex_rs2_data[17] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _21660_ (.RESET_B(net5401),
    .D(net1086),
    .Q(\soc_inst.cpu_core.ex_rs2_data[18] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _21661_ (.RESET_B(net5441),
    .D(net312),
    .Q(\soc_inst.cpu_core.ex_rs2_data[19] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _21662_ (.RESET_B(net5309),
    .D(net1649),
    .Q(\soc_inst.cpu_core.ex_rs2_data[20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _21663_ (.RESET_B(net5402),
    .D(_01375_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[21] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _21664_ (.RESET_B(net5293),
    .D(net2236),
    .Q(\soc_inst.cpu_core.ex_rs2_data[22] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _21665_ (.RESET_B(net5310),
    .D(net1973),
    .Q(\soc_inst.cpu_core.ex_rs2_data[23] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _21666_ (.RESET_B(net5299),
    .D(net498),
    .Q(\soc_inst.cpu_core.ex_rs2_data[24] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _21667_ (.RESET_B(net5367),
    .D(_01379_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[25] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _21668_ (.RESET_B(net5296),
    .D(_01380_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[26] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _21669_ (.RESET_B(net5384),
    .D(net317),
    .Q(\soc_inst.cpu_core.ex_rs2_data[27] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _21670_ (.RESET_B(net5367),
    .D(net1875),
    .Q(\soc_inst.cpu_core.ex_rs2_data[28] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _21671_ (.RESET_B(net5296),
    .D(_01383_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[29] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _21672_ (.RESET_B(net5296),
    .D(_01384_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[30] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _21673_ (.RESET_B(net5440),
    .D(net864),
    .Q(\soc_inst.cpu_core.ex_rs2_data[31] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _21674_ (.RESET_B(net5235),
    .D(_01386_),
    .Q(\soc_inst.cpu_core.ex_alu_result[0] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _21675_ (.RESET_B(net5235),
    .D(_01387_),
    .Q(\soc_inst.cpu_core.ex_alu_result[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _21676_ (.RESET_B(net5237),
    .D(_01388_),
    .Q(\soc_inst.cpu_core.ex_alu_result[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21677_ (.RESET_B(net5238),
    .D(_01389_),
    .Q(\soc_inst.cpu_core.ex_alu_result[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21678_ (.RESET_B(net5256),
    .D(_01390_),
    .Q(\soc_inst.cpu_core.ex_alu_result[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _21679_ (.RESET_B(net5262),
    .D(net2924),
    .Q(\soc_inst.cpu_core.ex_alu_result[5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _21680_ (.RESET_B(net5211),
    .D(_01392_),
    .Q(\soc_inst.cpu_core.ex_alu_result[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _21681_ (.RESET_B(net5238),
    .D(_01393_),
    .Q(\soc_inst.cpu_core.ex_alu_result[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _21682_ (.RESET_B(net5240),
    .D(net2818),
    .Q(\soc_inst.cpu_core.ex_alu_result[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _21683_ (.RESET_B(net5240),
    .D(_01395_),
    .Q(\soc_inst.cpu_core.ex_alu_result[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21684_ (.RESET_B(net5255),
    .D(_01396_),
    .Q(\soc_inst.cpu_core.ex_alu_result[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _21685_ (.RESET_B(net5238),
    .D(_01397_),
    .Q(\soc_inst.cpu_core.ex_alu_result[11] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21686_ (.RESET_B(net5235),
    .D(net2834),
    .Q(\soc_inst.cpu_core.ex_alu_result[12] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21687_ (.RESET_B(net5232),
    .D(_01399_),
    .Q(\soc_inst.cpu_core.ex_alu_result[13] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21688_ (.RESET_B(net5232),
    .D(_01400_),
    .Q(\soc_inst.cpu_core.ex_alu_result[14] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21689_ (.RESET_B(net5232),
    .D(_01401_),
    .Q(\soc_inst.cpu_core.ex_alu_result[15] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21690_ (.RESET_B(net5250),
    .D(_01402_),
    .Q(\soc_inst.cpu_core.ex_alu_result[16] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _21691_ (.RESET_B(net5248),
    .D(_01403_),
    .Q(\soc_inst.cpu_core.ex_alu_result[17] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _21692_ (.RESET_B(net5248),
    .D(_01404_),
    .Q(\soc_inst.cpu_core.ex_alu_result[18] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _21693_ (.RESET_B(net5248),
    .D(_01405_),
    .Q(\soc_inst.cpu_core.ex_alu_result[19] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _21694_ (.RESET_B(net5248),
    .D(_01406_),
    .Q(\soc_inst.cpu_core.ex_alu_result[20] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _21695_ (.RESET_B(net5244),
    .D(_01407_),
    .Q(\soc_inst.cpu_core.ex_alu_result[21] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _21696_ (.RESET_B(net5243),
    .D(_01408_),
    .Q(\soc_inst.cpu_core.ex_alu_result[22] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21697_ (.RESET_B(net5242),
    .D(_01409_),
    .Q(\soc_inst.cpu_core.ex_alu_result[23] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _21698_ (.RESET_B(net5245),
    .D(_01410_),
    .Q(\soc_inst.cpu_core.ex_alu_result[24] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _21699_ (.RESET_B(net5265),
    .D(_01411_),
    .Q(\soc_inst.cpu_core.ex_alu_result[25] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _21700_ (.RESET_B(net5238),
    .D(_01412_),
    .Q(\soc_inst.cpu_core.ex_alu_result[26] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _21701_ (.RESET_B(net5259),
    .D(_01413_),
    .Q(\soc_inst.cpu_core.ex_alu_result[27] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _21702_ (.RESET_B(net5244),
    .D(_01414_),
    .Q(\soc_inst.cpu_core.ex_alu_result[28] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _21703_ (.RESET_B(net5251),
    .D(_01415_),
    .Q(\soc_inst.cpu_core.ex_alu_result[29] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _21704_ (.RESET_B(net5244),
    .D(_01416_),
    .Q(\soc_inst.cpu_core.ex_alu_result[30] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _21705_ (.RESET_B(net5235),
    .D(_01417_),
    .Q(\soc_inst.cpu_core.ex_alu_result[31] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _21706_ (.RESET_B(net5372),
    .D(_00025_),
    .Q(\soc_inst.core_mem_we ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _21707_ (.RESET_B(net5358),
    .D(net351),
    .Q(\soc_inst.cpu_core.ex_mem_we ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _21708_ (.RESET_B(net5363),
    .D(_01419_),
    .Q(\soc_inst.cpu_core.ex_mem_re ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _21709_ (.RESET_B(net5177),
    .D(_01420_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21710_ (.RESET_B(net5192),
    .D(_01421_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _21711_ (.RESET_B(net5183),
    .D(_01422_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _21712_ (.RESET_B(net5191),
    .D(_01423_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _21713_ (.RESET_B(net5217),
    .D(_01424_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _21714_ (.RESET_B(net5200),
    .D(_01425_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _21715_ (.RESET_B(net5216),
    .D(_01426_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _21716_ (.RESET_B(net5192),
    .D(_01427_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _21717_ (.RESET_B(net5149),
    .D(_01428_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _21718_ (.RESET_B(net5205),
    .D(_01429_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _21719_ (.RESET_B(net5176),
    .D(_01430_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _21720_ (.RESET_B(net5180),
    .D(_01431_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _21721_ (.RESET_B(net5208),
    .D(_01432_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][12] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _21722_ (.RESET_B(net5145),
    .D(_01433_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _21723_ (.RESET_B(net5209),
    .D(_01434_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][14] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _21724_ (.RESET_B(net5169),
    .D(_01435_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][15] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _21725_ (.RESET_B(net5144),
    .D(_01436_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _21726_ (.RESET_B(net5159),
    .D(_01437_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _21727_ (.RESET_B(net5130),
    .D(_01438_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][18] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _21728_ (.RESET_B(net5137),
    .D(_01439_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][19] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _21729_ (.RESET_B(net5136),
    .D(_01440_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][20] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _21730_ (.RESET_B(net5161),
    .D(_01441_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _21731_ (.RESET_B(net5142),
    .D(_01442_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _21732_ (.RESET_B(net5130),
    .D(_01443_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _21733_ (.RESET_B(net5154),
    .D(_01444_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _21734_ (.RESET_B(net5204),
    .D(_01445_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][25] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _21735_ (.RESET_B(net5184),
    .D(_01446_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][26] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21736_ (.RESET_B(net5166),
    .D(_01447_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][27] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _21737_ (.RESET_B(net5140),
    .D(_01448_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _21738_ (.RESET_B(net5163),
    .D(_01449_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21739_ (.RESET_B(net5186),
    .D(_01450_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21740_ (.RESET_B(net5153),
    .D(_01451_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][31] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21741_ (.RESET_B(net5177),
    .D(_01452_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _21742_ (.RESET_B(net5192),
    .D(_01453_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _21743_ (.RESET_B(net5183),
    .D(_01454_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _21744_ (.RESET_B(net5191),
    .D(_01455_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _21745_ (.RESET_B(net5217),
    .D(_01456_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _21746_ (.RESET_B(net5199),
    .D(_01457_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _21747_ (.RESET_B(net5216),
    .D(_01458_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][6] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _21748_ (.RESET_B(net5199),
    .D(_01459_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _21749_ (.RESET_B(net5148),
    .D(_01460_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _21750_ (.RESET_B(net5205),
    .D(_01461_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][9] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21751_ (.RESET_B(net5175),
    .D(_01462_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21752_ (.RESET_B(net5180),
    .D(_01463_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _21753_ (.RESET_B(net5208),
    .D(_01464_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][12] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _21754_ (.RESET_B(net5145),
    .D(_01465_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _21755_ (.RESET_B(net5209),
    .D(_01466_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _21756_ (.RESET_B(net5168),
    .D(_01467_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _21757_ (.RESET_B(net5144),
    .D(_01468_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _21758_ (.RESET_B(net5160),
    .D(_01469_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _21759_ (.RESET_B(net5130),
    .D(_01470_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _21760_ (.RESET_B(net5138),
    .D(_01471_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][19] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _21761_ (.RESET_B(net5136),
    .D(_01472_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][20] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _21762_ (.RESET_B(net5159),
    .D(_01473_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _21763_ (.RESET_B(net5142),
    .D(_01474_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][22] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21764_ (.RESET_B(net5132),
    .D(_01475_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _21765_ (.RESET_B(net5155),
    .D(_01476_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _21766_ (.RESET_B(net5207),
    .D(_01477_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][25] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _21767_ (.RESET_B(net5179),
    .D(_01478_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][26] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _21768_ (.RESET_B(net5166),
    .D(_01479_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][27] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _21769_ (.RESET_B(net5140),
    .D(_01480_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _21770_ (.RESET_B(net5162),
    .D(_01481_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21771_ (.RESET_B(net5186),
    .D(_01482_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _21772_ (.RESET_B(net5150),
    .D(_01483_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][31] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _21773_ (.RESET_B(net5177),
    .D(_01484_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _21774_ (.RESET_B(net5196),
    .D(_01485_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21775_ (.RESET_B(net5188),
    .D(_01486_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _21776_ (.RESET_B(net5194),
    .D(_01487_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _21777_ (.RESET_B(net5219),
    .D(_01488_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _21778_ (.RESET_B(net5201),
    .D(_01489_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _21779_ (.RESET_B(net5218),
    .D(_01490_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21780_ (.RESET_B(net5201),
    .D(_01491_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _21781_ (.RESET_B(net5148),
    .D(_01492_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _21782_ (.RESET_B(net5205),
    .D(_01493_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _21783_ (.RESET_B(net5175),
    .D(_01494_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _21784_ (.RESET_B(net5180),
    .D(_01495_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][11] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _21785_ (.RESET_B(net5208),
    .D(_01496_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][12] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _21786_ (.RESET_B(net5146),
    .D(_01497_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _21787_ (.RESET_B(net5209),
    .D(_01498_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][14] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _21788_ (.RESET_B(net5169),
    .D(_01499_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _21789_ (.RESET_B(net5144),
    .D(_01500_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _21790_ (.RESET_B(net5160),
    .D(_01501_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _21791_ (.RESET_B(net5129),
    .D(_01502_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _21792_ (.RESET_B(net5158),
    .D(_01503_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _21793_ (.RESET_B(net5131),
    .D(_01504_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _21794_ (.RESET_B(net5158),
    .D(_01505_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][21] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _21795_ (.RESET_B(net5164),
    .D(_01506_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][22] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21796_ (.RESET_B(net5132),
    .D(_01507_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _21797_ (.RESET_B(net5154),
    .D(_01508_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21798_ (.RESET_B(net5204),
    .D(_01509_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21799_ (.RESET_B(net5179),
    .D(_01510_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _21800_ (.RESET_B(net5156),
    .D(_01511_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21801_ (.RESET_B(net5141),
    .D(_01512_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][28] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _21802_ (.RESET_B(net5163),
    .D(_01513_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21803_ (.RESET_B(net5186),
    .D(_01514_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _21804_ (.RESET_B(net5152),
    .D(_01515_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][31] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _21805_ (.RESET_B(net5177),
    .D(_01516_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _21806_ (.RESET_B(net5201),
    .D(_01517_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _21807_ (.RESET_B(net5188),
    .D(_01518_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _21808_ (.RESET_B(net5194),
    .D(_01519_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _21809_ (.RESET_B(net5219),
    .D(_01520_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][4] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _21810_ (.RESET_B(net5202),
    .D(_01521_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][5] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _21811_ (.RESET_B(net5219),
    .D(_01522_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21812_ (.RESET_B(net5199),
    .D(_01523_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _21813_ (.RESET_B(net5148),
    .D(_01524_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _21814_ (.RESET_B(net5170),
    .D(_01525_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _21815_ (.RESET_B(net5177),
    .D(_01526_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][10] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _21816_ (.RESET_B(net5180),
    .D(_01527_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _21817_ (.RESET_B(net5210),
    .D(_01528_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][12] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _21818_ (.RESET_B(net5146),
    .D(_01529_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _21819_ (.RESET_B(net5213),
    .D(_01530_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _21820_ (.RESET_B(net5168),
    .D(_01531_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21821_ (.RESET_B(net5144),
    .D(_01532_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _21822_ (.RESET_B(net5174),
    .D(_01533_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _21823_ (.RESET_B(net5129),
    .D(_01534_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][18] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _21824_ (.RESET_B(net5137),
    .D(_01535_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][19] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _21825_ (.RESET_B(net5136),
    .D(_01536_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][20] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _21826_ (.RESET_B(net5158),
    .D(_01537_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][21] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21827_ (.RESET_B(net5164),
    .D(_01538_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][22] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21828_ (.RESET_B(net5132),
    .D(_01539_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _21829_ (.RESET_B(net5154),
    .D(_01540_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _21830_ (.RESET_B(net5204),
    .D(_01541_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][25] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21831_ (.RESET_B(net5179),
    .D(_01542_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _21832_ (.RESET_B(net5151),
    .D(_01543_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][27] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _21833_ (.RESET_B(net5141),
    .D(_01544_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][28] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _21834_ (.RESET_B(net5162),
    .D(_01545_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21835_ (.RESET_B(net5186),
    .D(_01546_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][30] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _21836_ (.RESET_B(net5152),
    .D(_01547_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _21837_ (.RESET_B(net5182),
    .D(_01548_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _21838_ (.RESET_B(net5193),
    .D(_01549_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21839_ (.RESET_B(net5190),
    .D(_01550_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21840_ (.RESET_B(net5194),
    .D(_01551_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _21841_ (.RESET_B(net5216),
    .D(_01552_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21842_ (.RESET_B(net5202),
    .D(_01553_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _21843_ (.RESET_B(net5218),
    .D(_01554_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21844_ (.RESET_B(net5196),
    .D(_01555_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][7] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21845_ (.RESET_B(net5148),
    .D(_01556_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _21846_ (.RESET_B(net5170),
    .D(_01557_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _21847_ (.RESET_B(net5175),
    .D(_01558_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21848_ (.RESET_B(net5193),
    .D(_01559_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _21849_ (.RESET_B(net5208),
    .D(_01560_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _21850_ (.RESET_B(net5145),
    .D(_01561_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _21851_ (.RESET_B(net5209),
    .D(_01562_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][14] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _21852_ (.RESET_B(net5168),
    .D(_01563_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21853_ (.RESET_B(net5144),
    .D(_01564_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _21854_ (.RESET_B(net5160),
    .D(_01565_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _21855_ (.RESET_B(net5129),
    .D(_01566_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _21856_ (.RESET_B(net5137),
    .D(_01567_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _21857_ (.RESET_B(net5139),
    .D(_01568_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _21858_ (.RESET_B(net5158),
    .D(_01569_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _21859_ (.RESET_B(net5164),
    .D(_01570_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21860_ (.RESET_B(net5132),
    .D(_01571_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _21861_ (.RESET_B(net5154),
    .D(_01572_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][24] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _21862_ (.RESET_B(net5204),
    .D(_01573_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][25] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21863_ (.RESET_B(net5179),
    .D(_01574_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][26] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _21864_ (.RESET_B(net5166),
    .D(_01575_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][27] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _21865_ (.RESET_B(net5140),
    .D(_01576_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _21866_ (.RESET_B(net5167),
    .D(_01577_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _21867_ (.RESET_B(net5186),
    .D(_01578_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][30] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _21868_ (.RESET_B(net5152),
    .D(_01579_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _21869_ (.RESET_B(net5178),
    .D(_01580_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21870_ (.RESET_B(net5192),
    .D(_01581_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21871_ (.RESET_B(net5188),
    .D(_01582_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _21872_ (.RESET_B(net5191),
    .D(_01583_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _21873_ (.RESET_B(net5216),
    .D(_01584_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _21874_ (.RESET_B(net5201),
    .D(_01585_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _21875_ (.RESET_B(net5200),
    .D(_01586_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _21876_ (.RESET_B(net5191),
    .D(_01587_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][7] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _21877_ (.RESET_B(net5150),
    .D(_01588_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _21878_ (.RESET_B(net5211),
    .D(_01589_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _21879_ (.RESET_B(net5176),
    .D(_01590_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21880_ (.RESET_B(net5181),
    .D(_01591_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _21881_ (.RESET_B(net5210),
    .D(_01592_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _21882_ (.RESET_B(net5145),
    .D(_01593_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _21883_ (.RESET_B(net5213),
    .D(_01594_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _21884_ (.RESET_B(net5168),
    .D(_01595_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _21885_ (.RESET_B(net5134),
    .D(_01596_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _21886_ (.RESET_B(net5162),
    .D(_01597_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][17] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21887_ (.RESET_B(net5130),
    .D(_01598_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][18] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _21888_ (.RESET_B(net5138),
    .D(_01599_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][19] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _21889_ (.RESET_B(net5131),
    .D(_01600_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][20] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _21890_ (.RESET_B(net5164),
    .D(_01601_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][21] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21891_ (.RESET_B(net5142),
    .D(_01602_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][22] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _21892_ (.RESET_B(net5133),
    .D(_01603_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _21893_ (.RESET_B(net5154),
    .D(_01604_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][24] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21894_ (.RESET_B(net5204),
    .D(_01605_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _21895_ (.RESET_B(net5179),
    .D(_01606_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][26] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _21896_ (.RESET_B(net5166),
    .D(_01607_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][27] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21897_ (.RESET_B(net5141),
    .D(_01608_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][28] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _21898_ (.RESET_B(net5163),
    .D(_01609_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21899_ (.RESET_B(net5186),
    .D(_01610_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][30] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _21900_ (.RESET_B(net5152),
    .D(_01611_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][31] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _21901_ (.RESET_B(net5177),
    .D(_01612_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _21902_ (.RESET_B(net5196),
    .D(_01613_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21903_ (.RESET_B(net5188),
    .D(_01614_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21904_ (.RESET_B(net5194),
    .D(_01615_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][3] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _21905_ (.RESET_B(net5219),
    .D(_01616_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21906_ (.RESET_B(net5202),
    .D(_01617_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _21907_ (.RESET_B(net5218),
    .D(_01618_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21908_ (.RESET_B(net5194),
    .D(_01619_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][7] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _21909_ (.RESET_B(net5149),
    .D(_01620_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21910_ (.RESET_B(net5170),
    .D(_01621_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _21911_ (.RESET_B(net5175),
    .D(_01622_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21912_ (.RESET_B(net5180),
    .D(_01623_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][11] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _21913_ (.RESET_B(net5208),
    .D(_01624_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _21914_ (.RESET_B(net5146),
    .D(_01625_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21915_ (.RESET_B(net5206),
    .D(_01626_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21916_ (.RESET_B(net5168),
    .D(_01627_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _21917_ (.RESET_B(net5147),
    .D(_01628_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21918_ (.RESET_B(net5162),
    .D(_01629_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][17] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _21919_ (.RESET_B(net5129),
    .D(_01630_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _21920_ (.RESET_B(net5137),
    .D(_01631_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][19] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _21921_ (.RESET_B(net5136),
    .D(_01632_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _21922_ (.RESET_B(net5159),
    .D(_01633_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _21923_ (.RESET_B(net5151),
    .D(_01634_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][22] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _21924_ (.RESET_B(net5133),
    .D(_01635_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _21925_ (.RESET_B(net5155),
    .D(_01636_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _21926_ (.RESET_B(net5185),
    .D(_01637_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _21927_ (.RESET_B(net5179),
    .D(_01638_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][26] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21928_ (.RESET_B(net5166),
    .D(_01639_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][27] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _21929_ (.RESET_B(net5141),
    .D(_01640_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _21930_ (.RESET_B(net5163),
    .D(_01641_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _21931_ (.RESET_B(net5187),
    .D(_01642_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][30] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _21932_ (.RESET_B(net5153),
    .D(_01643_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21933_ (.RESET_B(net5182),
    .D(_01644_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _21934_ (.RESET_B(net5196),
    .D(_01645_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21935_ (.RESET_B(net5183),
    .D(_01646_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _21936_ (.RESET_B(net5191),
    .D(_01647_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _21937_ (.RESET_B(net5217),
    .D(_01648_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _21938_ (.RESET_B(net5200),
    .D(_01649_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _21939_ (.RESET_B(net5219),
    .D(_01650_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _21940_ (.RESET_B(net5195),
    .D(_01651_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21941_ (.RESET_B(net5148),
    .D(_01652_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _21942_ (.RESET_B(net5211),
    .D(_01653_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _21943_ (.RESET_B(net5176),
    .D(_01654_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21944_ (.RESET_B(net5180),
    .D(_01655_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _21945_ (.RESET_B(net5210),
    .D(_01656_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _21946_ (.RESET_B(net5146),
    .D(_01657_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21947_ (.RESET_B(net5209),
    .D(_01658_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _21948_ (.RESET_B(net5169),
    .D(_01659_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _21949_ (.RESET_B(net5147),
    .D(_01660_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21950_ (.RESET_B(net5160),
    .D(_01661_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _21951_ (.RESET_B(net5130),
    .D(_01662_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _21952_ (.RESET_B(net5138),
    .D(_01663_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _21953_ (.RESET_B(net5136),
    .D(_01664_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _21954_ (.RESET_B(net5161),
    .D(_01665_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _21955_ (.RESET_B(net5143),
    .D(_01666_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _21956_ (.RESET_B(net5132),
    .D(_01667_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _21957_ (.RESET_B(net5155),
    .D(_01668_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _21958_ (.RESET_B(net5185),
    .D(_01669_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _21959_ (.RESET_B(net5179),
    .D(_01670_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _21960_ (.RESET_B(net5156),
    .D(_01671_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _21961_ (.RESET_B(net5141),
    .D(_01672_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _21962_ (.RESET_B(net5162),
    .D(_01673_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _21963_ (.RESET_B(net5187),
    .D(_01674_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][30] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _21964_ (.RESET_B(net5153),
    .D(_01675_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _21965_ (.RESET_B(net5177),
    .D(_01676_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _21966_ (.RESET_B(net5196),
    .D(_01677_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _21967_ (.RESET_B(net5183),
    .D(_01678_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21968_ (.RESET_B(net5194),
    .D(_01679_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _21969_ (.RESET_B(net5219),
    .D(_01680_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _21970_ (.RESET_B(net5202),
    .D(_01681_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _21971_ (.RESET_B(net5218),
    .D(_01682_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _21972_ (.RESET_B(net5193),
    .D(_01683_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _21973_ (.RESET_B(net5150),
    .D(_01684_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _21974_ (.RESET_B(net5205),
    .D(_01685_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _21975_ (.RESET_B(net5175),
    .D(_01686_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _21976_ (.RESET_B(net5181),
    .D(_01687_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][11] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _21977_ (.RESET_B(net5209),
    .D(_01688_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][12] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _21978_ (.RESET_B(net5146),
    .D(_01689_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _21979_ (.RESET_B(net5213),
    .D(_01690_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][14] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _21980_ (.RESET_B(net5169),
    .D(_01691_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _21981_ (.RESET_B(net5144),
    .D(_01692_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _21982_ (.RESET_B(net5160),
    .D(_01693_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _21983_ (.RESET_B(net5129),
    .D(_01694_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][18] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _21984_ (.RESET_B(net5137),
    .D(_01695_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][19] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _21985_ (.RESET_B(net5131),
    .D(_01696_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][20] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _21986_ (.RESET_B(net5159),
    .D(_01697_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _21987_ (.RESET_B(net5142),
    .D(_01698_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _21988_ (.RESET_B(net5132),
    .D(_01699_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _21989_ (.RESET_B(net5154),
    .D(_01700_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _21990_ (.RESET_B(net5204),
    .D(_01701_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][25] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _21991_ (.RESET_B(net5184),
    .D(_01702_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][26] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _21992_ (.RESET_B(net5151),
    .D(_01703_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _21993_ (.RESET_B(net5135),
    .D(_01704_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][28] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _21994_ (.RESET_B(net5167),
    .D(_01705_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][29] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _21995_ (.RESET_B(net5187),
    .D(_01706_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][30] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _21996_ (.RESET_B(net5152),
    .D(_01707_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][31] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _21997_ (.RESET_B(net5177),
    .D(_01708_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _21998_ (.RESET_B(net5192),
    .D(_01709_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _21999_ (.RESET_B(net5183),
    .D(_01710_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _22000_ (.RESET_B(net5191),
    .D(_01711_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _22001_ (.RESET_B(net5217),
    .D(_01712_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _22002_ (.RESET_B(net5200),
    .D(_01713_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _22003_ (.RESET_B(net5216),
    .D(_01714_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _22004_ (.RESET_B(net5192),
    .D(_01715_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][7] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _22005_ (.RESET_B(net5149),
    .D(_01716_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _22006_ (.RESET_B(net5205),
    .D(_01717_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _22007_ (.RESET_B(net5175),
    .D(_01718_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _22008_ (.RESET_B(net5180),
    .D(_01719_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _22009_ (.RESET_B(net5208),
    .D(_01720_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _22010_ (.RESET_B(net5146),
    .D(_01721_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _22011_ (.RESET_B(net5213),
    .D(_01722_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _22012_ (.RESET_B(net5169),
    .D(_01723_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][15] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _22013_ (.RESET_B(net5134),
    .D(_01724_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][16] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _22014_ (.RESET_B(net5174),
    .D(_01725_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _22015_ (.RESET_B(net5130),
    .D(_01726_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _22016_ (.RESET_B(net5137),
    .D(_01727_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _22017_ (.RESET_B(net5136),
    .D(_01728_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _22018_ (.RESET_B(net5158),
    .D(_01729_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][21] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _22019_ (.RESET_B(net5142),
    .D(_01730_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][22] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _22020_ (.RESET_B(net5133),
    .D(_01731_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _22021_ (.RESET_B(net5154),
    .D(_01732_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][24] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _22022_ (.RESET_B(net5185),
    .D(_01733_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][25] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _22023_ (.RESET_B(net5184),
    .D(_01734_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _22024_ (.RESET_B(net5166),
    .D(_01735_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][27] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _22025_ (.RESET_B(net5140),
    .D(_01736_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _22026_ (.RESET_B(net5162),
    .D(_01737_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][29] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _22027_ (.RESET_B(net5186),
    .D(_01738_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][30] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _22028_ (.RESET_B(net5150),
    .D(_01739_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][31] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _22029_ (.RESET_B(net5182),
    .D(_01740_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _22030_ (.RESET_B(net5196),
    .D(_01741_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _22031_ (.RESET_B(net5188),
    .D(_01742_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _22032_ (.RESET_B(net5194),
    .D(_01743_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][3] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _22033_ (.RESET_B(net5216),
    .D(_01744_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _22034_ (.RESET_B(net5201),
    .D(_01745_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _22035_ (.RESET_B(net5218),
    .D(_01746_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _22036_ (.RESET_B(net5195),
    .D(_01747_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][7] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _22037_ (.RESET_B(net5148),
    .D(_01748_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _22038_ (.RESET_B(net5170),
    .D(_01749_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _22039_ (.RESET_B(net5176),
    .D(_01750_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _22040_ (.RESET_B(net5181),
    .D(_01751_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _22041_ (.RESET_B(net5208),
    .D(_01752_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][12] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _22042_ (.RESET_B(net5145),
    .D(_01753_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _22043_ (.RESET_B(net5206),
    .D(_01754_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][14] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _22044_ (.RESET_B(net5168),
    .D(_01755_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _22045_ (.RESET_B(net5147),
    .D(_01756_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _22046_ (.RESET_B(net5159),
    .D(_01757_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][17] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _22047_ (.RESET_B(net5129),
    .D(_01758_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][18] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _22048_ (.RESET_B(net5137),
    .D(_01759_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _22049_ (.RESET_B(net5131),
    .D(_01760_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _22050_ (.RESET_B(net5158),
    .D(_01761_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _22051_ (.RESET_B(net5151),
    .D(_01762_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][22] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _22052_ (.RESET_B(net5133),
    .D(_01763_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][23] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _22053_ (.RESET_B(net5155),
    .D(_01764_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][24] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _22054_ (.RESET_B(net5207),
    .D(_01765_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][25] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _22055_ (.RESET_B(net5184),
    .D(_01766_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _22056_ (.RESET_B(net5166),
    .D(_01767_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][27] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _22057_ (.RESET_B(net5140),
    .D(_01768_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _22058_ (.RESET_B(net5167),
    .D(_01769_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _22059_ (.RESET_B(net5187),
    .D(_01770_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _22060_ (.RESET_B(net5153),
    .D(_01771_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][31] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _22061_ (.RESET_B(net5182),
    .D(_01772_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _22062_ (.RESET_B(net5193),
    .D(_01773_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _22063_ (.RESET_B(net5188),
    .D(_01774_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _22064_ (.RESET_B(net5191),
    .D(_01775_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _22065_ (.RESET_B(net5217),
    .D(_01776_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _22066_ (.RESET_B(net5201),
    .D(_01777_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _22067_ (.RESET_B(net5200),
    .D(_01778_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _22068_ (.RESET_B(net5199),
    .D(_01779_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][7] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _22069_ (.RESET_B(net5149),
    .D(_01780_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _22070_ (.RESET_B(net5205),
    .D(_01781_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _22071_ (.RESET_B(net5175),
    .D(_01782_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _22072_ (.RESET_B(net5181),
    .D(_01783_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][11] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _22073_ (.RESET_B(net5209),
    .D(_01784_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _22074_ (.RESET_B(net5145),
    .D(_01785_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _22075_ (.RESET_B(net5211),
    .D(_01786_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _22076_ (.RESET_B(net5168),
    .D(_01787_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _22077_ (.RESET_B(net5144),
    .D(_01788_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _22078_ (.RESET_B(net5159),
    .D(_01789_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _22079_ (.RESET_B(net5129),
    .D(_01790_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _22080_ (.RESET_B(net5158),
    .D(_01791_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][19] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _22081_ (.RESET_B(net5136),
    .D(_01792_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _22082_ (.RESET_B(net5158),
    .D(_01793_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _22083_ (.RESET_B(net5142),
    .D(_01794_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][22] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _22084_ (.RESET_B(net5132),
    .D(_01795_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _22085_ (.RESET_B(net5171),
    .D(_01796_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][24] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _22086_ (.RESET_B(net5204),
    .D(_01797_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][25] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _22087_ (.RESET_B(net5185),
    .D(_01798_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _22088_ (.RESET_B(net5151),
    .D(_01799_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][27] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _22089_ (.RESET_B(net5135),
    .D(_01800_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][28] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _22090_ (.RESET_B(net5167),
    .D(_01801_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _22091_ (.RESET_B(net5187),
    .D(_01802_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][30] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _22092_ (.RESET_B(net5152),
    .D(_01803_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][31] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _22093_ (.RESET_B(net5182),
    .D(_01804_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _22094_ (.RESET_B(net5196),
    .D(_01805_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _22095_ (.RESET_B(net5188),
    .D(_01806_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _22096_ (.RESET_B(net5194),
    .D(_01807_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _22097_ (.RESET_B(net5216),
    .D(_01808_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _22098_ (.RESET_B(net5199),
    .D(_01809_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _22099_ (.RESET_B(net5216),
    .D(_01810_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _22100_ (.RESET_B(net5195),
    .D(_01811_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][7] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _22101_ (.RESET_B(net5148),
    .D(_01812_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _22102_ (.RESET_B(net5205),
    .D(_01813_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _22103_ (.RESET_B(net5178),
    .D(_01814_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][10] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _22104_ (.RESET_B(net5181),
    .D(_01815_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _22105_ (.RESET_B(net5209),
    .D(_01816_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _22106_ (.RESET_B(net5145),
    .D(_01817_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _22107_ (.RESET_B(net5213),
    .D(_01818_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _22108_ (.RESET_B(net5169),
    .D(_01819_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][15] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _22109_ (.RESET_B(net5134),
    .D(_01820_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _22110_ (.RESET_B(net5160),
    .D(_01821_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][17] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _22111_ (.RESET_B(net5130),
    .D(_01822_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _22112_ (.RESET_B(net5138),
    .D(_01823_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][19] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _22113_ (.RESET_B(net5139),
    .D(_01824_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _22114_ (.RESET_B(net5161),
    .D(_01825_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][21] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _22115_ (.RESET_B(net5142),
    .D(_01826_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _22116_ (.RESET_B(net5133),
    .D(_01827_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _22117_ (.RESET_B(net5155),
    .D(_01828_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][24] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _22118_ (.RESET_B(net5204),
    .D(_01829_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][25] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _22119_ (.RESET_B(net5184),
    .D(_01830_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][26] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _22120_ (.RESET_B(net5166),
    .D(_01831_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][27] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _22121_ (.RESET_B(net5140),
    .D(_01832_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][28] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _22122_ (.RESET_B(net5167),
    .D(_01833_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _22123_ (.RESET_B(net5187),
    .D(_01834_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][30] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _22124_ (.RESET_B(net5152),
    .D(_01835_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _22125_ (.RESET_B(net5183),
    .D(_01836_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _22126_ (.RESET_B(net5192),
    .D(_01837_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _22127_ (.RESET_B(net5188),
    .D(_01838_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _22128_ (.RESET_B(net5199),
    .D(_01839_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _22129_ (.RESET_B(net5217),
    .D(_01840_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][4] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _22130_ (.RESET_B(net5213),
    .D(_01841_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _22131_ (.RESET_B(net5213),
    .D(_01842_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _22132_ (.RESET_B(net5199),
    .D(_01843_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _22133_ (.RESET_B(net5150),
    .D(_01844_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][8] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _22134_ (.RESET_B(net5211),
    .D(_01845_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _22135_ (.RESET_B(net5184),
    .D(_01846_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][10] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _22136_ (.RESET_B(net5199),
    .D(_01847_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][11] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _22137_ (.RESET_B(net5214),
    .D(_01848_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][12] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _22138_ (.RESET_B(net5151),
    .D(_01849_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _22139_ (.RESET_B(net5213),
    .D(_01850_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _22140_ (.RESET_B(net5173),
    .D(_01851_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][15] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _22141_ (.RESET_B(net5151),
    .D(_01852_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _22142_ (.RESET_B(net5165),
    .D(_01853_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][17] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _22143_ (.RESET_B(net5136),
    .D(_01854_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][18] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _22144_ (.RESET_B(net5162),
    .D(_01855_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _22145_ (.RESET_B(net5131),
    .D(_01856_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][20] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _22146_ (.RESET_B(net5160),
    .D(_01857_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][21] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _22147_ (.RESET_B(net5162),
    .D(_01858_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][22] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _22148_ (.RESET_B(net5140),
    .D(_01859_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][23] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _22149_ (.RESET_B(net5171),
    .D(_01860_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][24] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _22150_ (.RESET_B(net5205),
    .D(_01861_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][25] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _22151_ (.RESET_B(net5184),
    .D(_01862_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _22152_ (.RESET_B(net5155),
    .D(_01863_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][27] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _22153_ (.RESET_B(net5140),
    .D(_01864_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _22154_ (.RESET_B(net5167),
    .D(_01865_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _22155_ (.RESET_B(net5185),
    .D(_01866_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][30] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _22156_ (.RESET_B(net5170),
    .D(_01867_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][31] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _22157_ (.RESET_B(net5344),
    .D(_01868_),
    .Q(\soc_inst.cpu_core.csr_file.mie[7] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _22158_ (.RESET_B(net5344),
    .D(net644),
    .Q(\soc_inst.cpu_core.csr_file.mie[11] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _22159_ (.RESET_B(net5258),
    .D(_01870_),
    .Q(\soc_inst.cpu_core.ex_branch_target[0] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _22160_ (.RESET_B(net5295),
    .D(_01871_),
    .Q(\soc_inst.cpu_core.ex_branch_target[1] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _22161_ (.RESET_B(net5295),
    .D(_01872_),
    .Q(\soc_inst.cpu_core.ex_branch_target[2] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _22162_ (.RESET_B(net5295),
    .D(_01873_),
    .Q(\soc_inst.cpu_core.ex_branch_target[3] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _22163_ (.RESET_B(net5356),
    .D(_01874_),
    .Q(\soc_inst.cpu_core.ex_branch_target[4] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _22164_ (.RESET_B(net5358),
    .D(_01875_),
    .Q(\soc_inst.cpu_core.ex_branch_target[5] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _22165_ (.RESET_B(net5295),
    .D(_01876_),
    .Q(\soc_inst.cpu_core.ex_branch_target[6] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _22166_ (.RESET_B(net5356),
    .D(_01877_),
    .Q(\soc_inst.cpu_core.ex_branch_target[7] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _22167_ (.RESET_B(net5295),
    .D(net1462),
    .Q(\soc_inst.cpu_core.ex_branch_target[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _22168_ (.RESET_B(net5330),
    .D(net2209),
    .Q(\soc_inst.cpu_core.ex_branch_target[9] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _22169_ (.RESET_B(net5326),
    .D(_01880_),
    .Q(\soc_inst.cpu_core.ex_branch_target[10] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _22170_ (.RESET_B(net5260),
    .D(net1826),
    .Q(\soc_inst.cpu_core.ex_branch_target[11] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _22171_ (.RESET_B(net5258),
    .D(net1323),
    .Q(\soc_inst.cpu_core.ex_branch_target[12] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _22172_ (.RESET_B(net5326),
    .D(_01883_),
    .Q(\soc_inst.cpu_core.ex_branch_target[13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _22173_ (.RESET_B(net5257),
    .D(_01884_),
    .Q(\soc_inst.cpu_core.ex_branch_target[14] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _22174_ (.RESET_B(net5328),
    .D(_01885_),
    .Q(\soc_inst.cpu_core.ex_branch_target[15] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _22175_ (.RESET_B(net5250),
    .D(_01886_),
    .Q(\soc_inst.cpu_core.ex_branch_target[16] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _22176_ (.RESET_B(net5250),
    .D(net1302),
    .Q(\soc_inst.cpu_core.ex_branch_target[17] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _22177_ (.RESET_B(net5250),
    .D(_01888_),
    .Q(\soc_inst.cpu_core.ex_branch_target[18] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _22178_ (.RESET_B(net5251),
    .D(net2986),
    .Q(\soc_inst.cpu_core.ex_branch_target[19] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _22179_ (.RESET_B(net5249),
    .D(net2226),
    .Q(\soc_inst.cpu_core.ex_branch_target[20] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _22180_ (.RESET_B(net5247),
    .D(net2351),
    .Q(\soc_inst.cpu_core.ex_branch_target[21] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _22181_ (.RESET_B(net5313),
    .D(_01892_),
    .Q(\soc_inst.cpu_core.ex_branch_target[22] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _22182_ (.RESET_B(net5312),
    .D(_01893_),
    .Q(\soc_inst.cpu_core.ex_branch_target[23] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _22183_ (.RESET_B(net5245),
    .D(net1158),
    .Q(\soc_inst.cpu_core.ex_branch_target[24] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _22184_ (.RESET_B(net5245),
    .D(net1392),
    .Q(\soc_inst.cpu_core.ex_branch_target[25] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _22185_ (.RESET_B(net5258),
    .D(net937),
    .Q(\soc_inst.cpu_core.ex_branch_target[26] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _22186_ (.RESET_B(net5253),
    .D(net1877),
    .Q(\soc_inst.cpu_core.ex_branch_target[27] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _22187_ (.RESET_B(net5313),
    .D(_01898_),
    .Q(\soc_inst.cpu_core.ex_branch_target[28] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _22188_ (.RESET_B(net5251),
    .D(net1822),
    .Q(\soc_inst.cpu_core.ex_branch_target[29] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _22189_ (.RESET_B(net5254),
    .D(net1460),
    .Q(\soc_inst.cpu_core.ex_branch_target[30] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _22190_ (.RESET_B(net5257),
    .D(net1531),
    .Q(\soc_inst.cpu_core.ex_branch_target[31] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _22191_ (.RESET_B(net5225),
    .D(_01902_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _22192_ (.RESET_B(net5225),
    .D(net2927),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _22193_ (.RESET_B(net5378),
    .D(net602),
    .Q(\soc_inst.cpu_core.csr_file.mtval[5] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _22194_ (.RESET_B(net5382),
    .D(net615),
    .Q(\soc_inst.cpu_core.csr_file.mtval[6] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _22195_ (.RESET_B(net5346),
    .D(net579),
    .Q(\soc_inst.cpu_core.csr_file.mtval[7] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _22196_ (.RESET_B(net5352),
    .D(net1432),
    .Q(\soc_inst.cpu_core.csr_file.mtval[8] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _22197_ (.RESET_B(net5345),
    .D(net477),
    .Q(\soc_inst.cpu_core.csr_file.mtval[9] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _22198_ (.RESET_B(net5352),
    .D(net1568),
    .Q(\soc_inst.cpu_core.csr_file.mtval[10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _22199_ (.RESET_B(net5344),
    .D(net417),
    .Q(\soc_inst.cpu_core.csr_file.mtval[11] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _22200_ (.RESET_B(net5347),
    .D(net1521),
    .Q(\soc_inst.cpu_core.csr_file.mtval[12] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _22201_ (.RESET_B(net5328),
    .D(net459),
    .Q(\soc_inst.cpu_core.csr_file.mtval[13] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _22202_ (.RESET_B(net5350),
    .D(net1446),
    .Q(\soc_inst.cpu_core.csr_file.mtval[14] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _22203_ (.RESET_B(net5336),
    .D(net2039),
    .Q(\soc_inst.cpu_core.csr_file.mtval[15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _22204_ (.RESET_B(net5340),
    .D(net1272),
    .Q(\soc_inst.cpu_core.csr_file.mtval[16] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _22205_ (.RESET_B(net5340),
    .D(net510),
    .Q(\soc_inst.cpu_core.csr_file.mtval[17] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _22206_ (.RESET_B(net5319),
    .D(net2023),
    .Q(\soc_inst.cpu_core.csr_file.mtval[18] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _22207_ (.RESET_B(net5318),
    .D(net577),
    .Q(\soc_inst.cpu_core.csr_file.mtval[19] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _22208_ (.RESET_B(net5336),
    .D(net456),
    .Q(\soc_inst.cpu_core.csr_file.mtval[20] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _22209_ (.RESET_B(net5315),
    .D(net1852),
    .Q(\soc_inst.cpu_core.csr_file.mtval[21] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _22210_ (.RESET_B(net5319),
    .D(_01921_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[22] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _22211_ (.RESET_B(net5315),
    .D(net1941),
    .Q(\soc_inst.cpu_core.csr_file.mtval[23] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _22212_ (.RESET_B(net5343),
    .D(net1504),
    .Q(\soc_inst.cpu_core.csr_file.mtval[24] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _22213_ (.RESET_B(net5340),
    .D(_01924_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[25] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _22214_ (.RESET_B(net5349),
    .D(net2596),
    .Q(\soc_inst.cpu_core.csr_file.mtval[26] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _22215_ (.RESET_B(net5341),
    .D(net2400),
    .Q(\soc_inst.cpu_core.csr_file.mtval[27] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _22216_ (.RESET_B(net5341),
    .D(_01927_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[28] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _22217_ (.RESET_B(net5340),
    .D(_01928_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[29] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _22218_ (.RESET_B(net5342),
    .D(net2547),
    .Q(\soc_inst.cpu_core.csr_file.mtval[30] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _22219_ (.RESET_B(net5343),
    .D(_01930_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[31] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _22220_ (.RESET_B(net5378),
    .D(_01931_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[5] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _22221_ (.RESET_B(net5378),
    .D(net838),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[6] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _22222_ (.RESET_B(net5345),
    .D(_01933_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[7] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _22223_ (.RESET_B(net5352),
    .D(_01934_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[8] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _22224_ (.RESET_B(net5345),
    .D(net666),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[9] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _22225_ (.RESET_B(net5378),
    .D(net950),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _22226_ (.RESET_B(net5344),
    .D(_01937_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[11] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _22227_ (.RESET_B(net5347),
    .D(net1073),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[12] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _22228_ (.RESET_B(net5329),
    .D(net946),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[13] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _22229_ (.RESET_B(net5352),
    .D(net540),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[14] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _22230_ (.RESET_B(net5347),
    .D(net931),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[15] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _22231_ (.RESET_B(net5338),
    .D(net619),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[16] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _22232_ (.RESET_B(net5338),
    .D(net734),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[17] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _22233_ (.RESET_B(net5334),
    .D(net1198),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[18] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _22234_ (.RESET_B(net5334),
    .D(net632),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[19] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _22235_ (.RESET_B(net5335),
    .D(net1579),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[20] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _22236_ (.RESET_B(net5315),
    .D(net1887),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[21] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _22237_ (.RESET_B(net5334),
    .D(net1409),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[22] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _22238_ (.RESET_B(net5317),
    .D(net1200),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[23] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _22239_ (.RESET_B(net5379),
    .D(net1091),
    .Q(\soc_inst.cpu_core.csr_file.mepc[5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _22240_ (.RESET_B(net5379),
    .D(_01951_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[6] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _22241_ (.RESET_B(net5346),
    .D(net2684),
    .Q(\soc_inst.cpu_core.csr_file.mepc[7] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _22242_ (.RESET_B(net5345),
    .D(net1017),
    .Q(\soc_inst.cpu_core.csr_file.mepc[8] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _22243_ (.RESET_B(net5346),
    .D(net1000),
    .Q(\soc_inst.cpu_core.csr_file.mepc[9] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _22244_ (.RESET_B(net5379),
    .D(net1209),
    .Q(\soc_inst.cpu_core.csr_file.mepc[10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _22245_ (.RESET_B(net5347),
    .D(net2485),
    .Q(\soc_inst.cpu_core.csr_file.mepc[11] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _22246_ (.RESET_B(net5347),
    .D(_01957_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[12] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _22247_ (.RESET_B(net5328),
    .D(net790),
    .Q(\soc_inst.cpu_core.csr_file.mepc[13] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _22248_ (.RESET_B(net5350),
    .D(_01959_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[14] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _22249_ (.RESET_B(net5329),
    .D(net833),
    .Q(\soc_inst.cpu_core.csr_file.mepc[15] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _22250_ (.RESET_B(net5335),
    .D(_01961_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[16] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _22251_ (.RESET_B(net5335),
    .D(_01962_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[17] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _22252_ (.RESET_B(net5316),
    .D(net1105),
    .Q(\soc_inst.cpu_core.csr_file.mepc[18] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _22253_ (.RESET_B(net5316),
    .D(net1308),
    .Q(\soc_inst.cpu_core.csr_file.mepc[19] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _22254_ (.RESET_B(net5335),
    .D(_01965_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[20] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _22255_ (.RESET_B(net5316),
    .D(net1714),
    .Q(\soc_inst.cpu_core.csr_file.mepc[21] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _22256_ (.RESET_B(net5318),
    .D(net926),
    .Q(\soc_inst.cpu_core.csr_file.mepc[22] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _22257_ (.RESET_B(net5316),
    .D(_01968_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[23] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _22258_ (.RESET_B(net5341),
    .D(net2249),
    .Q(\soc_inst.cpu_core.csr_file.mcause[31] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _22259_ (.RESET_B(net5414),
    .D(net85),
    .Q(\soc_inst.cpu_core.csr_file.mip_tip ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _22260_ (.RESET_B(net5447),
    .D(_01970_),
    .Q(\soc_inst.pwm_ena[1] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22261_ (.RESET_B(net5447),
    .D(_01971_),
    .Q(\soc_inst.pwm_ena[0] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22262_ (.RESET_B(net5331),
    .D(_00063_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _22263_ (.RESET_B(net5474),
    .D(net281),
    .Q(\soc_inst.i2c_inst.ack_received ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _22264_ (.RESET_B(net5466),
    .D(\soc_inst.i2c_ena ),
    .Q(\soc_inst.i2c_inst.status_reg[0] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _22265_ (.RESET_B(net5466),
    .D(net90),
    .Q(\soc_inst.i2c_inst.status_reg[1] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _22266_ (.RESET_B(net5467),
    .D(net89),
    .Q(\soc_inst.i2c_inst.status_reg[2] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _22267_ (.RESET_B(net5467),
    .D(net81),
    .Q(\soc_inst.i2c_inst.status_reg[3] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _22268_ (.RESET_B(net5456),
    .D(_01973_),
    .Q(\soc_inst.gpio_inst.int_pend_reg[6] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _22269_ (.RESET_B(net5459),
    .D(net564),
    .Q(\soc_inst.gpio_inst.int_pend_reg[5] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _22270_ (.RESET_B(net5458),
    .D(net359),
    .Q(\soc_inst.gpio_inst.int_pend_reg[4] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _22271_ (.RESET_B(net5460),
    .D(net382),
    .Q(\soc_inst.gpio_inst.int_pend_reg[3] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _22272_ (.RESET_B(net5458),
    .D(net485),
    .Q(\soc_inst.gpio_inst.int_pend_reg[2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _22273_ (.RESET_B(net5460),
    .D(_01978_),
    .Q(\soc_inst.gpio_inst.int_pend_reg[1] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _22274_ (.RESET_B(net5355),
    .D(_01979_),
    .Q(\soc_inst.cpu_core.id_pc[0] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _22275_ (.RESET_B(net5358),
    .D(_01980_),
    .Q(\soc_inst.cpu_core.id_pc[1] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _22276_ (.RESET_B(net5355),
    .D(_01981_),
    .Q(\soc_inst.cpu_core.id_pc[2] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _22277_ (.RESET_B(net5357),
    .D(_01982_),
    .Q(\soc_inst.cpu_core.id_pc[3] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _22278_ (.RESET_B(net5296),
    .D(_01983_),
    .Q(\soc_inst.cpu_core.id_pc[4] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _22279_ (.RESET_B(net5357),
    .D(_01984_),
    .Q(\soc_inst.cpu_core.id_pc[5] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _22280_ (.RESET_B(net5296),
    .D(_01985_),
    .Q(\soc_inst.cpu_core.id_pc[6] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _22281_ (.RESET_B(net5357),
    .D(_01986_),
    .Q(\soc_inst.cpu_core.id_pc[7] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _22282_ (.RESET_B(net5327),
    .D(_01987_),
    .Q(\soc_inst.cpu_core.id_pc[8] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _22283_ (.RESET_B(net5327),
    .D(_01988_),
    .Q(\soc_inst.cpu_core.id_pc[9] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _22284_ (.RESET_B(net5260),
    .D(_01989_),
    .Q(\soc_inst.cpu_core.id_pc[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _22285_ (.RESET_B(net5260),
    .D(_01990_),
    .Q(\soc_inst.cpu_core.id_pc[11] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _22286_ (.RESET_B(net5260),
    .D(_01991_),
    .Q(\soc_inst.cpu_core.id_pc[12] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _22287_ (.RESET_B(net5323),
    .D(_01992_),
    .Q(\soc_inst.cpu_core.id_pc[13] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _22288_ (.RESET_B(net5257),
    .D(_01993_),
    .Q(\soc_inst.cpu_core.id_pc[14] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _22289_ (.RESET_B(net5257),
    .D(_01994_),
    .Q(\soc_inst.cpu_core.id_pc[15] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _22290_ (.RESET_B(net5313),
    .D(_01995_),
    .Q(\soc_inst.cpu_core.id_pc[16] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _22291_ (.RESET_B(net5249),
    .D(_01996_),
    .Q(\soc_inst.cpu_core.id_pc[17] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _22292_ (.RESET_B(net5249),
    .D(_01997_),
    .Q(\soc_inst.cpu_core.id_pc[18] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _22293_ (.RESET_B(net5249),
    .D(_01998_),
    .Q(\soc_inst.cpu_core.id_pc[19] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _22294_ (.RESET_B(net5249),
    .D(_01999_),
    .Q(\soc_inst.cpu_core.id_pc[20] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _22295_ (.RESET_B(net5249),
    .D(_02000_),
    .Q(\soc_inst.cpu_core.id_pc[21] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _22296_ (.RESET_B(net5243),
    .D(_02001_),
    .Q(\soc_inst.cpu_core.id_pc[22] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _22297_ (.RESET_B(net5243),
    .D(_02002_),
    .Q(\soc_inst.cpu_core.id_pc[23] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _22298_ (.RESET_B(net5375),
    .D(_00332_),
    .Q(_00276_),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _22299_ (.RESET_B(net5375),
    .D(_00006_),
    .Q(\soc_inst.mem_ctrl.access_state[1] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _22300_ (.RESET_B(net5375),
    .D(_00007_),
    .Q(\soc_inst.mem_ctrl.access_state[2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _22301_ (.RESET_B(net5375),
    .D(net2567),
    .Q(\soc_inst.mem_ctrl.access_state[3] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _22302_ (.RESET_B(net5375),
    .D(_00009_),
    .Q(\soc_inst.mem_ctrl.access_state[4] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _22303_ (.RESET_B(net5422),
    .D(_02003_),
    .Q(_00277_),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _22304_ (.RESET_B(net5418),
    .D(_02004_),
    .Q(_00278_),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _22305_ (.RESET_B(net5419),
    .D(net1622),
    .Q(_00279_),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _22306_ (.RESET_B(net5419),
    .D(net1305),
    .Q(_00280_),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _22307_ (.RESET_B(net5445),
    .D(_02007_),
    .Q(_00281_),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _22308_ (.RESET_B(net5422),
    .D(_02008_),
    .Q(_00282_),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _22309_ (.RESET_B(net5445),
    .D(_02009_),
    .Q(_00283_),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _22310_ (.RESET_B(net5422),
    .D(_02010_),
    .Q(_00284_),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _22311_ (.RESET_B(net5418),
    .D(net1518),
    .Q(_00285_),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _22312_ (.RESET_B(net5418),
    .D(_02012_),
    .Q(_00286_),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _22313_ (.RESET_B(net5419),
    .D(net1422),
    .Q(_00287_),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22314_ (.RESET_B(net5410),
    .D(net1417),
    .Q(_00288_),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _22315_ (.RESET_B(net5410),
    .D(net1384),
    .Q(_00289_),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _22316_ (.RESET_B(net5412),
    .D(net1787),
    .Q(_00290_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22317_ (.RESET_B(net5410),
    .D(net2117),
    .Q(_00291_),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _22318_ (.RESET_B(net5412),
    .D(_02018_),
    .Q(_00292_),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22319_ (.RESET_B(net5346),
    .D(net2085),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[7] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _22320_ (.RESET_B(net5344),
    .D(net2383),
    .Q(_00293_),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _22321_ (.RESET_B(net5347),
    .D(net2075),
    .Q(_00294_),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _22322_ (.RESET_B(net48),
    .D(net2406),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[0] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _22323_ (.RESET_B(net46),
    .D(net2241),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _22324_ (.RESET_B(net44),
    .D(net1980),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[2] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _22325_ (.RESET_B(net42),
    .D(net1963),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[3] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _22326_ (.RESET_B(net40),
    .D(net376),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _22327_ (.RESET_B(net38),
    .D(_02027_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[5] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _22328_ (.RESET_B(net70),
    .D(_02028_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _22329_ (.RESET_B(net71),
    .D(_00019_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[0] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22330_ (.RESET_B(net72),
    .D(net939),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22331_ (.RESET_B(net73),
    .D(_00021_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[2] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _22332_ (.RESET_B(net36),
    .D(_00022_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[3] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22333_ (.RESET_B(net5448),
    .D(_02029_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _22334_ (.RESET_B(net5420),
    .D(_02030_),
    .Q(_00295_),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _22335_ (.RESET_B(net5420),
    .D(_02031_),
    .Q(_00296_),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _22336_ (.RESET_B(net5420),
    .D(_02032_),
    .Q(_00297_),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _22337_ (.RESET_B(net5420),
    .D(net1493),
    .Q(_00298_),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _22338_ (.RESET_B(net5448),
    .D(_02034_),
    .Q(_00299_),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _22339_ (.RESET_B(net5445),
    .D(_02035_),
    .Q(_00300_),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _22340_ (.RESET_B(net5445),
    .D(net1815),
    .Q(_00301_),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _22341_ (.RESET_B(net5414),
    .D(_02037_),
    .Q(_00302_),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _22342_ (.RESET_B(net5414),
    .D(net1488),
    .Q(_00303_),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _22343_ (.RESET_B(net5414),
    .D(_02039_),
    .Q(_00304_),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _22344_ (.RESET_B(net5418),
    .D(net1609),
    .Q(_00305_),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22345_ (.RESET_B(net5413),
    .D(_02041_),
    .Q(_00306_),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22346_ (.RESET_B(net5404),
    .D(net1362),
    .Q(_00307_),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _22347_ (.RESET_B(net5404),
    .D(net2009),
    .Q(_00308_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22348_ (.RESET_B(net5404),
    .D(net1133),
    .Q(_00309_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22349_ (.RESET_B(net5404),
    .D(_02045_),
    .Q(_00310_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22350_ (.RESET_B(net5405),
    .D(net1218),
    .Q(_00311_),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _22351_ (.RESET_B(net5405),
    .D(net1740),
    .Q(_00312_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22352_ (.RESET_B(net5405),
    .D(_02048_),
    .Q(_00313_),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _22353_ (.RESET_B(net5413),
    .D(net1022),
    .Q(_00314_),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _22354_ (.RESET_B(net5405),
    .D(net1497),
    .Q(_00315_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22355_ (.RESET_B(net5404),
    .D(net1926),
    .Q(_00316_),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _22356_ (.RESET_B(net5413),
    .D(net1390),
    .Q(_00317_),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _22357_ (.RESET_B(net5405),
    .D(net1857),
    .Q(_00318_),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _22358_ (.RESET_B(net5442),
    .D(_02054_),
    .Q(_00319_),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _22359_ (.RESET_B(net5441),
    .D(net2305),
    .Q(_00320_),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _22360_ (.RESET_B(net5441),
    .D(net533),
    .Q(_00321_),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _22361_ (.RESET_B(net5441),
    .D(net481),
    .Q(_00322_),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _22362_ (.RESET_B(net5442),
    .D(net611),
    .Q(_00323_),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _22363_ (.RESET_B(net5441),
    .D(net2312),
    .Q(_00324_),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _22364_ (.RESET_B(net5441),
    .D(net384),
    .Q(_00325_),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _22365_ (.RESET_B(net5441),
    .D(net423),
    .Q(_00326_),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _22366_ (.RESET_B(net5472),
    .D(_00168_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _22367_ (.RESET_B(net5483),
    .D(_02062_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[0] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _22368_ (.RESET_B(net5480),
    .D(_02063_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[1] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _22369_ (.RESET_B(net5481),
    .D(_02064_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[2] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _22370_ (.RESET_B(net5482),
    .D(_02065_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _22371_ (.RESET_B(net5482),
    .D(_02066_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _22372_ (.RESET_B(net5483),
    .D(_02067_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[5] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _22373_ (.RESET_B(net5482),
    .D(_02068_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _22374_ (.RESET_B(net5483),
    .D(_02069_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[7] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _22375_ (.RESET_B(net5448),
    .D(_00167_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _22376_ (.RESET_B(net5465),
    .D(_00166_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_rx_break_reg ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _22377_ (.RESET_B(net56),
    .D(_02070_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[7] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _22378_ (.RESET_B(net54),
    .D(net519),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[0] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _22379_ (.RESET_B(net52),
    .D(net1802),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[1] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _22380_ (.RESET_B(net50),
    .D(net2060),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _22381_ (.RESET_B(net47),
    .D(net871),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _22382_ (.RESET_B(net43),
    .D(_02075_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _22383_ (.RESET_B(net39),
    .D(_02076_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _22384_ (.RESET_B(net35),
    .D(net1450),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _22385_ (.RESET_B(net33),
    .D(_02078_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _22386_ (.RESET_B(net31),
    .D(net1366),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _22387_ (.RESET_B(net30),
    .D(_02080_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _22388_ (.RESET_B(net28),
    .D(net1313),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _22389_ (.RESET_B(net26),
    .D(_02082_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _22390_ (.RESET_B(net24),
    .D(_02083_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _22391_ (.RESET_B(net22),
    .D(_02084_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _22392_ (.RESET_B(net5469),
    .D(_02085_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _22393_ (.RESET_B(net5473),
    .D(_02086_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22394_ (.RESET_B(net5469),
    .D(net2653),
    .Q(_00327_),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22395_ (.RESET_B(net5436),
    .D(net2767),
    .Q(_00328_),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _22396_ (.RESET_B(net5469),
    .D(_02089_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _22397_ (.RESET_B(net5469),
    .D(_02090_),
    .Q(_00329_),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _22398_ (.RESET_B(net5436),
    .D(net2104),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _22399_ (.RESET_B(net5469),
    .D(_02092_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _22400_ (.RESET_B(net5435),
    .D(_02093_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _22401_ (.RESET_B(net5435),
    .D(_02094_),
    .Q(_00330_),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _22402_ (.RESET_B(net69),
    .D(_02095_),
    .Q(\soc_inst.uart_tx [0]),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _22403_ (.RESET_B(net5328),
    .D(_02096_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[13] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _22404_ (.RESET_B(net5350),
    .D(net2048),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[14] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _22405_ (.RESET_B(net5336),
    .D(_02098_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _22406_ (.RESET_B(net5338),
    .D(net2100),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[16] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _22407_ (.RESET_B(net5338),
    .D(net2003),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[17] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _22408_ (.RESET_B(net5317),
    .D(net2071),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[18] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _22409_ (.RESET_B(net5317),
    .D(net2013),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[19] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _22410_ (.RESET_B(net5335),
    .D(_02103_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[20] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _22411_ (.RESET_B(net5334),
    .D(_02104_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[21] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _22412_ (.RESET_B(net5334),
    .D(net2232),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[22] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _22413_ (.RESET_B(net5315),
    .D(net2121),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[23] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _22414_ (.RESET_B(net5348),
    .D(net473),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[24] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _22415_ (.RESET_B(net5339),
    .D(net2058),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[25] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _22416_ (.RESET_B(net5349),
    .D(net2110),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[26] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _22417_ (.RESET_B(net5339),
    .D(net2064),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[27] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _22418_ (.RESET_B(net5339),
    .D(net2437),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[28] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _22419_ (.RESET_B(net5339),
    .D(net1938),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[29] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _22420_ (.RESET_B(net5342),
    .D(net2411),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[30] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _22421_ (.RESET_B(net5348),
    .D(net2234),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[31] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _22422_ (.RESET_B(net65),
    .D(net606),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _22423_ (.RESET_B(net63),
    .D(net659),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _22424_ (.RESET_B(net62),
    .D(net1020),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _22425_ (.RESET_B(net60),
    .D(net663),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _22426_ (.RESET_B(net58),
    .D(net680),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _22427_ (.RESET_B(net55),
    .D(net1992),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _22428_ (.RESET_B(net51),
    .D(net1300),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _22429_ (.RESET_B(net45),
    .D(net1277),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _22430_ (.RESET_B(net37),
    .D(_02123_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[0] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _22431_ (.RESET_B(net32),
    .D(net1116),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[1] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _22432_ (.RESET_B(net29),
    .D(_02125_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[2] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _22433_ (.RESET_B(net25),
    .D(net657),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[3] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _22434_ (.RESET_B(net21),
    .D(net598),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[4] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _22435_ (.RESET_B(net19),
    .D(_02128_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _22436_ (.RESET_B(net17),
    .D(_02129_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[6] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _22437_ (.RESET_B(net15),
    .D(_02130_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _22438_ (.RESET_B(net74),
    .D(_02131_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _22439_ (.RESET_B(net64),
    .D(net524),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _22440_ (.RESET_B(net61),
    .D(_02133_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _22441_ (.RESET_B(net57),
    .D(_02134_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[3] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _22442_ (.RESET_B(net49),
    .D(net1699),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_sample ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _22443_ (.RESET_B(net34),
    .D(_02136_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22444_ (.RESET_B(net27),
    .D(net2182),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22445_ (.RESET_B(net20),
    .D(_02138_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _22446_ (.RESET_B(net16),
    .D(_02139_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _22447_ (.RESET_B(net66),
    .D(_02140_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _22448_ (.RESET_B(net59),
    .D(_02141_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _22449_ (.RESET_B(net41),
    .D(net2134),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _22450_ (.RESET_B(net23),
    .D(_02143_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _22451_ (.RESET_B(net14),
    .D(_02144_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _22452_ (.RESET_B(net53),
    .D(_02145_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _22453_ (.RESET_B(net18),
    .D(_02146_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg_0 ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _22454_ (.RESET_B(net75),
    .D(net571),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _22455_ (.RESET_B(net5476),
    .D(net491),
    .Q(\soc_inst.spi_inst.clk_counter[0] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _22456_ (.RESET_B(net5476),
    .D(net495),
    .Q(\soc_inst.spi_inst.clk_counter[1] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _22457_ (.RESET_B(net5475),
    .D(net585),
    .Q(\soc_inst.spi_inst.clk_counter[2] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _22458_ (.RESET_B(net5475),
    .D(net1919),
    .Q(\soc_inst.spi_inst.clk_counter[3] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _22459_ (.RESET_B(net5475),
    .D(net1936),
    .Q(\soc_inst.spi_inst.clk_counter[4] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _22460_ (.RESET_B(net5475),
    .D(net2379),
    .Q(\soc_inst.spi_inst.clk_counter[5] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _22461_ (.RESET_B(net5476),
    .D(net1995),
    .Q(\soc_inst.spi_inst.clk_counter[6] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _22462_ (.RESET_B(net5475),
    .D(net503),
    .Q(\soc_inst.spi_inst.clk_counter[7] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_tiehi _22437__15 (.L_HI(net15));
 sg13g2_tiehi _22446__16 (.L_HI(net16));
 sg13g2_tiehi _22436__17 (.L_HI(net17));
 sg13g2_tiehi _22453__18 (.L_HI(net18));
 sg13g2_tiehi _22435__19 (.L_HI(net19));
 sg13g2_tiehi _22445__20 (.L_HI(net20));
 sg13g2_tiehi _22434__21 (.L_HI(net21));
 sg13g2_tiehi _22391__22 (.L_HI(net22));
 sg13g2_tiehi _22450__23 (.L_HI(net23));
 sg13g2_tiehi _22390__24 (.L_HI(net24));
 sg13g2_tiehi _22433__25 (.L_HI(net25));
 sg13g2_tiehi _22389__26 (.L_HI(net26));
 sg13g2_tiehi _22444__27 (.L_HI(net27));
 sg13g2_tiehi _22388__28 (.L_HI(net28));
 sg13g2_tiehi _22432__29 (.L_HI(net29));
 sg13g2_tiehi _22387__30 (.L_HI(net30));
 sg13g2_tiehi _22386__31 (.L_HI(net31));
 sg13g2_tiehi _22431__32 (.L_HI(net32));
 sg13g2_tiehi _22385__33 (.L_HI(net33));
 sg13g2_tiehi _22443__34 (.L_HI(net34));
 sg13g2_tiehi _22384__35 (.L_HI(net35));
 sg13g2_tiehi _22332__36 (.L_HI(net36));
 sg13g2_tiehi _22430__37 (.L_HI(net37));
 sg13g2_tiehi _22327__38 (.L_HI(net38));
 sg13g2_tiehi _22383__39 (.L_HI(net39));
 sg13g2_tiehi _22326__40 (.L_HI(net40));
 sg13g2_tiehi _22449__41 (.L_HI(net41));
 sg13g2_tiehi _22325__42 (.L_HI(net42));
 sg13g2_tiehi _22382__43 (.L_HI(net43));
 sg13g2_tiehi _22324__44 (.L_HI(net44));
 sg13g2_tiehi _22429__45 (.L_HI(net45));
 sg13g2_tiehi _22323__46 (.L_HI(net46));
 sg13g2_tiehi _22381__47 (.L_HI(net47));
 sg13g2_tiehi _22322__48 (.L_HI(net48));
 sg13g2_tiehi _22442__49 (.L_HI(net49));
 sg13g2_tiehi _22380__50 (.L_HI(net50));
 sg13g2_tiehi _22428__51 (.L_HI(net51));
 sg13g2_tiehi _22379__52 (.L_HI(net52));
 sg13g2_tiehi _22452__53 (.L_HI(net53));
 sg13g2_tiehi _22378__54 (.L_HI(net54));
 sg13g2_tiehi _22427__55 (.L_HI(net55));
 sg13g2_tiehi _22377__56 (.L_HI(net56));
 sg13g2_tiehi _22441__57 (.L_HI(net57));
 sg13g2_tiehi _22426__58 (.L_HI(net58));
 sg13g2_tiehi _22448__59 (.L_HI(net59));
 sg13g2_tiehi _22425__60 (.L_HI(net60));
 sg13g2_tiehi _22440__61 (.L_HI(net61));
 sg13g2_tiehi _22424__62 (.L_HI(net62));
 sg13g2_tiehi _22423__63 (.L_HI(net63));
 sg13g2_tiehi _22439__64 (.L_HI(net64));
 sg13g2_tiehi _22422__65 (.L_HI(net65));
 sg13g2_tiehi _22447__66 (.L_HI(net66));
 sg13g2_tiehi _21060__67 (.L_HI(net67));
 sg13g2_tiehi _21059__68 (.L_HI(net68));
 sg13g2_tiehi _22402__69 (.L_HI(net69));
 sg13g2_tiehi _22328__70 (.L_HI(net70));
 sg13g2_tiehi _22329__71 (.L_HI(net71));
 sg13g2_tiehi _22330__72 (.L_HI(net72));
 sg13g2_tiehi _22331__73 (.L_HI(net73));
 sg13g2_tiehi _22438__74 (.L_HI(net74));
 sg13g2_tiehi _22454__75 (.L_HI(net75));
 sg13g2_tiehi tt_um_SotaSoC_76 (.L_HI(net76));
 sg13g2_tiehi tt_um_SotaSoC_77 (.L_HI(net77));
 sg13g2_tiehi tt_um_SotaSoC_78 (.L_HI(net78));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 _22528_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_8 _22529_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_8 _22530_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_8 _22531_ (.A(\soc_inst.flash_cs_n ),
    .X(uio_out[0]));
 sg13g2_buf_8 _22532_ (.A(\soc_inst.bus_spi_sclk ),
    .X(uio_out[3]));
 sg13g2_buf_8 _22533_ (.A(\soc_inst.mem_ctrl.ram_cs_n ),
    .X(uio_out[6]));
 sg13g2_buf_8 _22534_ (.A(\soc_inst.cpu_core.error_flag_reg ),
    .X(uo_out[0]));
 sg13g2_buf_16 _22535_ (.X(uo_out[1]),
    .A(\soc_inst.uart_tx [0]));
 sg13g2_buf_16 _22536_ (.X(uo_out[3]),
    .A(\soc_inst.gpio_inst.gpio_out[1] ));
 sg13g2_buf_8 fanout3683 (.A(net3685),
    .X(net3683));
 sg13g2_buf_8 fanout3684 (.A(net3685),
    .X(net3684));
 sg13g2_buf_8 fanout3685 (.A(net3686),
    .X(net3685));
 sg13g2_buf_2 fanout3686 (.A(net3689),
    .X(net3686));
 sg13g2_buf_8 fanout3687 (.A(net3688),
    .X(net3687));
 sg13g2_buf_8 fanout3688 (.A(net3689),
    .X(net3688));
 sg13g2_buf_2 fanout3689 (.A(_08318_),
    .X(net3689));
 sg13g2_buf_8 fanout3690 (.A(net3691),
    .X(net3690));
 sg13g2_buf_2 fanout3691 (.A(net3693),
    .X(net3691));
 sg13g2_buf_8 fanout3692 (.A(net3693),
    .X(net3692));
 sg13g2_buf_1 fanout3693 (.A(_08318_),
    .X(net3693));
 sg13g2_buf_8 fanout3694 (.A(net3695),
    .X(net3694));
 sg13g2_buf_8 fanout3695 (.A(net3697),
    .X(net3695));
 sg13g2_buf_8 fanout3696 (.A(net3697),
    .X(net3696));
 sg13g2_buf_8 fanout3697 (.A(net3700),
    .X(net3697));
 sg13g2_buf_8 fanout3698 (.A(net3699),
    .X(net3698));
 sg13g2_buf_8 fanout3699 (.A(net3700),
    .X(net3699));
 sg13g2_buf_8 fanout3700 (.A(_07718_),
    .X(net3700));
 sg13g2_buf_8 fanout3701 (.A(net3702),
    .X(net3701));
 sg13g2_buf_2 fanout3702 (.A(net3703),
    .X(net3702));
 sg13g2_buf_8 fanout3703 (.A(_07718_),
    .X(net3703));
 sg13g2_buf_8 fanout3704 (.A(net3705),
    .X(net3704));
 sg13g2_buf_2 fanout3705 (.A(net3706),
    .X(net3705));
 sg13g2_buf_1 fanout3706 (.A(_07667_),
    .X(net3706));
 sg13g2_buf_8 fanout3707 (.A(net3711),
    .X(net3707));
 sg13g2_buf_2 fanout3708 (.A(net3709),
    .X(net3708));
 sg13g2_buf_8 fanout3709 (.A(net3710),
    .X(net3709));
 sg13g2_buf_8 fanout3710 (.A(net3711),
    .X(net3710));
 sg13g2_buf_2 fanout3711 (.A(_07667_),
    .X(net3711));
 sg13g2_buf_8 fanout3712 (.A(_04408_),
    .X(net3712));
 sg13g2_buf_1 fanout3713 (.A(_04408_),
    .X(net3713));
 sg13g2_buf_8 fanout3714 (.A(net3715),
    .X(net3714));
 sg13g2_buf_8 fanout3715 (.A(_04326_),
    .X(net3715));
 sg13g2_buf_8 fanout3716 (.A(net3717),
    .X(net3716));
 sg13g2_buf_8 fanout3717 (.A(_06594_),
    .X(net3717));
 sg13g2_buf_8 fanout3718 (.A(net3719),
    .X(net3718));
 sg13g2_buf_8 fanout3719 (.A(_04996_),
    .X(net3719));
 sg13g2_buf_8 fanout3720 (.A(_09250_),
    .X(net3720));
 sg13g2_buf_8 fanout3721 (.A(_09250_),
    .X(net3721));
 sg13g2_buf_8 fanout3722 (.A(net3723),
    .X(net3722));
 sg13g2_buf_8 fanout3723 (.A(net3729),
    .X(net3723));
 sg13g2_buf_8 fanout3724 (.A(net3728),
    .X(net3724));
 sg13g2_buf_1 fanout3725 (.A(net3728),
    .X(net3725));
 sg13g2_buf_8 fanout3726 (.A(net3727),
    .X(net3726));
 sg13g2_buf_2 fanout3727 (.A(net3728),
    .X(net3727));
 sg13g2_buf_8 fanout3728 (.A(net3729),
    .X(net3728));
 sg13g2_buf_8 fanout3729 (.A(_09249_),
    .X(net3729));
 sg13g2_buf_8 fanout3730 (.A(net3733),
    .X(net3730));
 sg13g2_buf_1 fanout3731 (.A(net3733),
    .X(net3731));
 sg13g2_buf_2 fanout3732 (.A(net3733),
    .X(net3732));
 sg13g2_buf_8 fanout3733 (.A(_08782_),
    .X(net3733));
 sg13g2_buf_8 fanout3734 (.A(_08782_),
    .X(net3734));
 sg13g2_buf_1 fanout3735 (.A(net3736),
    .X(net3735));
 sg13g2_buf_8 fanout3736 (.A(_08782_),
    .X(net3736));
 sg13g2_buf_8 fanout3737 (.A(_06529_),
    .X(net3737));
 sg13g2_buf_8 fanout3738 (.A(_06529_),
    .X(net3738));
 sg13g2_buf_8 fanout3739 (.A(net3741),
    .X(net3739));
 sg13g2_buf_8 fanout3740 (.A(net3741),
    .X(net3740));
 sg13g2_buf_8 fanout3741 (.A(_04975_),
    .X(net3741));
 sg13g2_buf_8 fanout3742 (.A(_04801_),
    .X(net3742));
 sg13g2_buf_8 fanout3743 (.A(net3745),
    .X(net3743));
 sg13g2_buf_8 fanout3744 (.A(net3745),
    .X(net3744));
 sg13g2_buf_8 fanout3745 (.A(_04801_),
    .X(net3745));
 sg13g2_buf_8 fanout3746 (.A(_08470_),
    .X(net3746));
 sg13g2_buf_8 fanout3747 (.A(_08470_),
    .X(net3747));
 sg13g2_buf_8 fanout3748 (.A(net3750),
    .X(net3748));
 sg13g2_buf_8 fanout3749 (.A(net3750),
    .X(net3749));
 sg13g2_buf_8 fanout3750 (.A(_08469_),
    .X(net3750));
 sg13g2_buf_2 fanout3751 (.A(net3754),
    .X(net3751));
 sg13g2_buf_8 fanout3752 (.A(net3754),
    .X(net3752));
 sg13g2_buf_1 fanout3753 (.A(net3754),
    .X(net3753));
 sg13g2_buf_8 fanout3754 (.A(_06760_),
    .X(net3754));
 sg13g2_buf_8 fanout3755 (.A(_04994_),
    .X(net3755));
 sg13g2_buf_8 fanout3756 (.A(_04994_),
    .X(net3756));
 sg13g2_buf_8 fanout3757 (.A(net3761),
    .X(net3757));
 sg13g2_buf_8 fanout3758 (.A(net3761),
    .X(net3758));
 sg13g2_buf_8 fanout3759 (.A(net3760),
    .X(net3759));
 sg13g2_buf_8 fanout3760 (.A(net3761),
    .X(net3760));
 sg13g2_buf_8 fanout3761 (.A(_08466_),
    .X(net3761));
 sg13g2_buf_8 fanout3762 (.A(net3766),
    .X(net3762));
 sg13g2_buf_1 fanout3763 (.A(net3766),
    .X(net3763));
 sg13g2_buf_8 fanout3764 (.A(net3765),
    .X(net3764));
 sg13g2_buf_8 fanout3765 (.A(net3766),
    .X(net3765));
 sg13g2_buf_8 fanout3766 (.A(_07629_),
    .X(net3766));
 sg13g2_buf_8 fanout3767 (.A(net3769),
    .X(net3767));
 sg13g2_buf_8 fanout3768 (.A(net3769),
    .X(net3768));
 sg13g2_buf_8 fanout3769 (.A(net3778),
    .X(net3769));
 sg13g2_buf_8 fanout3770 (.A(net3778),
    .X(net3770));
 sg13g2_buf_8 fanout3771 (.A(net3776),
    .X(net3771));
 sg13g2_buf_2 fanout3772 (.A(net3776),
    .X(net3772));
 sg13g2_buf_8 fanout3773 (.A(net3774),
    .X(net3773));
 sg13g2_buf_8 fanout3774 (.A(net3776),
    .X(net3774));
 sg13g2_buf_1 fanout3775 (.A(net3776),
    .X(net3775));
 sg13g2_buf_2 fanout3776 (.A(net3777),
    .X(net3776));
 sg13g2_buf_8 fanout3777 (.A(net3778),
    .X(net3777));
 sg13g2_buf_8 fanout3778 (.A(_07531_),
    .X(net3778));
 sg13g2_buf_8 fanout3779 (.A(net3780),
    .X(net3779));
 sg13g2_buf_8 fanout3780 (.A(net3781),
    .X(net3780));
 sg13g2_buf_2 fanout3781 (.A(net3782),
    .X(net3781));
 sg13g2_buf_1 fanout3782 (.A(net3784),
    .X(net3782));
 sg13g2_buf_8 fanout3783 (.A(net3784),
    .X(net3783));
 sg13g2_buf_2 fanout3784 (.A(_07086_),
    .X(net3784));
 sg13g2_buf_8 fanout3785 (.A(net3786),
    .X(net3785));
 sg13g2_buf_8 fanout3786 (.A(_06817_),
    .X(net3786));
 sg13g2_buf_2 fanout3787 (.A(net3789),
    .X(net3787));
 sg13g2_buf_8 fanout3788 (.A(net3789),
    .X(net3788));
 sg13g2_buf_8 fanout3789 (.A(_06745_),
    .X(net3789));
 sg13g2_buf_2 fanout3790 (.A(net3791),
    .X(net3790));
 sg13g2_buf_1 fanout3791 (.A(net3792),
    .X(net3791));
 sg13g2_buf_8 fanout3792 (.A(net3797),
    .X(net3792));
 sg13g2_buf_8 fanout3793 (.A(net3794),
    .X(net3793));
 sg13g2_buf_8 fanout3794 (.A(net3795),
    .X(net3794));
 sg13g2_buf_8 fanout3795 (.A(net3796),
    .X(net3795));
 sg13g2_buf_8 fanout3796 (.A(net3797),
    .X(net3796));
 sg13g2_buf_8 fanout3797 (.A(_06658_),
    .X(net3797));
 sg13g2_buf_8 fanout3798 (.A(net3799),
    .X(net3798));
 sg13g2_buf_8 fanout3799 (.A(net3801),
    .X(net3799));
 sg13g2_buf_8 fanout3800 (.A(net3801),
    .X(net3800));
 sg13g2_buf_8 fanout3801 (.A(_06657_),
    .X(net3801));
 sg13g2_buf_2 fanout3802 (.A(net3803),
    .X(net3802));
 sg13g2_buf_8 fanout3803 (.A(net3805),
    .X(net3803));
 sg13g2_buf_2 fanout3804 (.A(net3805),
    .X(net3804));
 sg13g2_buf_1 fanout3805 (.A(_06657_),
    .X(net3805));
 sg13g2_buf_2 fanout3806 (.A(net3807),
    .X(net3806));
 sg13g2_buf_2 fanout3807 (.A(net3808),
    .X(net3807));
 sg13g2_buf_8 fanout3808 (.A(net3809),
    .X(net3808));
 sg13g2_buf_8 fanout3809 (.A(_07810_),
    .X(net3809));
 sg13g2_buf_2 fanout3810 (.A(net3814),
    .X(net3810));
 sg13g2_buf_2 fanout3811 (.A(net3813),
    .X(net3811));
 sg13g2_buf_1 fanout3812 (.A(net3813),
    .X(net3812));
 sg13g2_buf_1 fanout3813 (.A(net3814),
    .X(net3813));
 sg13g2_buf_1 fanout3814 (.A(net3816),
    .X(net3814));
 sg13g2_buf_8 fanout3815 (.A(net3816),
    .X(net3815));
 sg13g2_buf_8 fanout3816 (.A(_07809_),
    .X(net3816));
 sg13g2_buf_8 fanout3817 (.A(net3818),
    .X(net3817));
 sg13g2_buf_8 fanout3818 (.A(_07524_),
    .X(net3818));
 sg13g2_buf_8 fanout3819 (.A(_07508_),
    .X(net3819));
 sg13g2_buf_2 fanout3820 (.A(_07508_),
    .X(net3820));
 sg13g2_buf_8 fanout3821 (.A(net3823),
    .X(net3821));
 sg13g2_buf_1 fanout3822 (.A(net3823),
    .X(net3822));
 sg13g2_buf_2 fanout3823 (.A(_07500_),
    .X(net3823));
 sg13g2_buf_8 fanout3824 (.A(_07484_),
    .X(net3824));
 sg13g2_buf_8 fanout3825 (.A(_07484_),
    .X(net3825));
 sg13g2_buf_8 fanout3826 (.A(net3828),
    .X(net3826));
 sg13g2_buf_1 fanout3827 (.A(net3828),
    .X(net3827));
 sg13g2_buf_2 fanout3828 (.A(_07476_),
    .X(net3828));
 sg13g2_buf_8 fanout3829 (.A(net3830),
    .X(net3829));
 sg13g2_buf_8 fanout3830 (.A(_07468_),
    .X(net3830));
 sg13g2_buf_8 fanout3831 (.A(net3832),
    .X(net3831));
 sg13g2_buf_8 fanout3832 (.A(_07406_),
    .X(net3832));
 sg13g2_buf_8 fanout3833 (.A(net3834),
    .X(net3833));
 sg13g2_buf_8 fanout3834 (.A(_07350_),
    .X(net3834));
 sg13g2_buf_8 fanout3835 (.A(_07264_),
    .X(net3835));
 sg13g2_buf_8 fanout3836 (.A(_07264_),
    .X(net3836));
 sg13g2_buf_8 fanout3837 (.A(net3838),
    .X(net3837));
 sg13g2_buf_8 fanout3838 (.A(net3844),
    .X(net3838));
 sg13g2_buf_8 fanout3839 (.A(net3844),
    .X(net3839));
 sg13g2_buf_8 fanout3840 (.A(net3843),
    .X(net3840));
 sg13g2_buf_2 fanout3841 (.A(net3843),
    .X(net3841));
 sg13g2_buf_8 fanout3842 (.A(net3843),
    .X(net3842));
 sg13g2_buf_8 fanout3843 (.A(net3844),
    .X(net3843));
 sg13g2_buf_8 fanout3844 (.A(_06818_),
    .X(net3844));
 sg13g2_buf_2 fanout3845 (.A(net3846),
    .X(net3845));
 sg13g2_buf_8 fanout3846 (.A(_06796_),
    .X(net3846));
 sg13g2_buf_8 fanout3847 (.A(net3849),
    .X(net3847));
 sg13g2_buf_1 fanout3848 (.A(_06796_),
    .X(net3848));
 sg13g2_buf_8 fanout3849 (.A(_06796_),
    .X(net3849));
 sg13g2_buf_8 fanout3850 (.A(net3852),
    .X(net3850));
 sg13g2_buf_8 fanout3851 (.A(net3852),
    .X(net3851));
 sg13g2_buf_8 fanout3852 (.A(_06746_),
    .X(net3852));
 sg13g2_buf_8 fanout3853 (.A(net3854),
    .X(net3853));
 sg13g2_buf_8 fanout3854 (.A(net3856),
    .X(net3854));
 sg13g2_buf_8 fanout3855 (.A(net3856),
    .X(net3855));
 sg13g2_buf_8 fanout3856 (.A(_06720_),
    .X(net3856));
 sg13g2_buf_2 fanout3857 (.A(net3859),
    .X(net3857));
 sg13g2_buf_1 fanout3858 (.A(net3859),
    .X(net3858));
 sg13g2_buf_8 fanout3859 (.A(_06655_),
    .X(net3859));
 sg13g2_buf_8 fanout3860 (.A(net3863),
    .X(net3860));
 sg13g2_buf_8 fanout3861 (.A(net3862),
    .X(net3861));
 sg13g2_buf_8 fanout3862 (.A(net3863),
    .X(net3862));
 sg13g2_buf_8 fanout3863 (.A(_06654_),
    .X(net3863));
 sg13g2_buf_8 fanout3864 (.A(net3865),
    .X(net3864));
 sg13g2_buf_8 fanout3865 (.A(net3866),
    .X(net3865));
 sg13g2_buf_1 fanout3866 (.A(net3873),
    .X(net3866));
 sg13g2_buf_8 fanout3867 (.A(net3868),
    .X(net3867));
 sg13g2_buf_8 fanout3868 (.A(net3873),
    .X(net3868));
 sg13g2_buf_8 fanout3869 (.A(net3870),
    .X(net3869));
 sg13g2_buf_8 fanout3870 (.A(net3872),
    .X(net3870));
 sg13g2_buf_8 fanout3871 (.A(net3872),
    .X(net3871));
 sg13g2_buf_8 fanout3872 (.A(net3873),
    .X(net3872));
 sg13g2_buf_8 fanout3873 (.A(net3877),
    .X(net3873));
 sg13g2_buf_8 fanout3874 (.A(net3877),
    .X(net3874));
 sg13g2_buf_8 fanout3875 (.A(net3876),
    .X(net3875));
 sg13g2_buf_8 fanout3876 (.A(net3877),
    .X(net3876));
 sg13g2_buf_8 fanout3877 (.A(_06332_),
    .X(net3877));
 sg13g2_buf_8 fanout3878 (.A(net3879),
    .X(net3878));
 sg13g2_buf_8 fanout3879 (.A(_06331_),
    .X(net3879));
 sg13g2_buf_8 fanout3880 (.A(_02419_),
    .X(net3880));
 sg13g2_buf_8 fanout3881 (.A(_02399_),
    .X(net3881));
 sg13g2_buf_2 fanout3882 (.A(net3883),
    .X(net3882));
 sg13g2_buf_1 fanout3883 (.A(net3892),
    .X(net3883));
 sg13g2_buf_8 fanout3884 (.A(net3892),
    .X(net3884));
 sg13g2_buf_8 fanout3885 (.A(net3886),
    .X(net3885));
 sg13g2_buf_8 fanout3886 (.A(net3887),
    .X(net3886));
 sg13g2_buf_1 fanout3887 (.A(net3892),
    .X(net3887));
 sg13g2_buf_8 fanout3888 (.A(net3891),
    .X(net3888));
 sg13g2_buf_2 fanout3889 (.A(net3890),
    .X(net3889));
 sg13g2_buf_8 fanout3890 (.A(net3891),
    .X(net3890));
 sg13g2_buf_8 fanout3891 (.A(net3892),
    .X(net3891));
 sg13g2_buf_8 fanout3892 (.A(_09087_),
    .X(net3892));
 sg13g2_buf_8 fanout3893 (.A(_07516_),
    .X(net3893));
 sg13g2_buf_2 fanout3894 (.A(_07516_),
    .X(net3894));
 sg13g2_buf_8 fanout3895 (.A(_07492_),
    .X(net3895));
 sg13g2_buf_2 fanout3896 (.A(_07492_),
    .X(net3896));
 sg13g2_buf_8 fanout3897 (.A(net3898),
    .X(net3897));
 sg13g2_buf_1 fanout3898 (.A(net3899),
    .X(net3898));
 sg13g2_buf_1 fanout3899 (.A(_07460_),
    .X(net3899));
 sg13g2_buf_8 fanout3900 (.A(net3901),
    .X(net3900));
 sg13g2_buf_8 fanout3901 (.A(_07451_),
    .X(net3901));
 sg13g2_buf_8 fanout3902 (.A(net3903),
    .X(net3902));
 sg13g2_buf_8 fanout3903 (.A(_07442_),
    .X(net3903));
 sg13g2_buf_8 fanout3904 (.A(net3905),
    .X(net3904));
 sg13g2_buf_8 fanout3905 (.A(_07433_),
    .X(net3905));
 sg13g2_buf_8 fanout3906 (.A(net3908),
    .X(net3906));
 sg13g2_buf_1 fanout3907 (.A(net3908),
    .X(net3907));
 sg13g2_buf_1 fanout3908 (.A(_07424_),
    .X(net3908));
 sg13g2_buf_8 fanout3909 (.A(net3910),
    .X(net3909));
 sg13g2_buf_8 fanout3910 (.A(_07415_),
    .X(net3910));
 sg13g2_buf_8 fanout3911 (.A(net3913),
    .X(net3911));
 sg13g2_buf_1 fanout3912 (.A(net3913),
    .X(net3912));
 sg13g2_buf_8 fanout3913 (.A(_07397_),
    .X(net3913));
 sg13g2_buf_8 fanout3914 (.A(net3915),
    .X(net3914));
 sg13g2_buf_1 fanout3915 (.A(net3916),
    .X(net3915));
 sg13g2_buf_1 fanout3916 (.A(_07383_),
    .X(net3916));
 sg13g2_buf_8 fanout3917 (.A(_07372_),
    .X(net3917));
 sg13g2_buf_2 fanout3918 (.A(_07372_),
    .X(net3918));
 sg13g2_buf_8 fanout3919 (.A(net3921),
    .X(net3919));
 sg13g2_buf_1 fanout3920 (.A(net3921),
    .X(net3920));
 sg13g2_buf_2 fanout3921 (.A(_07361_),
    .X(net3921));
 sg13g2_buf_8 fanout3922 (.A(net3923),
    .X(net3922));
 sg13g2_buf_8 fanout3923 (.A(_07339_),
    .X(net3923));
 sg13g2_buf_8 fanout3924 (.A(net3925),
    .X(net3924));
 sg13g2_buf_8 fanout3925 (.A(_07327_),
    .X(net3925));
 sg13g2_buf_8 fanout3926 (.A(net3927),
    .X(net3926));
 sg13g2_buf_8 fanout3927 (.A(_07316_),
    .X(net3927));
 sg13g2_buf_8 fanout3928 (.A(net3929),
    .X(net3928));
 sg13g2_buf_8 fanout3929 (.A(_07305_),
    .X(net3929));
 sg13g2_buf_8 fanout3930 (.A(_07292_),
    .X(net3930));
 sg13g2_buf_8 fanout3931 (.A(_07292_),
    .X(net3931));
 sg13g2_buf_8 fanout3932 (.A(net3934),
    .X(net3932));
 sg13g2_buf_1 fanout3933 (.A(net3934),
    .X(net3933));
 sg13g2_buf_2 fanout3934 (.A(_07282_),
    .X(net3934));
 sg13g2_buf_8 fanout3935 (.A(net3937),
    .X(net3935));
 sg13g2_buf_1 fanout3936 (.A(net3937),
    .X(net3936));
 sg13g2_buf_8 fanout3937 (.A(_07273_),
    .X(net3937));
 sg13g2_buf_8 fanout3938 (.A(_07255_),
    .X(net3938));
 sg13g2_buf_1 fanout3939 (.A(_07255_),
    .X(net3939));
 sg13g2_buf_8 fanout3940 (.A(net3941),
    .X(net3940));
 sg13g2_buf_8 fanout3941 (.A(_07246_),
    .X(net3941));
 sg13g2_buf_8 fanout3942 (.A(net3943),
    .X(net3942));
 sg13g2_buf_8 fanout3943 (.A(_07236_),
    .X(net3943));
 sg13g2_buf_8 fanout3944 (.A(net3945),
    .X(net3944));
 sg13g2_buf_8 fanout3945 (.A(_07227_),
    .X(net3945));
 sg13g2_buf_8 fanout3946 (.A(_06718_),
    .X(net3946));
 sg13g2_buf_8 fanout3947 (.A(_06112_),
    .X(net3947));
 sg13g2_buf_8 fanout3948 (.A(net3949),
    .X(net3948));
 sg13g2_buf_2 fanout3949 (.A(_05332_),
    .X(net3949));
 sg13g2_buf_8 fanout3950 (.A(net3951),
    .X(net3950));
 sg13g2_buf_8 fanout3951 (.A(net3952),
    .X(net3951));
 sg13g2_buf_1 fanout3952 (.A(_05235_),
    .X(net3952));
 sg13g2_buf_8 fanout3953 (.A(net3956),
    .X(net3953));
 sg13g2_buf_8 fanout3954 (.A(net3955),
    .X(net3954));
 sg13g2_buf_2 fanout3955 (.A(net3956),
    .X(net3955));
 sg13g2_buf_1 fanout3956 (.A(net3957),
    .X(net3956));
 sg13g2_buf_2 fanout3957 (.A(net3958),
    .X(net3957));
 sg13g2_buf_8 fanout3958 (.A(_05172_),
    .X(net3958));
 sg13g2_buf_8 fanout3959 (.A(net3961),
    .X(net3959));
 sg13g2_buf_2 fanout3960 (.A(net3961),
    .X(net3960));
 sg13g2_buf_8 fanout3961 (.A(_05172_),
    .X(net3961));
 sg13g2_buf_2 fanout3962 (.A(net3963),
    .X(net3962));
 sg13g2_buf_1 fanout3963 (.A(_05172_),
    .X(net3963));
 sg13g2_buf_8 fanout3964 (.A(_05149_),
    .X(net3964));
 sg13g2_buf_8 fanout3965 (.A(net3966),
    .X(net3965));
 sg13g2_buf_2 fanout3966 (.A(net3969),
    .X(net3966));
 sg13g2_buf_8 fanout3967 (.A(net3969),
    .X(net3967));
 sg13g2_buf_8 fanout3968 (.A(net3969),
    .X(net3968));
 sg13g2_buf_8 fanout3969 (.A(_05118_),
    .X(net3969));
 sg13g2_buf_8 fanout3970 (.A(_02402_),
    .X(net3970));
 sg13g2_buf_8 fanout3971 (.A(net3972),
    .X(net3971));
 sg13g2_buf_8 fanout3972 (.A(_08401_),
    .X(net3972));
 sg13g2_buf_8 fanout3973 (.A(net3974),
    .X(net3973));
 sg13g2_buf_8 fanout3974 (.A(net3975),
    .X(net3974));
 sg13g2_buf_2 fanout3975 (.A(_08401_),
    .X(net3975));
 sg13g2_buf_8 fanout3976 (.A(_08226_),
    .X(net3976));
 sg13g2_buf_1 fanout3977 (.A(_08226_),
    .X(net3977));
 sg13g2_buf_8 fanout3978 (.A(_07929_),
    .X(net3978));
 sg13g2_buf_8 fanout3979 (.A(net3980),
    .X(net3979));
 sg13g2_buf_8 fanout3980 (.A(_07211_),
    .X(net3980));
 sg13g2_buf_2 fanout3981 (.A(net3982),
    .X(net3981));
 sg13g2_buf_8 fanout3982 (.A(_07133_),
    .X(net3982));
 sg13g2_buf_2 fanout3983 (.A(net3984),
    .X(net3983));
 sg13g2_buf_1 fanout3984 (.A(net3985),
    .X(net3984));
 sg13g2_buf_1 fanout3985 (.A(_07119_),
    .X(net3985));
 sg13g2_buf_8 fanout3986 (.A(net3987),
    .X(net3986));
 sg13g2_buf_8 fanout3987 (.A(_07070_),
    .X(net3987));
 sg13g2_buf_2 fanout3988 (.A(net3991),
    .X(net3988));
 sg13g2_buf_2 fanout3989 (.A(net3990),
    .X(net3989));
 sg13g2_buf_2 fanout3990 (.A(net3991),
    .X(net3990));
 sg13g2_buf_1 fanout3991 (.A(_06823_),
    .X(net3991));
 sg13g2_buf_2 fanout3992 (.A(net3995),
    .X(net3992));
 sg13g2_buf_2 fanout3993 (.A(net3994),
    .X(net3993));
 sg13g2_buf_2 fanout3994 (.A(net3995),
    .X(net3994));
 sg13g2_buf_1 fanout3995 (.A(_06643_),
    .X(net3995));
 sg13g2_buf_2 fanout3996 (.A(net3997),
    .X(net3996));
 sg13g2_buf_8 fanout3997 (.A(net4000),
    .X(net3997));
 sg13g2_buf_8 fanout3998 (.A(net4000),
    .X(net3998));
 sg13g2_buf_8 fanout3999 (.A(net4000),
    .X(net3999));
 sg13g2_buf_8 fanout4000 (.A(_06593_),
    .X(net4000));
 sg13g2_buf_8 fanout4001 (.A(net4005),
    .X(net4001));
 sg13g2_buf_8 fanout4002 (.A(net4005),
    .X(net4002));
 sg13g2_buf_8 fanout4003 (.A(net4005),
    .X(net4003));
 sg13g2_buf_8 fanout4004 (.A(net4005),
    .X(net4004));
 sg13g2_buf_8 fanout4005 (.A(_06527_),
    .X(net4005));
 sg13g2_buf_8 fanout4006 (.A(net4008),
    .X(net4006));
 sg13g2_buf_1 fanout4007 (.A(net4008),
    .X(net4007));
 sg13g2_buf_8 fanout4008 (.A(_06434_),
    .X(net4008));
 sg13g2_buf_8 fanout4009 (.A(net4010),
    .X(net4009));
 sg13g2_buf_8 fanout4010 (.A(_06306_),
    .X(net4010));
 sg13g2_buf_8 fanout4011 (.A(_06304_),
    .X(net4011));
 sg13g2_buf_1 fanout4012 (.A(_06304_),
    .X(net4012));
 sg13g2_buf_8 fanout4013 (.A(net4014),
    .X(net4013));
 sg13g2_buf_8 fanout4014 (.A(_06304_),
    .X(net4014));
 sg13g2_buf_8 fanout4015 (.A(net4017),
    .X(net4015));
 sg13g2_buf_8 fanout4016 (.A(net4017),
    .X(net4016));
 sg13g2_buf_8 fanout4017 (.A(net4018),
    .X(net4017));
 sg13g2_buf_8 fanout4018 (.A(_05904_),
    .X(net4018));
 sg13g2_buf_8 fanout4019 (.A(net4022),
    .X(net4019));
 sg13g2_buf_8 fanout4020 (.A(net4021),
    .X(net4020));
 sg13g2_buf_8 fanout4021 (.A(net4022),
    .X(net4021));
 sg13g2_buf_8 fanout4022 (.A(_02480_),
    .X(net4022));
 sg13g2_buf_8 fanout4023 (.A(_09011_),
    .X(net4023));
 sg13g2_buf_8 fanout4024 (.A(net4027),
    .X(net4024));
 sg13g2_buf_8 fanout4025 (.A(net4026),
    .X(net4025));
 sg13g2_buf_1 fanout4026 (.A(net4027),
    .X(net4026));
 sg13g2_buf_2 fanout4027 (.A(_08829_),
    .X(net4027));
 sg13g2_buf_8 fanout4028 (.A(net4030),
    .X(net4028));
 sg13g2_buf_1 fanout4029 (.A(net4030),
    .X(net4029));
 sg13g2_buf_1 fanout4030 (.A(net4031),
    .X(net4030));
 sg13g2_buf_1 fanout4031 (.A(_08829_),
    .X(net4031));
 sg13g2_buf_8 fanout4032 (.A(net4034),
    .X(net4032));
 sg13g2_buf_1 fanout4033 (.A(net4034),
    .X(net4033));
 sg13g2_buf_8 fanout4034 (.A(net4035),
    .X(net4034));
 sg13g2_buf_2 fanout4035 (.A(_08828_),
    .X(net4035));
 sg13g2_buf_8 fanout4036 (.A(net4037),
    .X(net4036));
 sg13g2_buf_8 fanout4037 (.A(_08400_),
    .X(net4037));
 sg13g2_buf_8 fanout4038 (.A(net4039),
    .X(net4038));
 sg13g2_buf_8 fanout4039 (.A(net4040),
    .X(net4039));
 sg13g2_buf_2 fanout4040 (.A(_08400_),
    .X(net4040));
 sg13g2_buf_8 fanout4041 (.A(net4042),
    .X(net4041));
 sg13g2_buf_8 fanout4042 (.A(_08096_),
    .X(net4042));
 sg13g2_buf_8 fanout4043 (.A(_07862_),
    .X(net4043));
 sg13g2_buf_8 fanout4044 (.A(_07847_),
    .X(net4044));
 sg13g2_buf_8 fanout4045 (.A(net4048),
    .X(net4045));
 sg13g2_buf_1 fanout4046 (.A(net4048),
    .X(net4046));
 sg13g2_buf_2 fanout4047 (.A(net4048),
    .X(net4047));
 sg13g2_buf_8 fanout4048 (.A(_07835_),
    .X(net4048));
 sg13g2_buf_2 fanout4049 (.A(_06651_),
    .X(net4049));
 sg13g2_buf_1 fanout4050 (.A(net4051),
    .X(net4050));
 sg13g2_buf_8 fanout4051 (.A(_06651_),
    .X(net4051));
 sg13g2_buf_8 fanout4052 (.A(net4053),
    .X(net4052));
 sg13g2_buf_8 fanout4053 (.A(net4054),
    .X(net4053));
 sg13g2_buf_1 fanout4054 (.A(_06651_),
    .X(net4054));
 sg13g2_buf_8 fanout4055 (.A(net4056),
    .X(net4055));
 sg13g2_buf_8 fanout4056 (.A(net4057),
    .X(net4056));
 sg13g2_buf_8 fanout4057 (.A(_06640_),
    .X(net4057));
 sg13g2_buf_8 fanout4058 (.A(net4059),
    .X(net4058));
 sg13g2_buf_8 fanout4059 (.A(_06639_),
    .X(net4059));
 sg13g2_buf_8 fanout4060 (.A(_06435_),
    .X(net4060));
 sg13g2_buf_8 fanout4061 (.A(net4062),
    .X(net4061));
 sg13g2_buf_1 fanout4062 (.A(net4065),
    .X(net4062));
 sg13g2_buf_8 fanout4063 (.A(net4064),
    .X(net4063));
 sg13g2_buf_1 fanout4064 (.A(net4065),
    .X(net4064));
 sg13g2_buf_1 fanout4065 (.A(_06301_),
    .X(net4065));
 sg13g2_buf_8 fanout4066 (.A(_05886_),
    .X(net4066));
 sg13g2_buf_8 fanout4067 (.A(_03379_),
    .X(net4067));
 sg13g2_buf_8 fanout4068 (.A(net4069),
    .X(net4068));
 sg13g2_buf_8 fanout4069 (.A(net4072),
    .X(net4069));
 sg13g2_buf_8 fanout4070 (.A(net4071),
    .X(net4070));
 sg13g2_buf_8 fanout4071 (.A(net4072),
    .X(net4071));
 sg13g2_buf_8 fanout4072 (.A(_02539_),
    .X(net4072));
 sg13g2_buf_8 fanout4073 (.A(_02365_),
    .X(net4073));
 sg13g2_buf_1 fanout4074 (.A(_02365_),
    .X(net4074));
 sg13g2_buf_8 fanout4075 (.A(net4079),
    .X(net4075));
 sg13g2_buf_8 fanout4076 (.A(net4079),
    .X(net4076));
 sg13g2_buf_8 fanout4077 (.A(net4078),
    .X(net4077));
 sg13g2_buf_8 fanout4078 (.A(net4079),
    .X(net4078));
 sg13g2_buf_8 fanout4079 (.A(_09988_),
    .X(net4079));
 sg13g2_buf_8 fanout4080 (.A(_09594_),
    .X(net4080));
 sg13g2_buf_2 fanout4081 (.A(_09594_),
    .X(net4081));
 sg13g2_buf_8 fanout4082 (.A(net4084),
    .X(net4082));
 sg13g2_buf_8 fanout4083 (.A(net4084),
    .X(net4083));
 sg13g2_buf_8 fanout4084 (.A(_09594_),
    .X(net4084));
 sg13g2_buf_8 fanout4085 (.A(net4086),
    .X(net4085));
 sg13g2_buf_2 fanout4086 (.A(net4087),
    .X(net4086));
 sg13g2_buf_2 fanout4087 (.A(_07387_),
    .X(net4087));
 sg13g2_buf_8 fanout4088 (.A(net4089),
    .X(net4088));
 sg13g2_buf_2 fanout4089 (.A(net4090),
    .X(net4089));
 sg13g2_buf_1 fanout4090 (.A(net4091),
    .X(net4090));
 sg13g2_buf_1 fanout4091 (.A(_06816_),
    .X(net4091));
 sg13g2_buf_8 fanout4092 (.A(net4094),
    .X(net4092));
 sg13g2_buf_8 fanout4093 (.A(net4094),
    .X(net4093));
 sg13g2_buf_8 fanout4094 (.A(_06816_),
    .X(net4094));
 sg13g2_buf_8 fanout4095 (.A(net4096),
    .X(net4095));
 sg13g2_buf_8 fanout4096 (.A(net4100),
    .X(net4096));
 sg13g2_buf_8 fanout4097 (.A(net4099),
    .X(net4097));
 sg13g2_buf_8 fanout4098 (.A(net4099),
    .X(net4098));
 sg13g2_buf_8 fanout4099 (.A(net4100),
    .X(net4099));
 sg13g2_buf_8 fanout4100 (.A(_06795_),
    .X(net4100));
 sg13g2_buf_8 fanout4101 (.A(net4103),
    .X(net4101));
 sg13g2_buf_8 fanout4102 (.A(net4103),
    .X(net4102));
 sg13g2_buf_8 fanout4103 (.A(_06642_),
    .X(net4103));
 sg13g2_buf_8 fanout4104 (.A(net4105),
    .X(net4104));
 sg13g2_buf_8 fanout4105 (.A(net4106),
    .X(net4105));
 sg13g2_buf_8 fanout4106 (.A(_06641_),
    .X(net4106));
 sg13g2_buf_8 fanout4107 (.A(net4108),
    .X(net4107));
 sg13g2_buf_2 fanout4108 (.A(_04298_),
    .X(net4108));
 sg13g2_buf_8 fanout4109 (.A(_04297_),
    .X(net4109));
 sg13g2_buf_1 fanout4110 (.A(_04297_),
    .X(net4110));
 sg13g2_buf_8 fanout4111 (.A(net4112),
    .X(net4111));
 sg13g2_buf_8 fanout4112 (.A(_02674_),
    .X(net4112));
 sg13g2_buf_8 fanout4113 (.A(net4114),
    .X(net4113));
 sg13g2_buf_8 fanout4114 (.A(net4115),
    .X(net4114));
 sg13g2_buf_1 fanout4115 (.A(_02477_),
    .X(net4115));
 sg13g2_buf_8 fanout4116 (.A(net4118),
    .X(net4116));
 sg13g2_buf_1 fanout4117 (.A(net4118),
    .X(net4117));
 sg13g2_buf_8 fanout4118 (.A(_02477_),
    .X(net4118));
 sg13g2_buf_8 fanout4119 (.A(_09231_),
    .X(net4119));
 sg13g2_buf_8 fanout4120 (.A(net4121),
    .X(net4120));
 sg13g2_buf_8 fanout4121 (.A(_09230_),
    .X(net4121));
 sg13g2_buf_8 fanout4122 (.A(net4123),
    .X(net4122));
 sg13g2_buf_8 fanout4123 (.A(net4124),
    .X(net4123));
 sg13g2_buf_8 fanout4124 (.A(_09211_),
    .X(net4124));
 sg13g2_buf_8 fanout4125 (.A(net4126),
    .X(net4125));
 sg13g2_buf_8 fanout4126 (.A(net4133),
    .X(net4126));
 sg13g2_buf_8 fanout4127 (.A(net4128),
    .X(net4127));
 sg13g2_buf_8 fanout4128 (.A(net4129),
    .X(net4128));
 sg13g2_buf_8 fanout4129 (.A(net4132),
    .X(net4129));
 sg13g2_buf_8 fanout4130 (.A(net4131),
    .X(net4130));
 sg13g2_buf_8 fanout4131 (.A(net4132),
    .X(net4131));
 sg13g2_buf_8 fanout4132 (.A(net4133),
    .X(net4132));
 sg13g2_buf_8 fanout4133 (.A(_09210_),
    .X(net4133));
 sg13g2_buf_8 fanout4134 (.A(net4135),
    .X(net4134));
 sg13g2_buf_8 fanout4135 (.A(_09089_),
    .X(net4135));
 sg13g2_buf_8 fanout4136 (.A(_08797_),
    .X(net4136));
 sg13g2_buf_1 fanout4137 (.A(_08797_),
    .X(net4137));
 sg13g2_buf_8 fanout4138 (.A(net4139),
    .X(net4138));
 sg13g2_buf_8 fanout4139 (.A(net4140),
    .X(net4139));
 sg13g2_buf_2 fanout4140 (.A(net4141),
    .X(net4140));
 sg13g2_buf_8 fanout4141 (.A(_08625_),
    .X(net4141));
 sg13g2_buf_8 fanout4142 (.A(net4143),
    .X(net4142));
 sg13g2_buf_8 fanout4143 (.A(_08597_),
    .X(net4143));
 sg13g2_buf_8 fanout4144 (.A(net4145),
    .X(net4144));
 sg13g2_buf_8 fanout4145 (.A(_08593_),
    .X(net4145));
 sg13g2_buf_8 fanout4146 (.A(_08593_),
    .X(net4146));
 sg13g2_buf_8 fanout4147 (.A(net4151),
    .X(net4147));
 sg13g2_buf_8 fanout4148 (.A(net4149),
    .X(net4148));
 sg13g2_buf_8 fanout4149 (.A(net4150),
    .X(net4149));
 sg13g2_buf_8 fanout4150 (.A(net4151),
    .X(net4150));
 sg13g2_buf_8 fanout4151 (.A(_08589_),
    .X(net4151));
 sg13g2_buf_8 fanout4152 (.A(net4153),
    .X(net4152));
 sg13g2_buf_8 fanout4153 (.A(_08587_),
    .X(net4153));
 sg13g2_buf_8 fanout4154 (.A(net4162),
    .X(net4154));
 sg13g2_buf_8 fanout4155 (.A(net4162),
    .X(net4155));
 sg13g2_buf_8 fanout4156 (.A(net4161),
    .X(net4156));
 sg13g2_buf_8 fanout4157 (.A(net4158),
    .X(net4157));
 sg13g2_buf_8 fanout4158 (.A(net4161),
    .X(net4158));
 sg13g2_buf_8 fanout4159 (.A(net4160),
    .X(net4159));
 sg13g2_buf_8 fanout4160 (.A(net4161),
    .X(net4160));
 sg13g2_buf_2 fanout4161 (.A(net4162),
    .X(net4161));
 sg13g2_buf_2 fanout4162 (.A(_08583_),
    .X(net4162));
 sg13g2_buf_8 fanout4163 (.A(net4164),
    .X(net4163));
 sg13g2_buf_1 fanout4164 (.A(net4165),
    .X(net4164));
 sg13g2_buf_8 fanout4165 (.A(net4166),
    .X(net4165));
 sg13g2_buf_8 fanout4166 (.A(_07669_),
    .X(net4166));
 sg13g2_buf_8 fanout4167 (.A(_07610_),
    .X(net4167));
 sg13g2_buf_1 fanout4168 (.A(_07610_),
    .X(net4168));
 sg13g2_buf_8 fanout4169 (.A(net4170),
    .X(net4169));
 sg13g2_buf_8 fanout4170 (.A(net4171),
    .X(net4170));
 sg13g2_buf_8 fanout4171 (.A(net4172),
    .X(net4171));
 sg13g2_buf_8 fanout4172 (.A(_07610_),
    .X(net4172));
 sg13g2_buf_8 fanout4173 (.A(_07607_),
    .X(net4173));
 sg13g2_buf_8 fanout4174 (.A(net4176),
    .X(net4174));
 sg13g2_buf_1 fanout4175 (.A(net4176),
    .X(net4175));
 sg13g2_buf_1 fanout4176 (.A(_07547_),
    .X(net4176));
 sg13g2_buf_8 fanout4177 (.A(_07295_),
    .X(net4177));
 sg13g2_buf_8 fanout4178 (.A(_07210_),
    .X(net4178));
 sg13g2_buf_8 fanout4179 (.A(_07210_),
    .X(net4179));
 sg13g2_buf_8 fanout4180 (.A(net4183),
    .X(net4180));
 sg13g2_buf_8 fanout4181 (.A(net4182),
    .X(net4181));
 sg13g2_buf_8 fanout4182 (.A(net4183),
    .X(net4182));
 sg13g2_buf_8 fanout4183 (.A(_06711_),
    .X(net4183));
 sg13g2_buf_8 fanout4184 (.A(net4188),
    .X(net4184));
 sg13g2_buf_1 fanout4185 (.A(net4188),
    .X(net4185));
 sg13g2_buf_8 fanout4186 (.A(net4188),
    .X(net4186));
 sg13g2_buf_8 fanout4187 (.A(net4188),
    .X(net4187));
 sg13g2_buf_8 fanout4188 (.A(_06697_),
    .X(net4188));
 sg13g2_buf_8 fanout4189 (.A(net4194),
    .X(net4189));
 sg13g2_buf_1 fanout4190 (.A(net4194),
    .X(net4190));
 sg13g2_buf_8 fanout4191 (.A(net4192),
    .X(net4191));
 sg13g2_buf_8 fanout4192 (.A(net4193),
    .X(net4192));
 sg13g2_buf_8 fanout4193 (.A(net4194),
    .X(net4193));
 sg13g2_buf_8 fanout4194 (.A(_06691_),
    .X(net4194));
 sg13g2_buf_8 fanout4195 (.A(net4198),
    .X(net4195));
 sg13g2_buf_1 fanout4196 (.A(net4198),
    .X(net4196));
 sg13g2_buf_8 fanout4197 (.A(net4198),
    .X(net4197));
 sg13g2_buf_8 fanout4198 (.A(_06627_),
    .X(net4198));
 sg13g2_buf_8 fanout4199 (.A(net4200),
    .X(net4199));
 sg13g2_buf_8 fanout4200 (.A(net4201),
    .X(net4200));
 sg13g2_buf_8 fanout4201 (.A(_06627_),
    .X(net4201));
 sg13g2_buf_8 fanout4202 (.A(_06472_),
    .X(net4202));
 sg13g2_buf_8 fanout4203 (.A(net4205),
    .X(net4203));
 sg13g2_buf_1 fanout4204 (.A(net4205),
    .X(net4204));
 sg13g2_buf_8 fanout4205 (.A(_06445_),
    .X(net4205));
 sg13g2_buf_8 fanout4206 (.A(_06297_),
    .X(net4206));
 sg13g2_buf_1 fanout4207 (.A(_06297_),
    .X(net4207));
 sg13g2_buf_8 fanout4208 (.A(_03406_),
    .X(net4208));
 sg13g2_buf_8 fanout4209 (.A(_03227_),
    .X(net4209));
 sg13g2_buf_8 fanout4210 (.A(_03017_),
    .X(net4210));
 sg13g2_buf_8 fanout4211 (.A(net4212),
    .X(net4211));
 sg13g2_buf_8 fanout4212 (.A(_02946_),
    .X(net4212));
 sg13g2_buf_8 fanout4213 (.A(net4214),
    .X(net4213));
 sg13g2_buf_8 fanout4214 (.A(_02910_),
    .X(net4214));
 sg13g2_buf_8 fanout4215 (.A(_02774_),
    .X(net4215));
 sg13g2_buf_8 fanout4216 (.A(net4217),
    .X(net4216));
 sg13g2_buf_8 fanout4217 (.A(_09229_),
    .X(net4217));
 sg13g2_buf_8 fanout4218 (.A(net4219),
    .X(net4218));
 sg13g2_buf_8 fanout4219 (.A(_08387_),
    .X(net4219));
 sg13g2_buf_8 fanout4220 (.A(net4221),
    .X(net4220));
 sg13g2_buf_8 fanout4221 (.A(_08386_),
    .X(net4221));
 sg13g2_buf_8 fanout4222 (.A(net4223),
    .X(net4222));
 sg13g2_buf_1 fanout4223 (.A(net4224),
    .X(net4223));
 sg13g2_buf_8 fanout4224 (.A(net4225),
    .X(net4224));
 sg13g2_buf_8 fanout4225 (.A(_07668_),
    .X(net4225));
 sg13g2_buf_8 fanout4226 (.A(net4227),
    .X(net4226));
 sg13g2_buf_8 fanout4227 (.A(_07385_),
    .X(net4227));
 sg13g2_buf_8 fanout4228 (.A(_07294_),
    .X(net4228));
 sg13g2_buf_8 fanout4229 (.A(net4230),
    .X(net4229));
 sg13g2_buf_8 fanout4230 (.A(net4231),
    .X(net4230));
 sg13g2_buf_8 fanout4231 (.A(_06751_),
    .X(net4231));
 sg13g2_buf_8 fanout4232 (.A(_06716_),
    .X(net4232));
 sg13g2_buf_8 fanout4233 (.A(net4234),
    .X(net4233));
 sg13g2_buf_1 fanout4234 (.A(net4235),
    .X(net4234));
 sg13g2_buf_8 fanout4235 (.A(net4236),
    .X(net4235));
 sg13g2_buf_8 fanout4236 (.A(_06709_),
    .X(net4236));
 sg13g2_buf_2 fanout4237 (.A(net4238),
    .X(net4237));
 sg13g2_buf_8 fanout4238 (.A(net4239),
    .X(net4238));
 sg13g2_buf_8 fanout4239 (.A(_06708_),
    .X(net4239));
 sg13g2_buf_8 fanout4240 (.A(net4241),
    .X(net4240));
 sg13g2_buf_8 fanout4241 (.A(net4246),
    .X(net4241));
 sg13g2_buf_2 fanout4242 (.A(net4243),
    .X(net4242));
 sg13g2_buf_8 fanout4243 (.A(net4246),
    .X(net4243));
 sg13g2_buf_8 fanout4244 (.A(net4245),
    .X(net4244));
 sg13g2_buf_8 fanout4245 (.A(net4246),
    .X(net4245));
 sg13g2_buf_8 fanout4246 (.A(_06680_),
    .X(net4246));
 sg13g2_buf_8 fanout4247 (.A(_06679_),
    .X(net4247));
 sg13g2_buf_8 fanout4248 (.A(_06679_),
    .X(net4248));
 sg13g2_buf_8 fanout4249 (.A(net4250),
    .X(net4249));
 sg13g2_buf_8 fanout4250 (.A(net4251),
    .X(net4250));
 sg13g2_buf_8 fanout4251 (.A(net4258),
    .X(net4251));
 sg13g2_buf_8 fanout4252 (.A(net4254),
    .X(net4252));
 sg13g2_buf_1 fanout4253 (.A(net4254),
    .X(net4253));
 sg13g2_buf_8 fanout4254 (.A(net4258),
    .X(net4254));
 sg13g2_buf_8 fanout4255 (.A(net4256),
    .X(net4255));
 sg13g2_buf_8 fanout4256 (.A(net4257),
    .X(net4256));
 sg13g2_buf_8 fanout4257 (.A(net4258),
    .X(net4257));
 sg13g2_buf_8 fanout4258 (.A(_06671_),
    .X(net4258));
 sg13g2_buf_8 fanout4259 (.A(_06591_),
    .X(net4259));
 sg13g2_buf_8 fanout4260 (.A(_06591_),
    .X(net4260));
 sg13g2_buf_8 fanout4261 (.A(_06524_),
    .X(net4261));
 sg13g2_buf_8 fanout4262 (.A(net4263),
    .X(net4262));
 sg13g2_buf_8 fanout4263 (.A(net4264),
    .X(net4263));
 sg13g2_buf_8 fanout4264 (.A(_06521_),
    .X(net4264));
 sg13g2_buf_8 fanout4265 (.A(net4268),
    .X(net4265));
 sg13g2_buf_8 fanout4266 (.A(net4268),
    .X(net4266));
 sg13g2_buf_8 fanout4267 (.A(net4268),
    .X(net4267));
 sg13g2_buf_8 fanout4268 (.A(_06433_),
    .X(net4268));
 sg13g2_buf_8 fanout4269 (.A(net4270),
    .X(net4269));
 sg13g2_buf_8 fanout4270 (.A(_06433_),
    .X(net4270));
 sg13g2_buf_8 fanout4271 (.A(net4272),
    .X(net4271));
 sg13g2_buf_8 fanout4272 (.A(_06432_),
    .X(net4272));
 sg13g2_buf_2 fanout4273 (.A(_06432_),
    .X(net4273));
 sg13g2_buf_8 fanout4274 (.A(net4276),
    .X(net4274));
 sg13g2_buf_1 fanout4275 (.A(net4276),
    .X(net4275));
 sg13g2_buf_8 fanout4276 (.A(_06429_),
    .X(net4276));
 sg13g2_buf_8 fanout4277 (.A(_06295_),
    .X(net4277));
 sg13g2_buf_8 fanout4278 (.A(_06047_),
    .X(net4278));
 sg13g2_buf_1 fanout4279 (.A(_06047_),
    .X(net4279));
 sg13g2_buf_8 fanout4280 (.A(_06046_),
    .X(net4280));
 sg13g2_buf_8 fanout4281 (.A(net4284),
    .X(net4281));
 sg13g2_buf_8 fanout4282 (.A(net4284),
    .X(net4282));
 sg13g2_buf_8 fanout4283 (.A(net4284),
    .X(net4283));
 sg13g2_buf_8 fanout4284 (.A(_04142_),
    .X(net4284));
 sg13g2_buf_8 fanout4285 (.A(net4286),
    .X(net4285));
 sg13g2_buf_8 fanout4286 (.A(net4287),
    .X(net4286));
 sg13g2_buf_8 fanout4287 (.A(_04142_),
    .X(net4287));
 sg13g2_buf_8 fanout4288 (.A(net4290),
    .X(net4288));
 sg13g2_buf_8 fanout4289 (.A(net4290),
    .X(net4289));
 sg13g2_buf_8 fanout4290 (.A(_04142_),
    .X(net4290));
 sg13g2_buf_8 fanout4291 (.A(net4292),
    .X(net4291));
 sg13g2_buf_8 fanout4292 (.A(net4295),
    .X(net4292));
 sg13g2_buf_8 fanout4293 (.A(net4295),
    .X(net4293));
 sg13g2_buf_8 fanout4294 (.A(net4295),
    .X(net4294));
 sg13g2_buf_8 fanout4295 (.A(_04109_),
    .X(net4295));
 sg13g2_buf_8 fanout4296 (.A(net4300),
    .X(net4296));
 sg13g2_buf_8 fanout4297 (.A(net4300),
    .X(net4297));
 sg13g2_buf_8 fanout4298 (.A(net4299),
    .X(net4298));
 sg13g2_buf_8 fanout4299 (.A(net4300),
    .X(net4299));
 sg13g2_buf_8 fanout4300 (.A(_04109_),
    .X(net4300));
 sg13g2_buf_8 fanout4301 (.A(net4305),
    .X(net4301));
 sg13g2_buf_8 fanout4302 (.A(net4305),
    .X(net4302));
 sg13g2_buf_8 fanout4303 (.A(net4305),
    .X(net4303));
 sg13g2_buf_8 fanout4304 (.A(net4305),
    .X(net4304));
 sg13g2_buf_8 fanout4305 (.A(_04076_),
    .X(net4305));
 sg13g2_buf_8 fanout4306 (.A(net4307),
    .X(net4306));
 sg13g2_buf_8 fanout4307 (.A(net4310),
    .X(net4307));
 sg13g2_buf_8 fanout4308 (.A(net4309),
    .X(net4308));
 sg13g2_buf_8 fanout4309 (.A(net4310),
    .X(net4309));
 sg13g2_buf_8 fanout4310 (.A(_04076_),
    .X(net4310));
 sg13g2_buf_8 fanout4311 (.A(net4315),
    .X(net4311));
 sg13g2_buf_8 fanout4312 (.A(net4315),
    .X(net4312));
 sg13g2_buf_8 fanout4313 (.A(net4315),
    .X(net4313));
 sg13g2_buf_8 fanout4314 (.A(net4315),
    .X(net4314));
 sg13g2_buf_8 fanout4315 (.A(net4321),
    .X(net4315));
 sg13g2_buf_8 fanout4316 (.A(net4318),
    .X(net4316));
 sg13g2_buf_1 fanout4317 (.A(net4318),
    .X(net4317));
 sg13g2_buf_8 fanout4318 (.A(net4321),
    .X(net4318));
 sg13g2_buf_8 fanout4319 (.A(net4321),
    .X(net4319));
 sg13g2_buf_8 fanout4320 (.A(net4321),
    .X(net4320));
 sg13g2_buf_8 fanout4321 (.A(_04043_),
    .X(net4321));
 sg13g2_buf_8 fanout4322 (.A(net4323),
    .X(net4322));
 sg13g2_buf_8 fanout4323 (.A(net4331),
    .X(net4323));
 sg13g2_buf_8 fanout4324 (.A(net4325),
    .X(net4324));
 sg13g2_buf_8 fanout4325 (.A(net4331),
    .X(net4325));
 sg13g2_buf_8 fanout4326 (.A(net4328),
    .X(net4326));
 sg13g2_buf_1 fanout4327 (.A(net4328),
    .X(net4327));
 sg13g2_buf_8 fanout4328 (.A(net4331),
    .X(net4328));
 sg13g2_buf_8 fanout4329 (.A(net4330),
    .X(net4329));
 sg13g2_buf_8 fanout4330 (.A(net4331),
    .X(net4330));
 sg13g2_buf_8 fanout4331 (.A(_04010_),
    .X(net4331));
 sg13g2_buf_8 fanout4332 (.A(net4333),
    .X(net4332));
 sg13g2_buf_8 fanout4333 (.A(net4336),
    .X(net4333));
 sg13g2_buf_8 fanout4334 (.A(net4336),
    .X(net4334));
 sg13g2_buf_8 fanout4335 (.A(net4336),
    .X(net4335));
 sg13g2_buf_8 fanout4336 (.A(_03977_),
    .X(net4336));
 sg13g2_buf_8 fanout4337 (.A(net4341),
    .X(net4337));
 sg13g2_buf_8 fanout4338 (.A(net4341),
    .X(net4338));
 sg13g2_buf_8 fanout4339 (.A(net4341),
    .X(net4339));
 sg13g2_buf_8 fanout4340 (.A(net4341),
    .X(net4340));
 sg13g2_buf_8 fanout4341 (.A(_03977_),
    .X(net4341));
 sg13g2_buf_8 fanout4342 (.A(net4346),
    .X(net4342));
 sg13g2_buf_8 fanout4343 (.A(net4346),
    .X(net4343));
 sg13g2_buf_8 fanout4344 (.A(net4345),
    .X(net4344));
 sg13g2_buf_8 fanout4345 (.A(net4346),
    .X(net4345));
 sg13g2_buf_8 fanout4346 (.A(_03944_),
    .X(net4346));
 sg13g2_buf_8 fanout4347 (.A(net4351),
    .X(net4347));
 sg13g2_buf_8 fanout4348 (.A(net4351),
    .X(net4348));
 sg13g2_buf_8 fanout4349 (.A(net4350),
    .X(net4349));
 sg13g2_buf_8 fanout4350 (.A(net4351),
    .X(net4350));
 sg13g2_buf_8 fanout4351 (.A(_03944_),
    .X(net4351));
 sg13g2_buf_8 fanout4352 (.A(net4356),
    .X(net4352));
 sg13g2_buf_8 fanout4353 (.A(net4356),
    .X(net4353));
 sg13g2_buf_8 fanout4354 (.A(net4355),
    .X(net4354));
 sg13g2_buf_8 fanout4355 (.A(net4356),
    .X(net4355));
 sg13g2_buf_8 fanout4356 (.A(_03910_),
    .X(net4356));
 sg13g2_buf_8 fanout4357 (.A(net4361),
    .X(net4357));
 sg13g2_buf_8 fanout4358 (.A(net4361),
    .X(net4358));
 sg13g2_buf_8 fanout4359 (.A(net4361),
    .X(net4359));
 sg13g2_buf_8 fanout4360 (.A(net4361),
    .X(net4360));
 sg13g2_buf_8 fanout4361 (.A(_03910_),
    .X(net4361));
 sg13g2_buf_8 fanout4362 (.A(net4363),
    .X(net4362));
 sg13g2_buf_8 fanout4363 (.A(net4366),
    .X(net4363));
 sg13g2_buf_8 fanout4364 (.A(net4365),
    .X(net4364));
 sg13g2_buf_8 fanout4365 (.A(net4366),
    .X(net4365));
 sg13g2_buf_8 fanout4366 (.A(net4372),
    .X(net4366));
 sg13g2_buf_8 fanout4367 (.A(net4369),
    .X(net4367));
 sg13g2_buf_1 fanout4368 (.A(net4369),
    .X(net4368));
 sg13g2_buf_8 fanout4369 (.A(net4372),
    .X(net4369));
 sg13g2_buf_8 fanout4370 (.A(net4372),
    .X(net4370));
 sg13g2_buf_2 fanout4371 (.A(net4372),
    .X(net4371));
 sg13g2_buf_8 fanout4372 (.A(_03877_),
    .X(net4372));
 sg13g2_buf_8 fanout4373 (.A(net4377),
    .X(net4373));
 sg13g2_buf_8 fanout4374 (.A(net4377),
    .X(net4374));
 sg13g2_buf_8 fanout4375 (.A(net4377),
    .X(net4375));
 sg13g2_buf_8 fanout4376 (.A(net4377),
    .X(net4376));
 sg13g2_buf_8 fanout4377 (.A(_03844_),
    .X(net4377));
 sg13g2_buf_8 fanout4378 (.A(net4382),
    .X(net4378));
 sg13g2_buf_8 fanout4379 (.A(net4382),
    .X(net4379));
 sg13g2_buf_8 fanout4380 (.A(net4382),
    .X(net4380));
 sg13g2_buf_1 fanout4381 (.A(net4382),
    .X(net4381));
 sg13g2_buf_8 fanout4382 (.A(_03844_),
    .X(net4382));
 sg13g2_buf_8 fanout4383 (.A(net4392),
    .X(net4383));
 sg13g2_buf_8 fanout4384 (.A(net4392),
    .X(net4384));
 sg13g2_buf_8 fanout4385 (.A(net4386),
    .X(net4385));
 sg13g2_buf_8 fanout4386 (.A(net4392),
    .X(net4386));
 sg13g2_buf_8 fanout4387 (.A(net4388),
    .X(net4387));
 sg13g2_buf_8 fanout4388 (.A(net4391),
    .X(net4388));
 sg13g2_buf_8 fanout4389 (.A(net4390),
    .X(net4389));
 sg13g2_buf_8 fanout4390 (.A(net4391),
    .X(net4390));
 sg13g2_buf_8 fanout4391 (.A(net4392),
    .X(net4391));
 sg13g2_buf_8 fanout4392 (.A(_03811_),
    .X(net4392));
 sg13g2_buf_8 fanout4393 (.A(net4394),
    .X(net4393));
 sg13g2_buf_8 fanout4394 (.A(net4397),
    .X(net4394));
 sg13g2_buf_8 fanout4395 (.A(net4396),
    .X(net4395));
 sg13g2_buf_8 fanout4396 (.A(net4397),
    .X(net4396));
 sg13g2_buf_8 fanout4397 (.A(_03777_),
    .X(net4397));
 sg13g2_buf_8 fanout4398 (.A(net4399),
    .X(net4398));
 sg13g2_buf_8 fanout4399 (.A(net4402),
    .X(net4399));
 sg13g2_buf_8 fanout4400 (.A(net4402),
    .X(net4400));
 sg13g2_buf_8 fanout4401 (.A(net4402),
    .X(net4401));
 sg13g2_buf_8 fanout4402 (.A(_03777_),
    .X(net4402));
 sg13g2_buf_8 fanout4403 (.A(net4407),
    .X(net4403));
 sg13g2_buf_8 fanout4404 (.A(net4407),
    .X(net4404));
 sg13g2_buf_8 fanout4405 (.A(net4406),
    .X(net4405));
 sg13g2_buf_8 fanout4406 (.A(net4407),
    .X(net4406));
 sg13g2_buf_8 fanout4407 (.A(_03744_),
    .X(net4407));
 sg13g2_buf_8 fanout4408 (.A(net4409),
    .X(net4408));
 sg13g2_buf_8 fanout4409 (.A(net4412),
    .X(net4409));
 sg13g2_buf_8 fanout4410 (.A(net4411),
    .X(net4410));
 sg13g2_buf_8 fanout4411 (.A(net4412),
    .X(net4411));
 sg13g2_buf_8 fanout4412 (.A(_03744_),
    .X(net4412));
 sg13g2_buf_8 fanout4413 (.A(net4423),
    .X(net4413));
 sg13g2_buf_2 fanout4414 (.A(net4423),
    .X(net4414));
 sg13g2_buf_8 fanout4415 (.A(net4416),
    .X(net4415));
 sg13g2_buf_8 fanout4416 (.A(net4423),
    .X(net4416));
 sg13g2_buf_8 fanout4417 (.A(net4422),
    .X(net4417));
 sg13g2_buf_8 fanout4418 (.A(net4422),
    .X(net4418));
 sg13g2_buf_8 fanout4419 (.A(net4421),
    .X(net4419));
 sg13g2_buf_1 fanout4420 (.A(net4421),
    .X(net4420));
 sg13g2_buf_8 fanout4421 (.A(net4422),
    .X(net4421));
 sg13g2_buf_8 fanout4422 (.A(net4423),
    .X(net4422));
 sg13g2_buf_8 fanout4423 (.A(_03710_),
    .X(net4423));
 sg13g2_buf_8 fanout4424 (.A(_03015_),
    .X(net4424));
 sg13g2_buf_8 fanout4425 (.A(net4427),
    .X(net4425));
 sg13g2_buf_8 fanout4426 (.A(net4427),
    .X(net4426));
 sg13g2_buf_8 fanout4427 (.A(_03014_),
    .X(net4427));
 sg13g2_buf_8 fanout4428 (.A(net4431),
    .X(net4428));
 sg13g2_buf_8 fanout4429 (.A(net4431),
    .X(net4429));
 sg13g2_buf_1 fanout4430 (.A(net4431),
    .X(net4430));
 sg13g2_buf_8 fanout4431 (.A(_03010_),
    .X(net4431));
 sg13g2_buf_8 fanout4432 (.A(_02949_),
    .X(net4432));
 sg13g2_buf_8 fanout4433 (.A(_02949_),
    .X(net4433));
 sg13g2_buf_8 fanout4434 (.A(net4436),
    .X(net4434));
 sg13g2_buf_8 fanout4435 (.A(net4436),
    .X(net4435));
 sg13g2_buf_8 fanout4436 (.A(_02948_),
    .X(net4436));
 sg13g2_buf_8 fanout4437 (.A(net4441),
    .X(net4437));
 sg13g2_buf_1 fanout4438 (.A(net4441),
    .X(net4438));
 sg13g2_buf_8 fanout4439 (.A(net4441),
    .X(net4439));
 sg13g2_buf_1 fanout4440 (.A(net4441),
    .X(net4440));
 sg13g2_buf_2 fanout4441 (.A(_02935_),
    .X(net4441));
 sg13g2_buf_8 fanout4442 (.A(_02830_),
    .X(net4442));
 sg13g2_buf_8 fanout4443 (.A(_02777_),
    .X(net4443));
 sg13g2_buf_8 fanout4444 (.A(_02671_),
    .X(net4444));
 sg13g2_buf_8 fanout4445 (.A(_02671_),
    .X(net4445));
 sg13g2_buf_8 fanout4446 (.A(net4447),
    .X(net4446));
 sg13g2_buf_8 fanout4447 (.A(_02670_),
    .X(net4447));
 sg13g2_buf_8 fanout4448 (.A(net4453),
    .X(net4448));
 sg13g2_buf_1 fanout4449 (.A(net4453),
    .X(net4449));
 sg13g2_buf_8 fanout4450 (.A(net4451),
    .X(net4450));
 sg13g2_buf_8 fanout4451 (.A(net4453),
    .X(net4451));
 sg13g2_buf_8 fanout4452 (.A(net4453),
    .X(net4452));
 sg13g2_buf_8 fanout4453 (.A(_02352_),
    .X(net4453));
 sg13g2_buf_8 fanout4454 (.A(net4458),
    .X(net4454));
 sg13g2_buf_8 fanout4455 (.A(net4458),
    .X(net4455));
 sg13g2_buf_8 fanout4456 (.A(net4458),
    .X(net4456));
 sg13g2_buf_8 fanout4457 (.A(net4458),
    .X(net4457));
 sg13g2_buf_8 fanout4458 (.A(_10014_),
    .X(net4458));
 sg13g2_buf_8 fanout4459 (.A(net4463),
    .X(net4459));
 sg13g2_buf_8 fanout4460 (.A(net4463),
    .X(net4460));
 sg13g2_buf_8 fanout4461 (.A(net4463),
    .X(net4461));
 sg13g2_buf_8 fanout4462 (.A(net4463),
    .X(net4462));
 sg13g2_buf_8 fanout4463 (.A(_10013_),
    .X(net4463));
 sg13g2_buf_8 fanout4464 (.A(net4468),
    .X(net4464));
 sg13g2_buf_8 fanout4465 (.A(net4468),
    .X(net4465));
 sg13g2_buf_8 fanout4466 (.A(net4468),
    .X(net4466));
 sg13g2_buf_8 fanout4467 (.A(net4468),
    .X(net4467));
 sg13g2_buf_8 fanout4468 (.A(_10012_),
    .X(net4468));
 sg13g2_buf_8 fanout4469 (.A(net4473),
    .X(net4469));
 sg13g2_buf_8 fanout4470 (.A(net4473),
    .X(net4470));
 sg13g2_buf_8 fanout4471 (.A(net4473),
    .X(net4471));
 sg13g2_buf_8 fanout4472 (.A(net4473),
    .X(net4472));
 sg13g2_buf_8 fanout4473 (.A(_10011_),
    .X(net4473));
 sg13g2_buf_8 fanout4474 (.A(net4478),
    .X(net4474));
 sg13g2_buf_8 fanout4475 (.A(net4478),
    .X(net4475));
 sg13g2_buf_8 fanout4476 (.A(net4478),
    .X(net4476));
 sg13g2_buf_8 fanout4477 (.A(net4478),
    .X(net4477));
 sg13g2_buf_8 fanout4478 (.A(_10010_),
    .X(net4478));
 sg13g2_buf_8 fanout4479 (.A(net4483),
    .X(net4479));
 sg13g2_buf_8 fanout4480 (.A(net4483),
    .X(net4480));
 sg13g2_buf_8 fanout4481 (.A(net4483),
    .X(net4481));
 sg13g2_buf_8 fanout4482 (.A(net4483),
    .X(net4482));
 sg13g2_buf_8 fanout4483 (.A(_10009_),
    .X(net4483));
 sg13g2_buf_8 fanout4484 (.A(net4488),
    .X(net4484));
 sg13g2_buf_8 fanout4485 (.A(net4488),
    .X(net4485));
 sg13g2_buf_8 fanout4486 (.A(net4487),
    .X(net4486));
 sg13g2_buf_8 fanout4487 (.A(net4488),
    .X(net4487));
 sg13g2_buf_8 fanout4488 (.A(_10008_),
    .X(net4488));
 sg13g2_buf_8 fanout4489 (.A(net4493),
    .X(net4489));
 sg13g2_buf_8 fanout4490 (.A(net4493),
    .X(net4490));
 sg13g2_buf_8 fanout4491 (.A(net4492),
    .X(net4491));
 sg13g2_buf_8 fanout4492 (.A(net4493),
    .X(net4492));
 sg13g2_buf_8 fanout4493 (.A(_10006_),
    .X(net4493));
 sg13g2_buf_8 fanout4494 (.A(net4498),
    .X(net4494));
 sg13g2_buf_8 fanout4495 (.A(net4498),
    .X(net4495));
 sg13g2_buf_8 fanout4496 (.A(net4498),
    .X(net4496));
 sg13g2_buf_8 fanout4497 (.A(net4498),
    .X(net4497));
 sg13g2_buf_8 fanout4498 (.A(_10004_),
    .X(net4498));
 sg13g2_buf_8 fanout4499 (.A(net4503),
    .X(net4499));
 sg13g2_buf_8 fanout4500 (.A(net4503),
    .X(net4500));
 sg13g2_buf_8 fanout4501 (.A(net4503),
    .X(net4501));
 sg13g2_buf_8 fanout4502 (.A(net4503),
    .X(net4502));
 sg13g2_buf_8 fanout4503 (.A(_10003_),
    .X(net4503));
 sg13g2_buf_8 fanout4504 (.A(net4508),
    .X(net4504));
 sg13g2_buf_8 fanout4505 (.A(net4508),
    .X(net4505));
 sg13g2_buf_8 fanout4506 (.A(net4508),
    .X(net4506));
 sg13g2_buf_8 fanout4507 (.A(net4508),
    .X(net4507));
 sg13g2_buf_8 fanout4508 (.A(_10002_),
    .X(net4508));
 sg13g2_buf_8 fanout4509 (.A(net4513),
    .X(net4509));
 sg13g2_buf_8 fanout4510 (.A(net4513),
    .X(net4510));
 sg13g2_buf_8 fanout4511 (.A(net4513),
    .X(net4511));
 sg13g2_buf_8 fanout4512 (.A(net4513),
    .X(net4512));
 sg13g2_buf_8 fanout4513 (.A(_10000_),
    .X(net4513));
 sg13g2_buf_8 fanout4514 (.A(net4518),
    .X(net4514));
 sg13g2_buf_8 fanout4515 (.A(net4518),
    .X(net4515));
 sg13g2_buf_8 fanout4516 (.A(net4518),
    .X(net4516));
 sg13g2_buf_8 fanout4517 (.A(net4518),
    .X(net4517));
 sg13g2_buf_8 fanout4518 (.A(_09996_),
    .X(net4518));
 sg13g2_buf_8 fanout4519 (.A(net4523),
    .X(net4519));
 sg13g2_buf_8 fanout4520 (.A(net4523),
    .X(net4520));
 sg13g2_buf_8 fanout4521 (.A(net4523),
    .X(net4521));
 sg13g2_buf_8 fanout4522 (.A(net4523),
    .X(net4522));
 sg13g2_buf_8 fanout4523 (.A(_09994_),
    .X(net4523));
 sg13g2_buf_8 fanout4524 (.A(net4528),
    .X(net4524));
 sg13g2_buf_8 fanout4525 (.A(net4528),
    .X(net4525));
 sg13g2_buf_8 fanout4526 (.A(net4528),
    .X(net4526));
 sg13g2_buf_8 fanout4527 (.A(net4528),
    .X(net4527));
 sg13g2_buf_8 fanout4528 (.A(_09616_),
    .X(net4528));
 sg13g2_buf_8 fanout4529 (.A(net4533),
    .X(net4529));
 sg13g2_buf_8 fanout4530 (.A(net4533),
    .X(net4530));
 sg13g2_buf_8 fanout4531 (.A(net4533),
    .X(net4531));
 sg13g2_buf_8 fanout4532 (.A(net4533),
    .X(net4532));
 sg13g2_buf_8 fanout4533 (.A(_09615_),
    .X(net4533));
 sg13g2_buf_8 fanout4534 (.A(net4538),
    .X(net4534));
 sg13g2_buf_8 fanout4535 (.A(net4538),
    .X(net4535));
 sg13g2_buf_8 fanout4536 (.A(net4538),
    .X(net4536));
 sg13g2_buf_8 fanout4537 (.A(net4538),
    .X(net4537));
 sg13g2_buf_8 fanout4538 (.A(_09614_),
    .X(net4538));
 sg13g2_buf_8 fanout4539 (.A(net4543),
    .X(net4539));
 sg13g2_buf_8 fanout4540 (.A(net4543),
    .X(net4540));
 sg13g2_buf_8 fanout4541 (.A(net4543),
    .X(net4541));
 sg13g2_buf_8 fanout4542 (.A(net4543),
    .X(net4542));
 sg13g2_buf_8 fanout4543 (.A(_09613_),
    .X(net4543));
 sg13g2_buf_8 fanout4544 (.A(net4548),
    .X(net4544));
 sg13g2_buf_8 fanout4545 (.A(net4548),
    .X(net4545));
 sg13g2_buf_8 fanout4546 (.A(net4547),
    .X(net4546));
 sg13g2_buf_8 fanout4547 (.A(net4548),
    .X(net4547));
 sg13g2_buf_8 fanout4548 (.A(_09612_),
    .X(net4548));
 sg13g2_buf_8 fanout4549 (.A(net4553),
    .X(net4549));
 sg13g2_buf_8 fanout4550 (.A(net4553),
    .X(net4550));
 sg13g2_buf_8 fanout4551 (.A(net4553),
    .X(net4551));
 sg13g2_buf_8 fanout4552 (.A(net4553),
    .X(net4552));
 sg13g2_buf_8 fanout4553 (.A(_09611_),
    .X(net4553));
 sg13g2_buf_8 fanout4554 (.A(net4558),
    .X(net4554));
 sg13g2_buf_8 fanout4555 (.A(net4558),
    .X(net4555));
 sg13g2_buf_8 fanout4556 (.A(net4558),
    .X(net4556));
 sg13g2_buf_8 fanout4557 (.A(net4558),
    .X(net4557));
 sg13g2_buf_8 fanout4558 (.A(_09610_),
    .X(net4558));
 sg13g2_buf_8 fanout4559 (.A(net4563),
    .X(net4559));
 sg13g2_buf_8 fanout4560 (.A(net4563),
    .X(net4560));
 sg13g2_buf_8 fanout4561 (.A(net4563),
    .X(net4561));
 sg13g2_buf_8 fanout4562 (.A(net4563),
    .X(net4562));
 sg13g2_buf_8 fanout4563 (.A(_09608_),
    .X(net4563));
 sg13g2_buf_8 fanout4564 (.A(net4568),
    .X(net4564));
 sg13g2_buf_8 fanout4565 (.A(net4568),
    .X(net4565));
 sg13g2_buf_8 fanout4566 (.A(net4567),
    .X(net4566));
 sg13g2_buf_8 fanout4567 (.A(net4568),
    .X(net4567));
 sg13g2_buf_8 fanout4568 (.A(_09607_),
    .X(net4568));
 sg13g2_buf_8 fanout4569 (.A(net4573),
    .X(net4569));
 sg13g2_buf_8 fanout4570 (.A(net4573),
    .X(net4570));
 sg13g2_buf_8 fanout4571 (.A(net4573),
    .X(net4571));
 sg13g2_buf_8 fanout4572 (.A(net4573),
    .X(net4572));
 sg13g2_buf_8 fanout4573 (.A(_09604_),
    .X(net4573));
 sg13g2_buf_8 fanout4574 (.A(net4578),
    .X(net4574));
 sg13g2_buf_8 fanout4575 (.A(net4578),
    .X(net4575));
 sg13g2_buf_8 fanout4576 (.A(net4577),
    .X(net4576));
 sg13g2_buf_8 fanout4577 (.A(net4578),
    .X(net4577));
 sg13g2_buf_8 fanout4578 (.A(_09602_),
    .X(net4578));
 sg13g2_buf_8 fanout4579 (.A(net4583),
    .X(net4579));
 sg13g2_buf_8 fanout4580 (.A(net4583),
    .X(net4580));
 sg13g2_buf_8 fanout4581 (.A(net4582),
    .X(net4581));
 sg13g2_buf_8 fanout4582 (.A(net4583),
    .X(net4582));
 sg13g2_buf_8 fanout4583 (.A(_09600_),
    .X(net4583));
 sg13g2_buf_8 fanout4584 (.A(net4588),
    .X(net4584));
 sg13g2_buf_8 fanout4585 (.A(net4588),
    .X(net4585));
 sg13g2_buf_8 fanout4586 (.A(net4588),
    .X(net4586));
 sg13g2_buf_8 fanout4587 (.A(net4588),
    .X(net4587));
 sg13g2_buf_8 fanout4588 (.A(_09599_),
    .X(net4588));
 sg13g2_buf_8 fanout4589 (.A(net4593),
    .X(net4589));
 sg13g2_buf_8 fanout4590 (.A(net4593),
    .X(net4590));
 sg13g2_buf_8 fanout4591 (.A(net4592),
    .X(net4591));
 sg13g2_buf_8 fanout4592 (.A(net4593),
    .X(net4592));
 sg13g2_buf_8 fanout4593 (.A(_09597_),
    .X(net4593));
 sg13g2_buf_8 fanout4594 (.A(_09277_),
    .X(net4594));
 sg13g2_buf_2 fanout4595 (.A(_09255_),
    .X(net4595));
 sg13g2_buf_8 fanout4596 (.A(_08991_),
    .X(net4596));
 sg13g2_buf_8 fanout4597 (.A(_08990_),
    .X(net4597));
 sg13g2_buf_8 fanout4598 (.A(_08820_),
    .X(net4598));
 sg13g2_buf_8 fanout4599 (.A(_08808_),
    .X(net4599));
 sg13g2_buf_1 fanout4600 (.A(_08808_),
    .X(net4600));
 sg13g2_buf_2 fanout4601 (.A(net4602),
    .X(net4601));
 sg13g2_buf_8 fanout4602 (.A(_08805_),
    .X(net4602));
 sg13g2_buf_8 fanout4603 (.A(net4604),
    .X(net4603));
 sg13g2_buf_8 fanout4604 (.A(net4608),
    .X(net4604));
 sg13g2_buf_8 fanout4605 (.A(net4606),
    .X(net4605));
 sg13g2_buf_8 fanout4606 (.A(net4607),
    .X(net4606));
 sg13g2_buf_8 fanout4607 (.A(net4608),
    .X(net4607));
 sg13g2_buf_8 fanout4608 (.A(net4611),
    .X(net4608));
 sg13g2_buf_8 fanout4609 (.A(net4610),
    .X(net4609));
 sg13g2_buf_8 fanout4610 (.A(net4611),
    .X(net4610));
 sg13g2_buf_8 fanout4611 (.A(_07604_),
    .X(net4611));
 sg13g2_buf_8 fanout4612 (.A(net4615),
    .X(net4612));
 sg13g2_buf_8 fanout4613 (.A(net4615),
    .X(net4613));
 sg13g2_buf_1 fanout4614 (.A(net4615),
    .X(net4614));
 sg13g2_buf_8 fanout4615 (.A(net4616),
    .X(net4615));
 sg13g2_buf_8 fanout4616 (.A(_07389_),
    .X(net4616));
 sg13g2_buf_8 fanout4617 (.A(net4623),
    .X(net4617));
 sg13g2_buf_8 fanout4618 (.A(net4623),
    .X(net4618));
 sg13g2_buf_8 fanout4619 (.A(net4620),
    .X(net4619));
 sg13g2_buf_8 fanout4620 (.A(net4621),
    .X(net4620));
 sg13g2_buf_8 fanout4621 (.A(net4622),
    .X(net4621));
 sg13g2_buf_2 fanout4622 (.A(net4623),
    .X(net4622));
 sg13g2_buf_8 fanout4623 (.A(_07388_),
    .X(net4623));
 sg13g2_buf_8 fanout4624 (.A(net4630),
    .X(net4624));
 sg13g2_buf_8 fanout4625 (.A(net4630),
    .X(net4625));
 sg13g2_buf_8 fanout4626 (.A(net4627),
    .X(net4626));
 sg13g2_buf_1 fanout4627 (.A(net4630),
    .X(net4627));
 sg13g2_buf_8 fanout4628 (.A(net4629),
    .X(net4628));
 sg13g2_buf_8 fanout4629 (.A(net4630),
    .X(net4629));
 sg13g2_buf_8 fanout4630 (.A(_07215_),
    .X(net4630));
 sg13g2_buf_8 fanout4631 (.A(net4635),
    .X(net4631));
 sg13g2_buf_8 fanout4632 (.A(net4635),
    .X(net4632));
 sg13g2_buf_8 fanout4633 (.A(net4635),
    .X(net4633));
 sg13g2_buf_8 fanout4634 (.A(net4635),
    .X(net4634));
 sg13g2_buf_8 fanout4635 (.A(_07214_),
    .X(net4635));
 sg13g2_buf_8 fanout4636 (.A(net4637),
    .X(net4636));
 sg13g2_buf_8 fanout4637 (.A(net4640),
    .X(net4637));
 sg13g2_buf_8 fanout4638 (.A(net4639),
    .X(net4638));
 sg13g2_buf_8 fanout4639 (.A(net4640),
    .X(net4639));
 sg13g2_buf_8 fanout4640 (.A(_07214_),
    .X(net4640));
 sg13g2_buf_8 fanout4641 (.A(net4644),
    .X(net4641));
 sg13g2_buf_8 fanout4642 (.A(net4644),
    .X(net4642));
 sg13g2_buf_8 fanout4643 (.A(net4644),
    .X(net4643));
 sg13g2_buf_8 fanout4644 (.A(_06522_),
    .X(net4644));
 sg13g2_buf_8 fanout4645 (.A(net4646),
    .X(net4645));
 sg13g2_buf_8 fanout4646 (.A(net4647),
    .X(net4646));
 sg13g2_buf_8 fanout4647 (.A(net4653),
    .X(net4647));
 sg13g2_buf_8 fanout4648 (.A(net4649),
    .X(net4648));
 sg13g2_buf_1 fanout4649 (.A(net4650),
    .X(net4649));
 sg13g2_buf_1 fanout4650 (.A(net4653),
    .X(net4650));
 sg13g2_buf_8 fanout4651 (.A(net4652),
    .X(net4651));
 sg13g2_buf_8 fanout4652 (.A(net4653),
    .X(net4652));
 sg13g2_buf_8 fanout4653 (.A(_06412_),
    .X(net4653));
 sg13g2_buf_8 fanout4654 (.A(_06292_),
    .X(net4654));
 sg13g2_buf_8 fanout4655 (.A(_06292_),
    .X(net4655));
 sg13g2_buf_8 fanout4656 (.A(_06291_),
    .X(net4656));
 sg13g2_buf_8 fanout4657 (.A(_06291_),
    .X(net4657));
 sg13g2_buf_8 fanout4658 (.A(_05333_),
    .X(net4658));
 sg13g2_buf_8 fanout4659 (.A(_02925_),
    .X(net4659));
 sg13g2_buf_8 fanout4660 (.A(net4663),
    .X(net4660));
 sg13g2_buf_8 fanout4661 (.A(net4662),
    .X(net4661));
 sg13g2_buf_8 fanout4662 (.A(net4663),
    .X(net4662));
 sg13g2_buf_8 fanout4663 (.A(_02613_),
    .X(net4663));
 sg13g2_buf_8 fanout4664 (.A(net4667),
    .X(net4664));
 sg13g2_buf_8 fanout4665 (.A(net4666),
    .X(net4665));
 sg13g2_buf_8 fanout4666 (.A(net4667),
    .X(net4666));
 sg13g2_buf_8 fanout4667 (.A(_09990_),
    .X(net4667));
 sg13g2_buf_8 fanout4668 (.A(net4674),
    .X(net4668));
 sg13g2_buf_8 fanout4669 (.A(net4674),
    .X(net4669));
 sg13g2_buf_8 fanout4670 (.A(net4674),
    .X(net4670));
 sg13g2_buf_8 fanout4671 (.A(net4674),
    .X(net4671));
 sg13g2_buf_8 fanout4672 (.A(net4674),
    .X(net4672));
 sg13g2_buf_8 fanout4673 (.A(net4674),
    .X(net4673));
 sg13g2_buf_8 fanout4674 (.A(_09989_),
    .X(net4674));
 sg13g2_buf_8 fanout4675 (.A(net4677),
    .X(net4675));
 sg13g2_buf_8 fanout4676 (.A(net4677),
    .X(net4676));
 sg13g2_buf_8 fanout4677 (.A(_09592_),
    .X(net4677));
 sg13g2_buf_8 fanout4678 (.A(net4680),
    .X(net4678));
 sg13g2_buf_8 fanout4679 (.A(net4680),
    .X(net4679));
 sg13g2_buf_8 fanout4680 (.A(_09592_),
    .X(net4680));
 sg13g2_buf_8 fanout4681 (.A(_09276_),
    .X(net4681));
 sg13g2_buf_8 fanout4682 (.A(net4683),
    .X(net4682));
 sg13g2_buf_8 fanout4683 (.A(_09273_),
    .X(net4683));
 sg13g2_buf_8 fanout4684 (.A(_09253_),
    .X(net4684));
 sg13g2_buf_1 fanout4685 (.A(_09253_),
    .X(net4685));
 sg13g2_buf_8 fanout4686 (.A(net4687),
    .X(net4686));
 sg13g2_buf_8 fanout4687 (.A(_09088_),
    .X(net4687));
 sg13g2_buf_8 fanout4688 (.A(net4689),
    .X(net4688));
 sg13g2_buf_8 fanout4689 (.A(net4690),
    .X(net4689));
 sg13g2_buf_8 fanout4690 (.A(_09088_),
    .X(net4690));
 sg13g2_buf_8 fanout4691 (.A(_08819_),
    .X(net4691));
 sg13g2_buf_8 fanout4692 (.A(net4693),
    .X(net4692));
 sg13g2_buf_8 fanout4693 (.A(_08818_),
    .X(net4693));
 sg13g2_buf_8 fanout4694 (.A(_08814_),
    .X(net4694));
 sg13g2_buf_1 fanout4695 (.A(_08814_),
    .X(net4695));
 sg13g2_buf_8 fanout4696 (.A(_08787_),
    .X(net4696));
 sg13g2_buf_2 fanout4697 (.A(_07825_),
    .X(net4697));
 sg13g2_buf_8 fanout4698 (.A(net4699),
    .X(net4698));
 sg13g2_buf_8 fanout4699 (.A(_07218_),
    .X(net4699));
 sg13g2_buf_8 fanout4700 (.A(_07218_),
    .X(net4700));
 sg13g2_buf_8 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_2 fanout4702 (.A(_06940_),
    .X(net4702));
 sg13g2_buf_8 fanout4703 (.A(net4706),
    .X(net4703));
 sg13g2_buf_8 fanout4704 (.A(net4705),
    .X(net4704));
 sg13g2_buf_8 fanout4705 (.A(net4706),
    .X(net4705));
 sg13g2_buf_8 fanout4706 (.A(_06749_),
    .X(net4706));
 sg13g2_buf_8 fanout4707 (.A(_06738_),
    .X(net4707));
 sg13g2_buf_8 fanout4708 (.A(_06675_),
    .X(net4708));
 sg13g2_buf_2 fanout4709 (.A(_06675_),
    .X(net4709));
 sg13g2_buf_8 fanout4710 (.A(net4711),
    .X(net4710));
 sg13g2_buf_8 fanout4711 (.A(_06674_),
    .X(net4711));
 sg13g2_buf_2 fanout4712 (.A(_06659_),
    .X(net4712));
 sg13g2_buf_8 fanout4713 (.A(net4715),
    .X(net4713));
 sg13g2_buf_8 fanout4714 (.A(net4715),
    .X(net4714));
 sg13g2_buf_8 fanout4715 (.A(_06410_),
    .X(net4715));
 sg13g2_buf_8 fanout4716 (.A(net4717),
    .X(net4716));
 sg13g2_buf_2 fanout4717 (.A(_06052_),
    .X(net4717));
 sg13g2_buf_8 fanout4718 (.A(net4719),
    .X(net4718));
 sg13g2_buf_2 fanout4719 (.A(net4720),
    .X(net4719));
 sg13g2_buf_1 fanout4720 (.A(net4727),
    .X(net4720));
 sg13g2_buf_8 fanout4721 (.A(net4722),
    .X(net4721));
 sg13g2_buf_8 fanout4722 (.A(net4727),
    .X(net4722));
 sg13g2_buf_8 fanout4723 (.A(net4725),
    .X(net4723));
 sg13g2_buf_1 fanout4724 (.A(net4725),
    .X(net4724));
 sg13g2_buf_1 fanout4725 (.A(net4726),
    .X(net4725));
 sg13g2_buf_8 fanout4726 (.A(net4727),
    .X(net4726));
 sg13g2_buf_8 fanout4727 (.A(_05835_),
    .X(net4727));
 sg13g2_buf_8 fanout4728 (.A(net4729),
    .X(net4728));
 sg13g2_buf_8 fanout4729 (.A(net4731),
    .X(net4729));
 sg13g2_buf_8 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_8 fanout4731 (.A(net4732),
    .X(net4731));
 sg13g2_buf_8 fanout4732 (.A(net4734),
    .X(net4732));
 sg13g2_buf_8 fanout4733 (.A(net4734),
    .X(net4733));
 sg13g2_buf_2 fanout4734 (.A(_05833_),
    .X(net4734));
 sg13g2_buf_8 fanout4735 (.A(net4736),
    .X(net4735));
 sg13g2_buf_8 fanout4736 (.A(net4737),
    .X(net4736));
 sg13g2_buf_8 fanout4737 (.A(_05831_),
    .X(net4737));
 sg13g2_buf_8 fanout4738 (.A(net4739),
    .X(net4738));
 sg13g2_buf_8 fanout4739 (.A(net4740),
    .X(net4739));
 sg13g2_buf_8 fanout4740 (.A(_05487_),
    .X(net4740));
 sg13g2_buf_8 fanout4741 (.A(net4743),
    .X(net4741));
 sg13g2_buf_8 fanout4742 (.A(net4743),
    .X(net4742));
 sg13g2_buf_8 fanout4743 (.A(net4750),
    .X(net4743));
 sg13g2_buf_8 fanout4744 (.A(net4745),
    .X(net4744));
 sg13g2_buf_8 fanout4745 (.A(net4746),
    .X(net4745));
 sg13g2_buf_8 fanout4746 (.A(net4750),
    .X(net4746));
 sg13g2_buf_8 fanout4747 (.A(net4748),
    .X(net4747));
 sg13g2_buf_8 fanout4748 (.A(net4749),
    .X(net4748));
 sg13g2_buf_1 fanout4749 (.A(net4750),
    .X(net4749));
 sg13g2_buf_8 fanout4750 (.A(_05480_),
    .X(net4750));
 sg13g2_buf_8 fanout4751 (.A(_05480_),
    .X(net4751));
 sg13g2_buf_8 fanout4752 (.A(_05480_),
    .X(net4752));
 sg13g2_buf_8 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_8 fanout4754 (.A(_05416_),
    .X(net4754));
 sg13g2_buf_8 fanout4755 (.A(net4756),
    .X(net4755));
 sg13g2_buf_8 fanout4756 (.A(_05415_),
    .X(net4756));
 sg13g2_buf_8 fanout4757 (.A(_05415_),
    .X(net4757));
 sg13g2_buf_8 fanout4758 (.A(net2955),
    .X(net4758));
 sg13g2_buf_8 fanout4759 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ),
    .X(net4759));
 sg13g2_buf_8 fanout4760 (.A(net4761),
    .X(net4760));
 sg13g2_buf_8 fanout4761 (.A(net4762),
    .X(net4761));
 sg13g2_buf_8 fanout4762 (.A(net1584),
    .X(net4762));
 sg13g2_buf_8 fanout4763 (.A(net4764),
    .X(net4763));
 sg13g2_buf_8 fanout4764 (.A(net4766),
    .X(net4764));
 sg13g2_buf_8 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_8 fanout4766 (.A(net4769),
    .X(net4766));
 sg13g2_buf_8 fanout4767 (.A(net4768),
    .X(net4767));
 sg13g2_buf_8 fanout4768 (.A(net4769),
    .X(net4768));
 sg13g2_buf_8 fanout4769 (.A(net4774),
    .X(net4769));
 sg13g2_buf_8 fanout4770 (.A(net4774),
    .X(net4770));
 sg13g2_buf_1 fanout4771 (.A(net4774),
    .X(net4771));
 sg13g2_buf_8 fanout4772 (.A(net4773),
    .X(net4772));
 sg13g2_buf_1 fanout4773 (.A(net4774),
    .X(net4773));
 sg13g2_buf_8 fanout4774 (.A(net2825),
    .X(net4774));
 sg13g2_buf_8 fanout4775 (.A(net4776),
    .X(net4775));
 sg13g2_buf_8 fanout4776 (.A(net4777),
    .X(net4776));
 sg13g2_buf_8 fanout4777 (.A(net4781),
    .X(net4777));
 sg13g2_buf_8 fanout4778 (.A(net4780),
    .X(net4778));
 sg13g2_buf_8 fanout4779 (.A(net4780),
    .X(net4779));
 sg13g2_buf_8 fanout4780 (.A(net4781),
    .X(net4780));
 sg13g2_buf_8 fanout4781 (.A(\soc_inst.mem_ctrl.access_state[1] ),
    .X(net4781));
 sg13g2_buf_8 fanout4782 (.A(net2926),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(net2973),
    .X(net4783));
 sg13g2_buf_1 fanout4784 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ),
    .X(net4784));
 sg13g2_buf_8 fanout4785 (.A(net4786),
    .X(net4785));
 sg13g2_buf_8 fanout4786 (.A(net2939),
    .X(net4786));
 sg13g2_buf_8 fanout4787 (.A(net2971),
    .X(net4787));
 sg13g2_buf_8 fanout4788 (.A(net4789),
    .X(net4788));
 sg13g2_buf_8 fanout4789 (.A(net4794),
    .X(net4789));
 sg13g2_buf_8 fanout4790 (.A(net4791),
    .X(net4790));
 sg13g2_buf_8 fanout4791 (.A(net4794),
    .X(net4791));
 sg13g2_buf_8 fanout4792 (.A(net4793),
    .X(net4792));
 sg13g2_buf_8 fanout4793 (.A(net4794),
    .X(net4793));
 sg13g2_buf_8 fanout4794 (.A(\soc_inst.pwm_inst.channel_idx [0]),
    .X(net4794));
 sg13g2_buf_8 fanout4795 (.A(net4796),
    .X(net4795));
 sg13g2_buf_8 fanout4796 (.A(\soc_inst.core_mem_addr[3] ),
    .X(net4796));
 sg13g2_buf_8 fanout4797 (.A(net4799),
    .X(net4797));
 sg13g2_buf_8 fanout4798 (.A(net4799),
    .X(net4798));
 sg13g2_buf_8 fanout4799 (.A(\soc_inst.core_mem_addr[2] ),
    .X(net4799));
 sg13g2_buf_8 fanout4800 (.A(net4801),
    .X(net4800));
 sg13g2_buf_8 fanout4801 (.A(\soc_inst.core_mem_re ),
    .X(net4801));
 sg13g2_buf_8 fanout4802 (.A(net4803),
    .X(net4802));
 sg13g2_buf_8 fanout4803 (.A(net4805),
    .X(net4803));
 sg13g2_buf_8 fanout4804 (.A(net4805),
    .X(net4804));
 sg13g2_buf_8 fanout4805 (.A(net4807),
    .X(net4805));
 sg13g2_buf_8 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_8 fanout4807 (.A(net2857),
    .X(net4807));
 sg13g2_buf_8 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_8 fanout4809 (.A(net4810),
    .X(net4809));
 sg13g2_buf_8 fanout4810 (.A(net4816),
    .X(net4810));
 sg13g2_buf_8 fanout4811 (.A(net4813),
    .X(net4811));
 sg13g2_buf_8 fanout4812 (.A(net4813),
    .X(net4812));
 sg13g2_buf_8 fanout4813 (.A(net4816),
    .X(net4813));
 sg13g2_buf_8 fanout4814 (.A(net4815),
    .X(net4814));
 sg13g2_buf_8 fanout4815 (.A(net4816),
    .X(net4815));
 sg13g2_buf_8 fanout4816 (.A(\soc_inst.cpu_core.alu.b[3] ),
    .X(net4816));
 sg13g2_buf_8 fanout4817 (.A(net4818),
    .X(net4817));
 sg13g2_buf_8 fanout4818 (.A(net4819),
    .X(net4818));
 sg13g2_buf_2 fanout4819 (.A(net4820),
    .X(net4819));
 sg13g2_buf_8 fanout4820 (.A(net4822),
    .X(net4820));
 sg13g2_buf_8 fanout4821 (.A(net4822),
    .X(net4821));
 sg13g2_buf_8 fanout4822 (.A(net4823),
    .X(net4822));
 sg13g2_buf_8 fanout4823 (.A(net2938),
    .X(net4823));
 sg13g2_buf_8 fanout4824 (.A(net4825),
    .X(net4824));
 sg13g2_buf_1 fanout4825 (.A(net4826),
    .X(net4825));
 sg13g2_buf_1 fanout4826 (.A(net4828),
    .X(net4826));
 sg13g2_buf_8 fanout4827 (.A(net4828),
    .X(net4827));
 sg13g2_buf_2 fanout4828 (.A(net4832),
    .X(net4828));
 sg13g2_buf_8 fanout4829 (.A(net4832),
    .X(net4829));
 sg13g2_buf_8 fanout4830 (.A(net4832),
    .X(net4830));
 sg13g2_buf_8 fanout4831 (.A(net4832),
    .X(net4831));
 sg13g2_buf_8 fanout4832 (.A(\soc_inst.cpu_core.alu.b[1] ),
    .X(net4832));
 sg13g2_buf_8 fanout4833 (.A(net4834),
    .X(net4833));
 sg13g2_buf_1 fanout4834 (.A(net4838),
    .X(net4834));
 sg13g2_buf_8 fanout4835 (.A(net4836),
    .X(net4835));
 sg13g2_buf_8 fanout4836 (.A(net4837),
    .X(net4836));
 sg13g2_buf_8 fanout4837 (.A(net4838),
    .X(net4837));
 sg13g2_buf_2 fanout4838 (.A(net2965),
    .X(net4838));
 sg13g2_buf_8 fanout4839 (.A(net4840),
    .X(net4839));
 sg13g2_buf_8 fanout4840 (.A(net4844),
    .X(net4840));
 sg13g2_buf_8 fanout4841 (.A(net4844),
    .X(net4841));
 sg13g2_buf_8 fanout4842 (.A(net4844),
    .X(net4842));
 sg13g2_buf_1 fanout4843 (.A(net4844),
    .X(net4843));
 sg13g2_buf_8 fanout4844 (.A(net4847),
    .X(net4844));
 sg13g2_buf_8 fanout4845 (.A(net4846),
    .X(net4845));
 sg13g2_buf_8 fanout4846 (.A(net4847),
    .X(net4846));
 sg13g2_buf_8 fanout4847 (.A(\soc_inst.cpu_core.alu.b[0] ),
    .X(net4847));
 sg13g2_buf_8 fanout4848 (.A(net4851),
    .X(net4848));
 sg13g2_buf_8 fanout4849 (.A(net4851),
    .X(net4849));
 sg13g2_buf_8 fanout4850 (.A(net4851),
    .X(net4850));
 sg13g2_buf_8 fanout4851 (.A(net2975),
    .X(net4851));
 sg13g2_buf_8 fanout4852 (.A(\soc_inst.cpu_core.alu.b[0] ),
    .X(net4852));
 sg13g2_buf_8 fanout4853 (.A(net4854),
    .X(net4853));
 sg13g2_buf_8 fanout4854 (.A(\soc_inst.cpu_core.alu.a[31] ),
    .X(net4854));
 sg13g2_buf_8 fanout4855 (.A(net2957),
    .X(net4855));
 sg13g2_buf_8 fanout4856 (.A(\soc_inst.cpu_core.alu.a[26] ),
    .X(net4856));
 sg13g2_buf_1 fanout4857 (.A(\soc_inst.cpu_core.alu.a[26] ),
    .X(net4857));
 sg13g2_buf_8 fanout4858 (.A(\soc_inst.cpu_core.alu.a[25] ),
    .X(net4858));
 sg13g2_buf_8 fanout4859 (.A(\soc_inst.cpu_core.alu.a[23] ),
    .X(net4859));
 sg13g2_buf_8 fanout4860 (.A(net2961),
    .X(net4860));
 sg13g2_buf_8 fanout4861 (.A(net2967),
    .X(net4861));
 sg13g2_buf_8 fanout4862 (.A(net2930),
    .X(net4862));
 sg13g2_buf_8 fanout4863 (.A(net2966),
    .X(net4863));
 sg13g2_buf_8 fanout4864 (.A(net2875),
    .X(net4864));
 sg13g2_buf_8 fanout4865 (.A(net2747),
    .X(net4865));
 sg13g2_buf_8 fanout4866 (.A(\soc_inst.core_mem_flag[2] ),
    .X(net4866));
 sg13g2_buf_8 fanout4867 (.A(\soc_inst.core_mem_flag[2] ),
    .X(net4867));
 sg13g2_buf_8 fanout4868 (.A(net4870),
    .X(net4868));
 sg13g2_buf_8 fanout4869 (.A(net4870),
    .X(net4869));
 sg13g2_buf_8 fanout4870 (.A(\soc_inst.core_mem_flag[2] ),
    .X(net4870));
 sg13g2_buf_8 fanout4871 (.A(net4874),
    .X(net4871));
 sg13g2_buf_8 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_8 fanout4873 (.A(net4874),
    .X(net4873));
 sg13g2_buf_8 fanout4874 (.A(\soc_inst.core_mem_flag[1] ),
    .X(net4874));
 sg13g2_buf_8 fanout4875 (.A(\soc_inst.core_mem_flag[1] ),
    .X(net4875));
 sg13g2_buf_8 fanout4876 (.A(net4877),
    .X(net4876));
 sg13g2_buf_8 fanout4877 (.A(net2638),
    .X(net4877));
 sg13g2_buf_8 fanout4878 (.A(net2942),
    .X(net4878));
 sg13g2_buf_8 fanout4879 (.A(net2716),
    .X(net4879));
 sg13g2_buf_8 fanout4880 (.A(net4882),
    .X(net4880));
 sg13g2_buf_1 fanout4881 (.A(net4882),
    .X(net4881));
 sg13g2_buf_8 fanout4882 (.A(net1614),
    .X(net4882));
 sg13g2_buf_8 fanout4883 (.A(net4888),
    .X(net4883));
 sg13g2_buf_8 fanout4884 (.A(net4888),
    .X(net4884));
 sg13g2_buf_8 fanout4885 (.A(net4887),
    .X(net4885));
 sg13g2_buf_8 fanout4886 (.A(net4888),
    .X(net4886));
 sg13g2_buf_1 fanout4887 (.A(net4888),
    .X(net4887));
 sg13g2_buf_8 fanout4888 (.A(net4951),
    .X(net4888));
 sg13g2_buf_8 fanout4889 (.A(net4890),
    .X(net4889));
 sg13g2_buf_8 fanout4890 (.A(net4896),
    .X(net4890));
 sg13g2_buf_8 fanout4891 (.A(net4895),
    .X(net4891));
 sg13g2_buf_8 fanout4892 (.A(net4894),
    .X(net4892));
 sg13g2_buf_1 fanout4893 (.A(net4894),
    .X(net4893));
 sg13g2_buf_1 fanout4894 (.A(net4895),
    .X(net4894));
 sg13g2_buf_1 fanout4895 (.A(net4896),
    .X(net4895));
 sg13g2_buf_2 fanout4896 (.A(net4951),
    .X(net4896));
 sg13g2_buf_8 fanout4897 (.A(net4899),
    .X(net4897));
 sg13g2_buf_8 fanout4898 (.A(net4899),
    .X(net4898));
 sg13g2_buf_8 fanout4899 (.A(net4909),
    .X(net4899));
 sg13g2_buf_8 fanout4900 (.A(net4909),
    .X(net4900));
 sg13g2_buf_8 fanout4901 (.A(net4909),
    .X(net4901));
 sg13g2_buf_8 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(net4904),
    .X(net4903));
 sg13g2_buf_8 fanout4904 (.A(net4909),
    .X(net4904));
 sg13g2_buf_8 fanout4905 (.A(net4908),
    .X(net4905));
 sg13g2_buf_1 fanout4906 (.A(net4908),
    .X(net4906));
 sg13g2_buf_8 fanout4907 (.A(net4908),
    .X(net4907));
 sg13g2_buf_8 fanout4908 (.A(net4909),
    .X(net4908));
 sg13g2_buf_8 fanout4909 (.A(net4951),
    .X(net4909));
 sg13g2_buf_8 fanout4910 (.A(net4911),
    .X(net4910));
 sg13g2_buf_8 fanout4911 (.A(net4912),
    .X(net4911));
 sg13g2_buf_8 fanout4912 (.A(net4926),
    .X(net4912));
 sg13g2_buf_8 fanout4913 (.A(net4916),
    .X(net4913));
 sg13g2_buf_8 fanout4914 (.A(net4915),
    .X(net4914));
 sg13g2_buf_8 fanout4915 (.A(net4916),
    .X(net4915));
 sg13g2_buf_8 fanout4916 (.A(net4917),
    .X(net4916));
 sg13g2_buf_8 fanout4917 (.A(net4926),
    .X(net4917));
 sg13g2_buf_8 fanout4918 (.A(net4921),
    .X(net4918));
 sg13g2_buf_1 fanout4919 (.A(net4921),
    .X(net4919));
 sg13g2_buf_8 fanout4920 (.A(net4921),
    .X(net4920));
 sg13g2_buf_2 fanout4921 (.A(net4925),
    .X(net4921));
 sg13g2_buf_8 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_8 fanout4923 (.A(net4925),
    .X(net4923));
 sg13g2_buf_8 fanout4924 (.A(net4925),
    .X(net4924));
 sg13g2_buf_2 fanout4925 (.A(net4926),
    .X(net4925));
 sg13g2_buf_8 fanout4926 (.A(net4951),
    .X(net4926));
 sg13g2_buf_8 fanout4927 (.A(net4929),
    .X(net4927));
 sg13g2_buf_1 fanout4928 (.A(net4929),
    .X(net4928));
 sg13g2_buf_8 fanout4929 (.A(net4934),
    .X(net4929));
 sg13g2_buf_8 fanout4930 (.A(net4931),
    .X(net4930));
 sg13g2_buf_8 fanout4931 (.A(net4933),
    .X(net4931));
 sg13g2_buf_8 fanout4932 (.A(net4933),
    .X(net4932));
 sg13g2_buf_8 fanout4933 (.A(net4934),
    .X(net4933));
 sg13g2_buf_8 fanout4934 (.A(net4950),
    .X(net4934));
 sg13g2_buf_8 fanout4935 (.A(net4937),
    .X(net4935));
 sg13g2_buf_8 fanout4936 (.A(net4937),
    .X(net4936));
 sg13g2_buf_8 fanout4937 (.A(net4942),
    .X(net4937));
 sg13g2_buf_8 fanout4938 (.A(net4939),
    .X(net4938));
 sg13g2_buf_8 fanout4939 (.A(net4942),
    .X(net4939));
 sg13g2_buf_8 fanout4940 (.A(net4942),
    .X(net4940));
 sg13g2_buf_8 fanout4941 (.A(net4942),
    .X(net4941));
 sg13g2_buf_8 fanout4942 (.A(net4949),
    .X(net4942));
 sg13g2_buf_8 fanout4943 (.A(net4949),
    .X(net4943));
 sg13g2_buf_1 fanout4944 (.A(net4949),
    .X(net4944));
 sg13g2_buf_8 fanout4945 (.A(net4948),
    .X(net4945));
 sg13g2_buf_8 fanout4946 (.A(net4948),
    .X(net4946));
 sg13g2_buf_8 fanout4947 (.A(net4948),
    .X(net4947));
 sg13g2_buf_8 fanout4948 (.A(net4949),
    .X(net4948));
 sg13g2_buf_8 fanout4949 (.A(net4950),
    .X(net4949));
 sg13g2_buf_8 fanout4950 (.A(net1614),
    .X(net4950));
 sg13g2_buf_8 fanout4951 (.A(net1752),
    .X(net4951));
 sg13g2_buf_8 fanout4952 (.A(net4953),
    .X(net4952));
 sg13g2_buf_1 fanout4953 (.A(net4954),
    .X(net4953));
 sg13g2_buf_8 fanout4954 (.A(net4956),
    .X(net4954));
 sg13g2_buf_8 fanout4955 (.A(net4956),
    .X(net4955));
 sg13g2_buf_8 fanout4956 (.A(net4966),
    .X(net4956));
 sg13g2_buf_8 fanout4957 (.A(net4959),
    .X(net4957));
 sg13g2_buf_8 fanout4958 (.A(net4959),
    .X(net4958));
 sg13g2_buf_8 fanout4959 (.A(net4966),
    .X(net4959));
 sg13g2_buf_8 fanout4960 (.A(net4963),
    .X(net4960));
 sg13g2_buf_8 fanout4961 (.A(net4962),
    .X(net4961));
 sg13g2_buf_8 fanout4962 (.A(net4963),
    .X(net4962));
 sg13g2_buf_8 fanout4963 (.A(net4966),
    .X(net4963));
 sg13g2_buf_8 fanout4964 (.A(net4965),
    .X(net4964));
 sg13g2_buf_8 fanout4965 (.A(net4966),
    .X(net4965));
 sg13g2_buf_8 fanout4966 (.A(net4998),
    .X(net4966));
 sg13g2_buf_8 fanout4967 (.A(net4968),
    .X(net4967));
 sg13g2_buf_8 fanout4968 (.A(net4969),
    .X(net4968));
 sg13g2_buf_8 fanout4969 (.A(net4998),
    .X(net4969));
 sg13g2_buf_8 fanout4970 (.A(net4977),
    .X(net4970));
 sg13g2_buf_1 fanout4971 (.A(net4977),
    .X(net4971));
 sg13g2_buf_8 fanout4972 (.A(net4977),
    .X(net4972));
 sg13g2_buf_8 fanout4973 (.A(net4975),
    .X(net4973));
 sg13g2_buf_8 fanout4974 (.A(net4976),
    .X(net4974));
 sg13g2_buf_8 fanout4975 (.A(net4976),
    .X(net4975));
 sg13g2_buf_8 fanout4976 (.A(net4977),
    .X(net4976));
 sg13g2_buf_8 fanout4977 (.A(net4986),
    .X(net4977));
 sg13g2_buf_8 fanout4978 (.A(net4979),
    .X(net4978));
 sg13g2_buf_8 fanout4979 (.A(net4980),
    .X(net4979));
 sg13g2_buf_8 fanout4980 (.A(net4981),
    .X(net4980));
 sg13g2_buf_8 fanout4981 (.A(net4986),
    .X(net4981));
 sg13g2_buf_8 fanout4982 (.A(net4983),
    .X(net4982));
 sg13g2_buf_1 fanout4983 (.A(net4984),
    .X(net4983));
 sg13g2_buf_8 fanout4984 (.A(net4985),
    .X(net4984));
 sg13g2_buf_8 fanout4985 (.A(net4986),
    .X(net4985));
 sg13g2_buf_8 fanout4986 (.A(net4998),
    .X(net4986));
 sg13g2_buf_8 fanout4987 (.A(net4988),
    .X(net4987));
 sg13g2_buf_8 fanout4988 (.A(net4992),
    .X(net4988));
 sg13g2_buf_8 fanout4989 (.A(net4990),
    .X(net4989));
 sg13g2_buf_8 fanout4990 (.A(net4991),
    .X(net4990));
 sg13g2_buf_8 fanout4991 (.A(net4992),
    .X(net4991));
 sg13g2_buf_8 fanout4992 (.A(net4997),
    .X(net4992));
 sg13g2_buf_8 fanout4993 (.A(net4994),
    .X(net4993));
 sg13g2_buf_8 fanout4994 (.A(net4997),
    .X(net4994));
 sg13g2_buf_8 fanout4995 (.A(net4996),
    .X(net4995));
 sg13g2_buf_2 fanout4996 (.A(net4997),
    .X(net4996));
 sg13g2_buf_8 fanout4997 (.A(net4998),
    .X(net4997));
 sg13g2_buf_8 fanout4998 (.A(net1613),
    .X(net4998));
 sg13g2_buf_8 fanout4999 (.A(\soc_inst.cpu_core.if_imm12[3] ),
    .X(net4999));
 sg13g2_buf_2 fanout5000 (.A(net2956),
    .X(net5000));
 sg13g2_buf_8 fanout5001 (.A(\soc_inst.cpu_core.if_imm12[2] ),
    .X(net5001));
 sg13g2_buf_8 fanout5002 (.A(net2434),
    .X(net5002));
 sg13g2_buf_8 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_8 fanout5004 (.A(net2889),
    .X(net5004));
 sg13g2_buf_8 fanout5005 (.A(\soc_inst.cpu_core.if_imm12[0] ),
    .X(net5005));
 sg13g2_buf_2 fanout5006 (.A(net2676),
    .X(net5006));
 sg13g2_buf_8 fanout5007 (.A(\soc_inst.cpu_core.if_instr[18] ),
    .X(net5007));
 sg13g2_buf_8 fanout5008 (.A(net1239),
    .X(net5008));
 sg13g2_buf_8 fanout5009 (.A(\soc_inst.cpu_core.if_instr[16] ),
    .X(net5009));
 sg13g2_buf_8 fanout5010 (.A(net1126),
    .X(net5010));
 sg13g2_buf_8 fanout5011 (.A(net5012),
    .X(net5011));
 sg13g2_buf_8 fanout5012 (.A(net2977),
    .X(net5012));
 sg13g2_buf_8 fanout5013 (.A(net5015),
    .X(net5013));
 sg13g2_buf_1 fanout5014 (.A(net5015),
    .X(net5014));
 sg13g2_buf_8 fanout5015 (.A(net5016),
    .X(net5015));
 sg13g2_buf_8 fanout5016 (.A(net2974),
    .X(net5016));
 sg13g2_buf_8 fanout5017 (.A(net2170),
    .X(net5017));
 sg13g2_buf_8 fanout5018 (.A(net770),
    .X(net5018));
 sg13g2_buf_8 fanout5019 (.A(\soc_inst.core_mem_wdata[14] ),
    .X(net5019));
 sg13g2_buf_8 fanout5020 (.A(\soc_inst.core_mem_wdata[13] ),
    .X(net5020));
 sg13g2_buf_8 fanout5021 (.A(\soc_inst.core_mem_wdata[12] ),
    .X(net5021));
 sg13g2_buf_8 fanout5022 (.A(net1620),
    .X(net5022));
 sg13g2_buf_8 fanout5023 (.A(net2194),
    .X(net5023));
 sg13g2_buf_8 fanout5024 (.A(net5025),
    .X(net5024));
 sg13g2_buf_8 fanout5025 (.A(net1012),
    .X(net5025));
 sg13g2_buf_8 fanout5026 (.A(net5027),
    .X(net5026));
 sg13g2_buf_8 fanout5027 (.A(net1968),
    .X(net5027));
 sg13g2_buf_8 fanout5028 (.A(net5030),
    .X(net5028));
 sg13g2_buf_8 fanout5029 (.A(net5030),
    .X(net5029));
 sg13g2_buf_8 fanout5030 (.A(net1036),
    .X(net5030));
 sg13g2_buf_8 fanout5031 (.A(net5032),
    .X(net5031));
 sg13g2_buf_8 fanout5032 (.A(\soc_inst.core_mem_wdata[6] ),
    .X(net5032));
 sg13g2_buf_8 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_8 fanout5034 (.A(net1023),
    .X(net5034));
 sg13g2_buf_8 fanout5035 (.A(net5037),
    .X(net5035));
 sg13g2_buf_8 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_8 fanout5037 (.A(net957),
    .X(net5037));
 sg13g2_buf_8 fanout5038 (.A(net5040),
    .X(net5038));
 sg13g2_buf_8 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_8 fanout5040 (.A(\soc_inst.core_mem_wdata[3] ),
    .X(net5040));
 sg13g2_buf_8 fanout5041 (.A(net5043),
    .X(net5041));
 sg13g2_buf_8 fanout5042 (.A(net5043),
    .X(net5042));
 sg13g2_buf_8 fanout5043 (.A(\soc_inst.core_mem_wdata[2] ),
    .X(net5043));
 sg13g2_buf_8 fanout5044 (.A(net5046),
    .X(net5044));
 sg13g2_buf_8 fanout5045 (.A(net5046),
    .X(net5045));
 sg13g2_buf_8 fanout5046 (.A(\soc_inst.core_mem_wdata[1] ),
    .X(net5046));
 sg13g2_buf_8 fanout5047 (.A(net5048),
    .X(net5047));
 sg13g2_buf_8 fanout5048 (.A(net5049),
    .X(net5048));
 sg13g2_buf_8 fanout5049 (.A(net5050),
    .X(net5049));
 sg13g2_buf_8 fanout5050 (.A(net1202),
    .X(net5050));
 sg13g2_buf_8 fanout5051 (.A(net5058),
    .X(net5051));
 sg13g2_buf_8 fanout5052 (.A(net5053),
    .X(net5052));
 sg13g2_buf_8 fanout5053 (.A(net5058),
    .X(net5053));
 sg13g2_buf_8 fanout5054 (.A(net5056),
    .X(net5054));
 sg13g2_buf_8 fanout5055 (.A(net5056),
    .X(net5055));
 sg13g2_buf_8 fanout5056 (.A(net5057),
    .X(net5056));
 sg13g2_buf_8 fanout5057 (.A(net5058),
    .X(net5057));
 sg13g2_buf_8 fanout5058 (.A(net2258),
    .X(net5058));
 sg13g2_buf_8 fanout5059 (.A(net2948),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(net2809),
    .X(net5060));
 sg13g2_buf_8 fanout5061 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .X(net5061));
 sg13g2_buf_8 fanout5062 (.A(net5063),
    .X(net5062));
 sg13g2_buf_8 fanout5063 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .X(net5063));
 sg13g2_buf_8 fanout5064 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .X(net5064));
 sg13g2_buf_8 fanout5065 (.A(net2952),
    .X(net5065));
 sg13g2_buf_8 fanout5066 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .X(net5066));
 sg13g2_buf_8 fanout5067 (.A(net5068),
    .X(net5067));
 sg13g2_buf_2 fanout5068 (.A(net5069),
    .X(net5068));
 sg13g2_buf_2 fanout5069 (.A(net5070),
    .X(net5069));
 sg13g2_buf_8 fanout5070 (.A(net5071),
    .X(net5070));
 sg13g2_buf_8 fanout5071 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ),
    .X(net5071));
 sg13g2_buf_8 fanout5072 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ),
    .X(net5072));
 sg13g2_buf_8 fanout5073 (.A(net2203),
    .X(net5073));
 sg13g2_buf_8 fanout5074 (.A(net5075),
    .X(net5074));
 sg13g2_buf_1 fanout5075 (.A(net5076),
    .X(net5075));
 sg13g2_buf_8 fanout5076 (.A(net2509),
    .X(net5076));
 sg13g2_buf_8 fanout5077 (.A(net5078),
    .X(net5077));
 sg13g2_buf_8 fanout5078 (.A(net5079),
    .X(net5078));
 sg13g2_buf_8 fanout5079 (.A(net5080),
    .X(net5079));
 sg13g2_buf_8 fanout5080 (.A(\soc_inst.mem_ctrl.spi_mem_inst.write_mosi ),
    .X(net5080));
 sg13g2_buf_8 fanout5081 (.A(net2862),
    .X(net5081));
 sg13g2_buf_8 fanout5082 (.A(net2847),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(\soc_inst.core_instr_data[15] ),
    .X(net5083));
 sg13g2_buf_8 fanout5084 (.A(net5085),
    .X(net5084));
 sg13g2_buf_8 fanout5085 (.A(net2603),
    .X(net5085));
 sg13g2_buf_8 fanout5086 (.A(net5088),
    .X(net5086));
 sg13g2_buf_1 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_8 fanout5088 (.A(net2206),
    .X(net5088));
 sg13g2_buf_8 fanout5089 (.A(net5091),
    .X(net5089));
 sg13g2_buf_1 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_8 fanout5091 (.A(net2460),
    .X(net5091));
 sg13g2_buf_8 fanout5092 (.A(net5093),
    .X(net5092));
 sg13g2_buf_8 fanout5093 (.A(net5094),
    .X(net5093));
 sg13g2_buf_1 fanout5094 (.A(net2906),
    .X(net5094));
 sg13g2_buf_8 fanout5095 (.A(net2705),
    .X(net5095));
 sg13g2_buf_2 fanout5096 (.A(\soc_inst.core_instr_data[10] ),
    .X(net5096));
 sg13g2_buf_8 fanout5097 (.A(net947),
    .X(net5097));
 sg13g2_buf_1 fanout5098 (.A(\soc_inst.core_instr_data[9] ),
    .X(net5098));
 sg13g2_buf_8 fanout5099 (.A(net5101),
    .X(net5099));
 sg13g2_buf_1 fanout5100 (.A(net5101),
    .X(net5100));
 sg13g2_buf_1 fanout5101 (.A(net689),
    .X(net5101));
 sg13g2_buf_8 fanout5102 (.A(net5103),
    .X(net5102));
 sg13g2_buf_8 fanout5103 (.A(net1211),
    .X(net5103));
 sg13g2_buf_8 fanout5104 (.A(net2941),
    .X(net5104));
 sg13g2_buf_1 fanout5105 (.A(net2941),
    .X(net5105));
 sg13g2_buf_8 fanout5106 (.A(net2890),
    .X(net5106));
 sg13g2_buf_1 fanout5107 (.A(net2890),
    .X(net5107));
 sg13g2_buf_8 fanout5108 (.A(net5109),
    .X(net5108));
 sg13g2_buf_2 fanout5109 (.A(net2819),
    .X(net5109));
 sg13g2_buf_8 fanout5110 (.A(net2784),
    .X(net5110));
 sg13g2_buf_8 fanout5111 (.A(net5112),
    .X(net5111));
 sg13g2_buf_8 fanout5112 (.A(net2552),
    .X(net5112));
 sg13g2_buf_8 fanout5113 (.A(net543),
    .X(net5113));
 sg13g2_buf_8 fanout5114 (.A(net2499),
    .X(net5114));
 sg13g2_buf_2 fanout5115 (.A(\soc_inst.i2c_inst.state[3] ),
    .X(net5115));
 sg13g2_buf_1 fanout5116 (.A(net2936),
    .X(net5116));
 sg13g2_buf_8 fanout5117 (.A(net5119),
    .X(net5117));
 sg13g2_buf_1 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_2 fanout5119 (.A(net279),
    .X(net5119));
 sg13g2_buf_8 fanout5120 (.A(\soc_inst.i2c_inst.state[0] ),
    .X(net5120));
 sg13g2_buf_8 fanout5121 (.A(net5122),
    .X(net5121));
 sg13g2_buf_8 fanout5122 (.A(net5123),
    .X(net5122));
 sg13g2_buf_8 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_2 fanout5124 (.A(\soc_inst.mem_ctrl.spi_mem_inst.stop ),
    .X(net5124));
 sg13g2_buf_8 fanout5125 (.A(net5126),
    .X(net5125));
 sg13g2_buf_8 fanout5126 (.A(net2963),
    .X(net5126));
 sg13g2_buf_8 fanout5127 (.A(net2937),
    .X(net5127));
 sg13g2_buf_8 fanout5128 (.A(net2950),
    .X(net5128));
 sg13g2_buf_8 fanout5129 (.A(net5130),
    .X(net5129));
 sg13g2_buf_8 fanout5130 (.A(net5131),
    .X(net5130));
 sg13g2_buf_8 fanout5131 (.A(net5135),
    .X(net5131));
 sg13g2_buf_8 fanout5132 (.A(net5133),
    .X(net5132));
 sg13g2_buf_8 fanout5133 (.A(net5134),
    .X(net5133));
 sg13g2_buf_8 fanout5134 (.A(net5135),
    .X(net5134));
 sg13g2_buf_8 fanout5135 (.A(net5157),
    .X(net5135));
 sg13g2_buf_8 fanout5136 (.A(net5139),
    .X(net5136));
 sg13g2_buf_8 fanout5137 (.A(net5139),
    .X(net5137));
 sg13g2_buf_1 fanout5138 (.A(net5139),
    .X(net5138));
 sg13g2_buf_8 fanout5139 (.A(net5157),
    .X(net5139));
 sg13g2_buf_8 fanout5140 (.A(net5143),
    .X(net5140));
 sg13g2_buf_8 fanout5141 (.A(net5143),
    .X(net5141));
 sg13g2_buf_8 fanout5142 (.A(net5143),
    .X(net5142));
 sg13g2_buf_8 fanout5143 (.A(net5157),
    .X(net5143));
 sg13g2_buf_8 fanout5144 (.A(net5147),
    .X(net5144));
 sg13g2_buf_8 fanout5145 (.A(net5147),
    .X(net5145));
 sg13g2_buf_8 fanout5146 (.A(net5147),
    .X(net5146));
 sg13g2_buf_8 fanout5147 (.A(net5157),
    .X(net5147));
 sg13g2_buf_8 fanout5148 (.A(net5149),
    .X(net5148));
 sg13g2_buf_8 fanout5149 (.A(net5150),
    .X(net5149));
 sg13g2_buf_8 fanout5150 (.A(net5157),
    .X(net5150));
 sg13g2_buf_8 fanout5151 (.A(net5156),
    .X(net5151));
 sg13g2_buf_8 fanout5152 (.A(net5156),
    .X(net5152));
 sg13g2_buf_2 fanout5153 (.A(net5156),
    .X(net5153));
 sg13g2_buf_8 fanout5154 (.A(net5155),
    .X(net5154));
 sg13g2_buf_8 fanout5155 (.A(net5156),
    .X(net5155));
 sg13g2_buf_8 fanout5156 (.A(net5157),
    .X(net5156));
 sg13g2_buf_8 fanout5157 (.A(net5308),
    .X(net5157));
 sg13g2_buf_8 fanout5158 (.A(net5161),
    .X(net5158));
 sg13g2_buf_8 fanout5159 (.A(net5160),
    .X(net5159));
 sg13g2_buf_8 fanout5160 (.A(net5161),
    .X(net5160));
 sg13g2_buf_8 fanout5161 (.A(net5165),
    .X(net5161));
 sg13g2_buf_8 fanout5162 (.A(net5164),
    .X(net5162));
 sg13g2_buf_1 fanout5163 (.A(net5164),
    .X(net5163));
 sg13g2_buf_8 fanout5164 (.A(net5165),
    .X(net5164));
 sg13g2_buf_8 fanout5165 (.A(net5174),
    .X(net5165));
 sg13g2_buf_8 fanout5166 (.A(net5171),
    .X(net5166));
 sg13g2_buf_8 fanout5167 (.A(net5171),
    .X(net5167));
 sg13g2_buf_8 fanout5168 (.A(net5170),
    .X(net5168));
 sg13g2_buf_8 fanout5169 (.A(net5170),
    .X(net5169));
 sg13g2_buf_8 fanout5170 (.A(net5171),
    .X(net5170));
 sg13g2_buf_8 fanout5171 (.A(net5173),
    .X(net5171));
 sg13g2_buf_8 fanout5172 (.A(net5173),
    .X(net5172));
 sg13g2_buf_8 fanout5173 (.A(net5174),
    .X(net5173));
 sg13g2_buf_8 fanout5174 (.A(net5308),
    .X(net5174));
 sg13g2_buf_8 fanout5175 (.A(net5178),
    .X(net5175));
 sg13g2_buf_1 fanout5176 (.A(net5178),
    .X(net5176));
 sg13g2_buf_8 fanout5177 (.A(net5178),
    .X(net5177));
 sg13g2_buf_8 fanout5178 (.A(net5179),
    .X(net5178));
 sg13g2_buf_8 fanout5179 (.A(net5190),
    .X(net5179));
 sg13g2_buf_8 fanout5180 (.A(net5182),
    .X(net5180));
 sg13g2_buf_8 fanout5181 (.A(net5182),
    .X(net5181));
 sg13g2_buf_8 fanout5182 (.A(net5183),
    .X(net5182));
 sg13g2_buf_8 fanout5183 (.A(net5190),
    .X(net5183));
 sg13g2_buf_8 fanout5184 (.A(net5185),
    .X(net5184));
 sg13g2_buf_8 fanout5185 (.A(net5189),
    .X(net5185));
 sg13g2_buf_8 fanout5186 (.A(net5189),
    .X(net5186));
 sg13g2_buf_8 fanout5187 (.A(net5189),
    .X(net5187));
 sg13g2_buf_8 fanout5188 (.A(net5189),
    .X(net5188));
 sg13g2_buf_8 fanout5189 (.A(net5190),
    .X(net5189));
 sg13g2_buf_8 fanout5190 (.A(net5228),
    .X(net5190));
 sg13g2_buf_8 fanout5191 (.A(net5193),
    .X(net5191));
 sg13g2_buf_8 fanout5192 (.A(net5193),
    .X(net5192));
 sg13g2_buf_8 fanout5193 (.A(net5198),
    .X(net5193));
 sg13g2_buf_8 fanout5194 (.A(net5195),
    .X(net5194));
 sg13g2_buf_8 fanout5195 (.A(net5198),
    .X(net5195));
 sg13g2_buf_8 fanout5196 (.A(net5198),
    .X(net5196));
 sg13g2_buf_1 fanout5197 (.A(net5198),
    .X(net5197));
 sg13g2_buf_8 fanout5198 (.A(net5203),
    .X(net5198));
 sg13g2_buf_8 fanout5199 (.A(net5203),
    .X(net5199));
 sg13g2_buf_8 fanout5200 (.A(net5203),
    .X(net5200));
 sg13g2_buf_8 fanout5201 (.A(net5202),
    .X(net5201));
 sg13g2_buf_8 fanout5202 (.A(net5203),
    .X(net5202));
 sg13g2_buf_8 fanout5203 (.A(net5228),
    .X(net5203));
 sg13g2_buf_8 fanout5204 (.A(net5207),
    .X(net5204));
 sg13g2_buf_8 fanout5205 (.A(net5207),
    .X(net5205));
 sg13g2_buf_2 fanout5206 (.A(net5207),
    .X(net5206));
 sg13g2_buf_8 fanout5207 (.A(net5215),
    .X(net5207));
 sg13g2_buf_8 fanout5208 (.A(net5210),
    .X(net5208));
 sg13g2_buf_8 fanout5209 (.A(net5210),
    .X(net5209));
 sg13g2_buf_8 fanout5210 (.A(net5215),
    .X(net5210));
 sg13g2_buf_8 fanout5211 (.A(net5215),
    .X(net5211));
 sg13g2_buf_8 fanout5212 (.A(net5215),
    .X(net5212));
 sg13g2_buf_8 fanout5213 (.A(net5214),
    .X(net5213));
 sg13g2_buf_8 fanout5214 (.A(net5215),
    .X(net5214));
 sg13g2_buf_8 fanout5215 (.A(net5228),
    .X(net5215));
 sg13g2_buf_8 fanout5216 (.A(net5221),
    .X(net5216));
 sg13g2_buf_8 fanout5217 (.A(net5221),
    .X(net5217));
 sg13g2_buf_8 fanout5218 (.A(net5220),
    .X(net5218));
 sg13g2_buf_8 fanout5219 (.A(net5220),
    .X(net5219));
 sg13g2_buf_8 fanout5220 (.A(net5221),
    .X(net5220));
 sg13g2_buf_8 fanout5221 (.A(net5227),
    .X(net5221));
 sg13g2_buf_8 fanout5222 (.A(net5224),
    .X(net5222));
 sg13g2_buf_2 fanout5223 (.A(net5224),
    .X(net5223));
 sg13g2_buf_8 fanout5224 (.A(net5227),
    .X(net5224));
 sg13g2_buf_8 fanout5225 (.A(net5227),
    .X(net5225));
 sg13g2_buf_8 fanout5226 (.A(net5227),
    .X(net5226));
 sg13g2_buf_8 fanout5227 (.A(net5228),
    .X(net5227));
 sg13g2_buf_8 fanout5228 (.A(net5308),
    .X(net5228));
 sg13g2_buf_8 fanout5229 (.A(net5241),
    .X(net5229));
 sg13g2_buf_8 fanout5230 (.A(net5234),
    .X(net5230));
 sg13g2_buf_8 fanout5231 (.A(net5234),
    .X(net5231));
 sg13g2_buf_8 fanout5232 (.A(net5234),
    .X(net5232));
 sg13g2_buf_2 fanout5233 (.A(net5234),
    .X(net5233));
 sg13g2_buf_8 fanout5234 (.A(net5241),
    .X(net5234));
 sg13g2_buf_8 fanout5235 (.A(net5239),
    .X(net5235));
 sg13g2_buf_8 fanout5236 (.A(net5239),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(net5239),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(net5239),
    .X(net5238));
 sg13g2_buf_8 fanout5239 (.A(net5240),
    .X(net5239));
 sg13g2_buf_8 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_8 fanout5241 (.A(net5307),
    .X(net5241));
 sg13g2_buf_8 fanout5242 (.A(net5246),
    .X(net5242));
 sg13g2_buf_8 fanout5243 (.A(net5246),
    .X(net5243));
 sg13g2_buf_8 fanout5244 (.A(net5245),
    .X(net5244));
 sg13g2_buf_8 fanout5245 (.A(net5246),
    .X(net5245));
 sg13g2_buf_8 fanout5246 (.A(net5252),
    .X(net5246));
 sg13g2_buf_8 fanout5247 (.A(net5252),
    .X(net5247));
 sg13g2_buf_1 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(net5252),
    .X(net5249));
 sg13g2_buf_8 fanout5250 (.A(net5251),
    .X(net5250));
 sg13g2_buf_8 fanout5251 (.A(net5252),
    .X(net5251));
 sg13g2_buf_8 fanout5252 (.A(net5307),
    .X(net5252));
 sg13g2_buf_8 fanout5253 (.A(net5254),
    .X(net5253));
 sg13g2_buf_8 fanout5254 (.A(net5261),
    .X(net5254));
 sg13g2_buf_8 fanout5255 (.A(net5261),
    .X(net5255));
 sg13g2_buf_8 fanout5256 (.A(net5261),
    .X(net5256));
 sg13g2_buf_8 fanout5257 (.A(net5259),
    .X(net5257));
 sg13g2_buf_8 fanout5258 (.A(net5259),
    .X(net5258));
 sg13g2_buf_8 fanout5259 (.A(net5260),
    .X(net5259));
 sg13g2_buf_8 fanout5260 (.A(net5261),
    .X(net5260));
 sg13g2_buf_8 fanout5261 (.A(net5307),
    .X(net5261));
 sg13g2_buf_8 fanout5262 (.A(net5266),
    .X(net5262));
 sg13g2_buf_8 fanout5263 (.A(net5266),
    .X(net5263));
 sg13g2_buf_8 fanout5264 (.A(net5266),
    .X(net5264));
 sg13g2_buf_8 fanout5265 (.A(net5266),
    .X(net5265));
 sg13g2_buf_8 fanout5266 (.A(net5287),
    .X(net5266));
 sg13g2_buf_8 fanout5267 (.A(net5269),
    .X(net5267));
 sg13g2_buf_8 fanout5268 (.A(net5269),
    .X(net5268));
 sg13g2_buf_8 fanout5269 (.A(net5287),
    .X(net5269));
 sg13g2_buf_8 fanout5270 (.A(net5274),
    .X(net5270));
 sg13g2_buf_1 fanout5271 (.A(net5274),
    .X(net5271));
 sg13g2_buf_8 fanout5272 (.A(net5274),
    .X(net5272));
 sg13g2_buf_2 fanout5273 (.A(net5274),
    .X(net5273));
 sg13g2_buf_2 fanout5274 (.A(net5287),
    .X(net5274));
 sg13g2_buf_8 fanout5275 (.A(net5276),
    .X(net5275));
 sg13g2_buf_8 fanout5276 (.A(net5281),
    .X(net5276));
 sg13g2_buf_8 fanout5277 (.A(net5281),
    .X(net5277));
 sg13g2_buf_2 fanout5278 (.A(net5281),
    .X(net5278));
 sg13g2_buf_8 fanout5279 (.A(net5280),
    .X(net5279));
 sg13g2_buf_8 fanout5280 (.A(net5281),
    .X(net5280));
 sg13g2_buf_8 fanout5281 (.A(net5287),
    .X(net5281));
 sg13g2_buf_8 fanout5282 (.A(net5286),
    .X(net5282));
 sg13g2_buf_8 fanout5283 (.A(net5286),
    .X(net5283));
 sg13g2_buf_8 fanout5284 (.A(net5285),
    .X(net5284));
 sg13g2_buf_8 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_8 fanout5286 (.A(net5287),
    .X(net5286));
 sg13g2_buf_8 fanout5287 (.A(net5306),
    .X(net5287));
 sg13g2_buf_8 fanout5288 (.A(net5291),
    .X(net5288));
 sg13g2_buf_8 fanout5289 (.A(net5291),
    .X(net5289));
 sg13g2_buf_8 fanout5290 (.A(net5291),
    .X(net5290));
 sg13g2_buf_8 fanout5291 (.A(net5294),
    .X(net5291));
 sg13g2_buf_8 fanout5292 (.A(net5293),
    .X(net5292));
 sg13g2_buf_8 fanout5293 (.A(net5294),
    .X(net5293));
 sg13g2_buf_8 fanout5294 (.A(net5306),
    .X(net5294));
 sg13g2_buf_8 fanout5295 (.A(net5298),
    .X(net5295));
 sg13g2_buf_8 fanout5296 (.A(net5298),
    .X(net5296));
 sg13g2_buf_1 fanout5297 (.A(net5298),
    .X(net5297));
 sg13g2_buf_8 fanout5298 (.A(net5306),
    .X(net5298));
 sg13g2_buf_8 fanout5299 (.A(net5304),
    .X(net5299));
 sg13g2_buf_8 fanout5300 (.A(net5304),
    .X(net5300));
 sg13g2_buf_8 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_8 fanout5302 (.A(net5303),
    .X(net5302));
 sg13g2_buf_8 fanout5303 (.A(net5304),
    .X(net5303));
 sg13g2_buf_8 fanout5304 (.A(net5305),
    .X(net5304));
 sg13g2_buf_8 fanout5305 (.A(net5306),
    .X(net5305));
 sg13g2_buf_8 fanout5306 (.A(net5307),
    .X(net5306));
 sg13g2_buf_8 fanout5307 (.A(net5308),
    .X(net5307));
 sg13g2_buf_8 fanout5308 (.A(rst_n),
    .X(net5308));
 sg13g2_buf_8 fanout5309 (.A(net5311),
    .X(net5309));
 sg13g2_buf_8 fanout5310 (.A(net5311),
    .X(net5310));
 sg13g2_buf_8 fanout5311 (.A(net5314),
    .X(net5311));
 sg13g2_buf_8 fanout5312 (.A(net5314),
    .X(net5312));
 sg13g2_buf_8 fanout5313 (.A(net5314),
    .X(net5313));
 sg13g2_buf_8 fanout5314 (.A(net5321),
    .X(net5314));
 sg13g2_buf_8 fanout5315 (.A(net5318),
    .X(net5315));
 sg13g2_buf_1 fanout5316 (.A(net5318),
    .X(net5316));
 sg13g2_buf_8 fanout5317 (.A(net5318),
    .X(net5317));
 sg13g2_buf_8 fanout5318 (.A(net5321),
    .X(net5318));
 sg13g2_buf_8 fanout5319 (.A(net5321),
    .X(net5319));
 sg13g2_buf_8 fanout5320 (.A(net5321),
    .X(net5320));
 sg13g2_buf_8 fanout5321 (.A(net5400),
    .X(net5321));
 sg13g2_buf_8 fanout5322 (.A(net5324),
    .X(net5322));
 sg13g2_buf_8 fanout5323 (.A(net5333),
    .X(net5323));
 sg13g2_buf_2 fanout5324 (.A(net5333),
    .X(net5324));
 sg13g2_buf_8 fanout5325 (.A(net5327),
    .X(net5325));
 sg13g2_buf_8 fanout5326 (.A(net5327),
    .X(net5326));
 sg13g2_buf_8 fanout5327 (.A(net5333),
    .X(net5327));
 sg13g2_buf_8 fanout5328 (.A(net5332),
    .X(net5328));
 sg13g2_buf_2 fanout5329 (.A(net5332),
    .X(net5329));
 sg13g2_buf_8 fanout5330 (.A(net5332),
    .X(net5330));
 sg13g2_buf_8 fanout5331 (.A(net5332),
    .X(net5331));
 sg13g2_buf_8 fanout5332 (.A(net5333),
    .X(net5332));
 sg13g2_buf_8 fanout5333 (.A(net5400),
    .X(net5333));
 sg13g2_buf_8 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_8 fanout5335 (.A(net5337),
    .X(net5335));
 sg13g2_buf_8 fanout5336 (.A(net5337),
    .X(net5336));
 sg13g2_buf_8 fanout5337 (.A(net5354),
    .X(net5337));
 sg13g2_buf_8 fanout5338 (.A(net5340),
    .X(net5338));
 sg13g2_buf_8 fanout5339 (.A(net5340),
    .X(net5339));
 sg13g2_buf_8 fanout5340 (.A(net5354),
    .X(net5340));
 sg13g2_buf_8 fanout5341 (.A(net5343),
    .X(net5341));
 sg13g2_buf_8 fanout5342 (.A(net5343),
    .X(net5342));
 sg13g2_buf_8 fanout5343 (.A(net5354),
    .X(net5343));
 sg13g2_buf_8 fanout5344 (.A(net5346),
    .X(net5344));
 sg13g2_buf_8 fanout5345 (.A(net5346),
    .X(net5345));
 sg13g2_buf_8 fanout5346 (.A(net5354),
    .X(net5346));
 sg13g2_buf_8 fanout5347 (.A(net5354),
    .X(net5347));
 sg13g2_buf_8 fanout5348 (.A(net5350),
    .X(net5348));
 sg13g2_buf_1 fanout5349 (.A(net5350),
    .X(net5349));
 sg13g2_buf_8 fanout5350 (.A(net5353),
    .X(net5350));
 sg13g2_buf_8 fanout5351 (.A(net5353),
    .X(net5351));
 sg13g2_buf_8 fanout5352 (.A(net5353),
    .X(net5352));
 sg13g2_buf_8 fanout5353 (.A(net5354),
    .X(net5353));
 sg13g2_buf_8 fanout5354 (.A(net5400),
    .X(net5354));
 sg13g2_buf_8 fanout5355 (.A(net5365),
    .X(net5355));
 sg13g2_buf_1 fanout5356 (.A(net5365),
    .X(net5356));
 sg13g2_buf_8 fanout5357 (.A(net5359),
    .X(net5357));
 sg13g2_buf_8 fanout5358 (.A(net5359),
    .X(net5358));
 sg13g2_buf_8 fanout5359 (.A(net5365),
    .X(net5359));
 sg13g2_buf_8 fanout5360 (.A(net5361),
    .X(net5360));
 sg13g2_buf_8 fanout5361 (.A(net5365),
    .X(net5361));
 sg13g2_buf_8 fanout5362 (.A(net5363),
    .X(net5362));
 sg13g2_buf_8 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_8 fanout5364 (.A(net5365),
    .X(net5364));
 sg13g2_buf_8 fanout5365 (.A(net5399),
    .X(net5365));
 sg13g2_buf_8 fanout5366 (.A(net5368),
    .X(net5366));
 sg13g2_buf_8 fanout5367 (.A(net5368),
    .X(net5367));
 sg13g2_buf_8 fanout5368 (.A(net5377),
    .X(net5368));
 sg13g2_buf_8 fanout5369 (.A(net5371),
    .X(net5369));
 sg13g2_buf_8 fanout5370 (.A(net5371),
    .X(net5370));
 sg13g2_buf_8 fanout5371 (.A(net5377),
    .X(net5371));
 sg13g2_buf_8 fanout5372 (.A(net5377),
    .X(net5372));
 sg13g2_buf_2 fanout5373 (.A(net5377),
    .X(net5373));
 sg13g2_buf_8 fanout5374 (.A(net5376),
    .X(net5374));
 sg13g2_buf_8 fanout5375 (.A(net5376),
    .X(net5375));
 sg13g2_buf_8 fanout5376 (.A(net5377),
    .X(net5376));
 sg13g2_buf_8 fanout5377 (.A(net5399),
    .X(net5377));
 sg13g2_buf_8 fanout5378 (.A(net5379),
    .X(net5378));
 sg13g2_buf_8 fanout5379 (.A(net5381),
    .X(net5379));
 sg13g2_buf_8 fanout5380 (.A(net5381),
    .X(net5380));
 sg13g2_buf_8 fanout5381 (.A(net5399),
    .X(net5381));
 sg13g2_buf_8 fanout5382 (.A(net5383),
    .X(net5382));
 sg13g2_buf_8 fanout5383 (.A(net5386),
    .X(net5383));
 sg13g2_buf_8 fanout5384 (.A(net5385),
    .X(net5384));
 sg13g2_buf_8 fanout5385 (.A(net5386),
    .X(net5385));
 sg13g2_buf_8 fanout5386 (.A(net5399),
    .X(net5386));
 sg13g2_buf_8 fanout5387 (.A(net5398),
    .X(net5387));
 sg13g2_buf_1 fanout5388 (.A(net5398),
    .X(net5388));
 sg13g2_buf_8 fanout5389 (.A(net5391),
    .X(net5389));
 sg13g2_buf_8 fanout5390 (.A(net5391),
    .X(net5390));
 sg13g2_buf_8 fanout5391 (.A(net5398),
    .X(net5391));
 sg13g2_buf_8 fanout5392 (.A(net5393),
    .X(net5392));
 sg13g2_buf_8 fanout5393 (.A(net5397),
    .X(net5393));
 sg13g2_buf_8 fanout5394 (.A(net5396),
    .X(net5394));
 sg13g2_buf_8 fanout5395 (.A(net5397),
    .X(net5395));
 sg13g2_buf_8 fanout5396 (.A(net5397),
    .X(net5396));
 sg13g2_buf_8 fanout5397 (.A(net5398),
    .X(net5397));
 sg13g2_buf_8 fanout5398 (.A(net5399),
    .X(net5398));
 sg13g2_buf_8 fanout5399 (.A(net5400),
    .X(net5399));
 sg13g2_buf_8 fanout5400 (.A(net5487),
    .X(net5400));
 sg13g2_buf_8 fanout5401 (.A(net5402),
    .X(net5401));
 sg13g2_buf_8 fanout5402 (.A(net5403),
    .X(net5402));
 sg13g2_buf_8 fanout5403 (.A(net5406),
    .X(net5403));
 sg13g2_buf_8 fanout5404 (.A(net5405),
    .X(net5404));
 sg13g2_buf_8 fanout5405 (.A(net5406),
    .X(net5405));
 sg13g2_buf_8 fanout5406 (.A(net5424),
    .X(net5406));
 sg13g2_buf_8 fanout5407 (.A(net5409),
    .X(net5407));
 sg13g2_buf_8 fanout5408 (.A(net5409),
    .X(net5408));
 sg13g2_buf_8 fanout5409 (.A(net5424),
    .X(net5409));
 sg13g2_buf_8 fanout5410 (.A(net5412),
    .X(net5410));
 sg13g2_buf_8 fanout5411 (.A(net5412),
    .X(net5411));
 sg13g2_buf_8 fanout5412 (.A(net5424),
    .X(net5412));
 sg13g2_buf_8 fanout5413 (.A(net5417),
    .X(net5413));
 sg13g2_buf_8 fanout5414 (.A(net5417),
    .X(net5414));
 sg13g2_buf_8 fanout5415 (.A(net5416),
    .X(net5415));
 sg13g2_buf_8 fanout5416 (.A(net5417),
    .X(net5416));
 sg13g2_buf_8 fanout5417 (.A(net5424),
    .X(net5417));
 sg13g2_buf_8 fanout5418 (.A(net5423),
    .X(net5418));
 sg13g2_buf_8 fanout5419 (.A(net5423),
    .X(net5419));
 sg13g2_buf_8 fanout5420 (.A(net5423),
    .X(net5420));
 sg13g2_buf_1 fanout5421 (.A(net5422),
    .X(net5421));
 sg13g2_buf_8 fanout5422 (.A(net5423),
    .X(net5422));
 sg13g2_buf_8 fanout5423 (.A(net5424),
    .X(net5423));
 sg13g2_buf_8 fanout5424 (.A(net5487),
    .X(net5424));
 sg13g2_buf_8 fanout5425 (.A(net5426),
    .X(net5425));
 sg13g2_buf_8 fanout5426 (.A(net5429),
    .X(net5426));
 sg13g2_buf_8 fanout5427 (.A(net5429),
    .X(net5427));
 sg13g2_buf_2 fanout5428 (.A(net5429),
    .X(net5428));
 sg13g2_buf_8 fanout5429 (.A(net5438),
    .X(net5429));
 sg13g2_buf_8 fanout5430 (.A(net5431),
    .X(net5430));
 sg13g2_buf_8 fanout5431 (.A(net5438),
    .X(net5431));
 sg13g2_buf_8 fanout5432 (.A(net5434),
    .X(net5432));
 sg13g2_buf_2 fanout5433 (.A(net5434),
    .X(net5433));
 sg13g2_buf_8 fanout5434 (.A(net5435),
    .X(net5434));
 sg13g2_buf_8 fanout5435 (.A(net5438),
    .X(net5435));
 sg13g2_buf_8 fanout5436 (.A(net5437),
    .X(net5436));
 sg13g2_buf_8 fanout5437 (.A(net5438),
    .X(net5437));
 sg13g2_buf_8 fanout5438 (.A(net5487),
    .X(net5438));
 sg13g2_buf_8 fanout5439 (.A(net5444),
    .X(net5439));
 sg13g2_buf_8 fanout5440 (.A(net5441),
    .X(net5440));
 sg13g2_buf_8 fanout5441 (.A(net5444),
    .X(net5441));
 sg13g2_buf_8 fanout5442 (.A(net5444),
    .X(net5442));
 sg13g2_buf_1 fanout5443 (.A(net5444),
    .X(net5443));
 sg13g2_buf_8 fanout5444 (.A(net5486),
    .X(net5444));
 sg13g2_buf_8 fanout5445 (.A(net5448),
    .X(net5445));
 sg13g2_buf_8 fanout5446 (.A(net5447),
    .X(net5446));
 sg13g2_buf_8 fanout5447 (.A(net5448),
    .X(net5447));
 sg13g2_buf_8 fanout5448 (.A(net5486),
    .X(net5448));
 sg13g2_buf_8 fanout5449 (.A(net5451),
    .X(net5449));
 sg13g2_buf_8 fanout5450 (.A(net5463),
    .X(net5450));
 sg13g2_buf_8 fanout5451 (.A(net5463),
    .X(net5451));
 sg13g2_buf_8 fanout5452 (.A(net5455),
    .X(net5452));
 sg13g2_buf_1 fanout5453 (.A(net5455),
    .X(net5453));
 sg13g2_buf_8 fanout5454 (.A(net5455),
    .X(net5454));
 sg13g2_buf_8 fanout5455 (.A(net5463),
    .X(net5455));
 sg13g2_buf_8 fanout5456 (.A(net5457),
    .X(net5456));
 sg13g2_buf_8 fanout5457 (.A(net5462),
    .X(net5457));
 sg13g2_buf_8 fanout5458 (.A(net5459),
    .X(net5458));
 sg13g2_buf_8 fanout5459 (.A(net5462),
    .X(net5459));
 sg13g2_buf_8 fanout5460 (.A(net5461),
    .X(net5460));
 sg13g2_buf_8 fanout5461 (.A(net5462),
    .X(net5461));
 sg13g2_buf_8 fanout5462 (.A(net5463),
    .X(net5462));
 sg13g2_buf_8 fanout5463 (.A(net5486),
    .X(net5463));
 sg13g2_buf_8 fanout5464 (.A(net5465),
    .X(net5464));
 sg13g2_buf_8 fanout5465 (.A(net5485),
    .X(net5465));
 sg13g2_buf_8 fanout5466 (.A(net5467),
    .X(net5466));
 sg13g2_buf_8 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_8 fanout5468 (.A(net5485),
    .X(net5468));
 sg13g2_buf_8 fanout5469 (.A(net5470),
    .X(net5469));
 sg13g2_buf_8 fanout5470 (.A(net5473),
    .X(net5470));
 sg13g2_buf_8 fanout5471 (.A(net5472),
    .X(net5471));
 sg13g2_buf_8 fanout5472 (.A(net5473),
    .X(net5472));
 sg13g2_buf_8 fanout5473 (.A(net5485),
    .X(net5473));
 sg13g2_buf_8 fanout5474 (.A(net5475),
    .X(net5474));
 sg13g2_buf_8 fanout5475 (.A(net5479),
    .X(net5475));
 sg13g2_buf_8 fanout5476 (.A(net5479),
    .X(net5476));
 sg13g2_buf_8 fanout5477 (.A(net5478),
    .X(net5477));
 sg13g2_buf_2 fanout5478 (.A(net5479),
    .X(net5478));
 sg13g2_buf_8 fanout5479 (.A(net5484),
    .X(net5479));
 sg13g2_buf_8 fanout5480 (.A(net5484),
    .X(net5480));
 sg13g2_buf_1 fanout5481 (.A(net5484),
    .X(net5481));
 sg13g2_buf_8 fanout5482 (.A(net5483),
    .X(net5482));
 sg13g2_buf_8 fanout5483 (.A(net5484),
    .X(net5483));
 sg13g2_buf_8 fanout5484 (.A(net5485),
    .X(net5484));
 sg13g2_buf_8 fanout5485 (.A(net5486),
    .X(net5485));
 sg13g2_buf_8 fanout5486 (.A(net5487),
    .X(net5486));
 sg13g2_buf_8 fanout5487 (.A(rst_n),
    .X(net5487));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tiehi _22451__14 (.L_HI(net14));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_8 clkbuf_6_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0_0_clk));
 sg13g2_buf_8 clkbuf_6_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1_0_clk));
 sg13g2_buf_8 clkbuf_6_2_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2_0_clk));
 sg13g2_buf_8 clkbuf_6_3_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3_0_clk));
 sg13g2_buf_8 clkbuf_6_4_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4_0_clk));
 sg13g2_buf_8 clkbuf_6_5_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5_0_clk));
 sg13g2_buf_8 clkbuf_6_6_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6_0_clk));
 sg13g2_buf_8 clkbuf_6_7_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7_0_clk));
 sg13g2_buf_8 clkbuf_6_8_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8_0_clk));
 sg13g2_buf_8 clkbuf_6_9_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9_0_clk));
 sg13g2_buf_8 clkbuf_6_10_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10_0_clk));
 sg13g2_buf_8 clkbuf_6_11_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11_0_clk));
 sg13g2_buf_8 clkbuf_6_12_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12_0_clk));
 sg13g2_buf_8 clkbuf_6_13_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13_0_clk));
 sg13g2_buf_8 clkbuf_6_14_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14_0_clk));
 sg13g2_buf_8 clkbuf_6_15_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15_0_clk));
 sg13g2_buf_8 clkbuf_6_16_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16_0_clk));
 sg13g2_buf_8 clkbuf_6_17_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17_0_clk));
 sg13g2_buf_8 clkbuf_6_18_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18_0_clk));
 sg13g2_buf_8 clkbuf_6_19_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19_0_clk));
 sg13g2_buf_8 clkbuf_6_20_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20_0_clk));
 sg13g2_buf_8 clkbuf_6_21_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21_0_clk));
 sg13g2_buf_8 clkbuf_6_22_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22_0_clk));
 sg13g2_buf_8 clkbuf_6_23_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23_0_clk));
 sg13g2_buf_8 clkbuf_6_24_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24_0_clk));
 sg13g2_buf_8 clkbuf_6_25_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25_0_clk));
 sg13g2_buf_8 clkbuf_6_26_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26_0_clk));
 sg13g2_buf_8 clkbuf_6_27_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27_0_clk));
 sg13g2_buf_8 clkbuf_6_28_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28_0_clk));
 sg13g2_buf_8 clkbuf_6_29_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29_0_clk));
 sg13g2_buf_8 clkbuf_6_30_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30_0_clk));
 sg13g2_buf_8 clkbuf_6_31_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31_0_clk));
 sg13g2_buf_8 clkbuf_6_32_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32_0_clk));
 sg13g2_buf_8 clkbuf_6_33_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33_0_clk));
 sg13g2_buf_8 clkbuf_6_34_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34_0_clk));
 sg13g2_buf_8 clkbuf_6_35_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35_0_clk));
 sg13g2_buf_8 clkbuf_6_36_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36_0_clk));
 sg13g2_buf_8 clkbuf_6_37_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37_0_clk));
 sg13g2_buf_8 clkbuf_6_38_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38_0_clk));
 sg13g2_buf_8 clkbuf_6_39_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39_0_clk));
 sg13g2_buf_8 clkbuf_6_40_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40_0_clk));
 sg13g2_buf_8 clkbuf_6_41_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41_0_clk));
 sg13g2_buf_8 clkbuf_6_42_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42_0_clk));
 sg13g2_buf_8 clkbuf_6_43_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43_0_clk));
 sg13g2_buf_8 clkbuf_6_44_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44_0_clk));
 sg13g2_buf_8 clkbuf_6_45_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45_0_clk));
 sg13g2_buf_8 clkbuf_6_46_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46_0_clk));
 sg13g2_buf_8 clkbuf_6_47_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47_0_clk));
 sg13g2_buf_8 clkbuf_6_48_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48_0_clk));
 sg13g2_buf_8 clkbuf_6_49_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49_0_clk));
 sg13g2_buf_8 clkbuf_6_50_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50_0_clk));
 sg13g2_buf_8 clkbuf_6_51_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51_0_clk));
 sg13g2_buf_8 clkbuf_6_52_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52_0_clk));
 sg13g2_buf_8 clkbuf_6_53_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53_0_clk));
 sg13g2_buf_8 clkbuf_6_54_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54_0_clk));
 sg13g2_buf_8 clkbuf_6_55_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55_0_clk));
 sg13g2_buf_8 clkbuf_6_56_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56_0_clk));
 sg13g2_buf_8 clkbuf_6_57_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57_0_clk));
 sg13g2_buf_8 clkbuf_6_58_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58_0_clk));
 sg13g2_buf_8 clkbuf_6_59_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59_0_clk));
 sg13g2_buf_8 clkbuf_6_60_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60_0_clk));
 sg13g2_buf_8 clkbuf_6_61_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61_0_clk));
 sg13g2_buf_8 clkbuf_6_62_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62_0_clk));
 sg13g2_buf_8 clkbuf_6_63_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_1_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_2_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_3_0_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_4_0_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_5_0_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_6_0_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_7_0_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_17_0_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_18_0_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_19_0_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_20_0_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_21_0_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_6_22_0_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_6_23_0_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_6_33_0_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_6_34_0_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_6_35_0_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_6_36_0_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_6_37_0_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_6_38_0_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_6_39_0_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_6_49_0_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_6_50_0_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_6_51_0_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_6_52_0_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_6_53_0_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_6_54_0_clk));
 sg13g2_buf_8 clkload27 (.A(clknet_6_55_0_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_leaf_259_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_250_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_251_clk));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_90_clk));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_85_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\soc_inst.cpu_core.csr_file.external_interrupt ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold2 (.A(\soc_inst.gpio_inst.gpio_sync1[6] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold3 (.A(\soc_inst.i2c_inst.transfer_done ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold4 (.A(\soc_inst.gpio_inst.gpio_sync1[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold5 (.A(\soc_inst.gpio_inst.gpio_sync1[4] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold6 (.A(\soc_inst.gpio_inst.gpio_sync1[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold7 (.A(\soc_inst.cpu_core.csr_file.timer_interrupt ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold8 (.A(\soc_inst.gpio_inst.gpio_sync1[3] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold9 (.A(\soc_inst.gpio_inst.gpio_sync1[0] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold10 (.A(\soc_inst.gpio_inst.gpio_sync1[5] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold11 (.A(\soc_inst.i2c_inst.arb_lost ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold12 (.A(\soc_inst.i2c_inst.ack_received ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold13 (.A(\soc_inst.mem_ctrl.spi_mem_inst.ram_in_quad_mode ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00002_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold15 (.A(\soc_inst.cpu_core.csr_file.mcause[15] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold16 (.A(\soc_inst.cpu_core.csr_file.mcause[8] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold17 (.A(\soc_inst.cpu_core.csr_file.mcause[11] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold18 (.A(\soc_inst.cpu_core.csr_file.mcause[22] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold19 (.A(\soc_inst.bus_spi_sclk ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold20 (.A(_00090_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold21 (.A(\soc_inst.cpu_core.csr_file.mcause[9] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold22 (.A(\soc_inst.cpu_core.csr_file.mcause[26] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold23 (.A(\soc_inst.cpu_core.csr_file.mcause[10] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold24 (.A(\soc_inst.cpu_core.csr_file.mcause[18] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold25 (.A(\soc_inst.cpu_core.csr_file.mcause[21] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold26 (.A(_00040_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold27 (.A(\soc_inst.cpu_core.csr_file.mcause[7] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold28 (.A(\soc_inst.mem_ctrl.next_instr_data[4] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold29 (.A(_00662_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold30 (.A(\soc_inst.mem_ctrl.next_instr_data[3] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold31 (.A(_00661_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold32 (.A(\soc_inst.cpu_core.csr_file.mcause[27] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold33 (.A(\soc_inst.cpu_core.csr_file.mscratch[7] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold34 (.A(_08475_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold35 (.A(\soc_inst.spi_inst.tx_shift_reg[19] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00146_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold37 (.A(\soc_inst.mem_ctrl.next_instr_data[18] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold38 (.A(_00676_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold39 (.A(\soc_inst.cpu_core.csr_file.mcause[5] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold40 (.A(\soc_inst.spi_inst.tx_shift_reg[15] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold41 (.A(_00141_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold42 (.A(\soc_inst.cpu_core.csr_file.mcause[23] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold43 (.A(_00042_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold44 (.A(\soc_inst.mem_ctrl.next_instr_data[21] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold45 (.A(_00679_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold46 (.A(\soc_inst.mem_ctrl.next_instr_data[5] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold47 (.A(_00663_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold48 (.A(\soc_inst.mem_ctrl.next_instr_data[19] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold49 (.A(_00677_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold50 (.A(\soc_inst.cpu_core.csr_file.mcause[24] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold51 (.A(\soc_inst.cpu_core.csr_file.mscratch[21] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold52 (.A(_08526_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold53 (.A(_00744_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold54 (.A(\soc_inst.cpu_core.csr_file.mscratch[15] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold55 (.A(_08502_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold56 (.A(_00738_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold57 (.A(\soc_inst.cpu_core.csr_file.mscratch[8] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold58 (.A(_08478_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold59 (.A(\soc_inst.spi_inst.tx_shift_reg[20] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00147_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold61 (.A(\soc_inst.mem_ctrl.next_instr_data[8] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00666_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold63 (.A(\soc_inst.cpu_core.csr_file.mscratch[10] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold64 (.A(_08482_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00733_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold66 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[11] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold67 (.A(_00844_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold68 (.A(\soc_inst.mem_ctrl.next_instr_data[24] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold69 (.A(_00682_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold70 (.A(\soc_inst.pwm_inst.channel_counter[1][0] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold71 (.A(\soc_inst.spi_inst.tx_shift_reg[11] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold72 (.A(_00137_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold73 (.A(\soc_inst.cpu_core.csr_file.mscratch[23] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold74 (.A(_08534_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00746_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold76 (.A(\soc_inst.cpu_core.csr_file.mscratch[9] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold77 (.A(_08480_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold78 (.A(_00732_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold79 (.A(\soc_inst.cpu_core.csr_file.mcause[29] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold80 (.A(_00228_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold81 (.A(_07132_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold82 (.A(_00404_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold83 (.A(\soc_inst.mem_ctrl.next_instr_data[17] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold84 (.A(_00675_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold85 (.A(\soc_inst.cpu_core.csr_file.mscratch[6] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold86 (.A(_08471_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold87 (.A(\soc_inst.spi_inst.tx_shift_reg[18] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold88 (.A(_00144_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold89 (.A(\soc_inst.cpu_core.csr_file.mscratch[5] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold90 (.A(_08467_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold91 (.A(\soc_inst.cpu_core.csr_file.mcause[6] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold92 (.A(\soc_inst.spi_inst.tx_shift_reg[6] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold93 (.A(_00163_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold94 (.A(\soc_inst.cpu_core.csr_file.mscratch[19] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold95 (.A(_08518_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00742_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold97 (.A(\soc_inst.cpu_core.csr_file.mscratch[14] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold98 (.A(_08498_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold99 (.A(_00737_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold100 (.A(\soc_inst.cpu_core.csr_file.mcause[14] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold101 (.A(\soc_inst.mem_ctrl.next_instr_data[10] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold102 (.A(_00668_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold103 (.A(\soc_inst.cpu_core.csr_file.mcause[25] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold104 (.A(\soc_inst.mem_ctrl.next_instr_data[6] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold105 (.A(_00664_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold106 (.A(\soc_inst.mem_ctrl.next_instr_data[23] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold107 (.A(_00681_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold108 (.A(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold109 (.A(\soc_inst.spi_inst.tx_shift_reg[16] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold110 (.A(_00142_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold111 (.A(\soc_inst.mem_ctrl.next_instr_data[30] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold112 (.A(_00688_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold113 (.A(\soc_inst.core_instr_data[23] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00614_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold115 (.A(\soc_inst.cpu_core.csr_file.mscratch[18] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold116 (.A(_08514_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00741_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold118 (.A(\soc_inst.cpu_core.mem_instr[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold119 (.A(_01071_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold120 (.A(\soc_inst.core_instr_data[16] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold121 (.A(_00607_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold122 (.A(\soc_inst.mem_ctrl.next_instr_data[11] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold123 (.A(_00669_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold124 (.A(\soc_inst.mem_ctrl.next_instr_data[2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold125 (.A(_00660_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold126 (.A(\soc_inst.mem_ctrl.next_instr_data[16] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold127 (.A(_00674_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold128 (.A(\soc_inst.cpu_core.csr_file.mscratch[16] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold129 (.A(_08506_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold130 (.A(_00739_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold131 (.A(\soc_inst.cpu_core.csr_file.mscratch[12] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold132 (.A(_08490_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold133 (.A(\soc_inst.mem_ctrl.next_instr_data[1] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold134 (.A(_00659_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold135 (.A(\soc_inst.mem_ctrl.spi_data_in[27] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold136 (.A(_00548_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold137 (.A(\soc_inst.spi_inst.tx_shift_reg[10] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold138 (.A(_00136_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold139 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[4] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold140 (.A(_00837_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold141 (.A(\soc_inst.cpu_core.csr_file.mscratch[13] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold142 (.A(_08494_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold143 (.A(_00736_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold144 (.A(\soc_inst.mem_ctrl.next_instr_data[27] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold145 (.A(_00685_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold146 (.A(\soc_inst.spi_inst.tx_shift_reg[0] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold147 (.A(_00145_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold148 (.A(\soc_inst.mem_ctrl.spi_data_in[29] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold149 (.A(_00550_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold150 (.A(\soc_inst.mem_ctrl.next_instr_data[12] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold151 (.A(_00670_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold152 (.A(\soc_inst.mem_ctrl.next_instr_data[26] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold153 (.A(_00684_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold154 (.A(\soc_inst.spi_inst.tx_shift_reg[26] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold155 (.A(_00153_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold156 (.A(\soc_inst.mem_ctrl.next_instr_data[13] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold157 (.A(_00671_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold158 (.A(\soc_inst.cpu_core.csr_file.mscratch[11] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold159 (.A(_08486_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold160 (.A(\soc_inst.spi_inst.tx_shift_reg[3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold161 (.A(_00160_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold162 (.A(\soc_inst.cpu_core.csr_file.mcause[28] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold163 (.A(\soc_inst.mem_ctrl.next_instr_data[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold164 (.A(_00658_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold165 (.A(\soc_inst.spi_inst.tx_shift_reg[5] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold166 (.A(_00162_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold167 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[5] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold168 (.A(_00838_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold169 (.A(\soc_inst.mem_ctrl.next_instr_data[28] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold170 (.A(_00686_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold171 (.A(\soc_inst.mem_ctrl.next_instr_data[31] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold172 (.A(_00689_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold173 (.A(\soc_inst.mem_ctrl.next_instr_data[22] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold174 (.A(_00680_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold175 (.A(\soc_inst.mem_ctrl.next_instr_data[29] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold176 (.A(_00687_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold177 (.A(\soc_inst.mem_ctrl.next_instr_data[15] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold178 (.A(_00673_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold179 (.A(\soc_inst.cpu_core.ex_rs1_data[4] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold180 (.A(_01294_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold181 (.A(\soc_inst.cpu_core.csr_file.mscratch[17] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold182 (.A(_08510_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold183 (.A(_00740_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold184 (.A(\soc_inst.mem_ctrl.next_instr_data[20] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold185 (.A(_00678_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold186 (.A(\soc_inst.mem_ctrl.spi_data_in[28] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold187 (.A(_00549_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold188 (.A(\soc_inst.core_instr_data[24] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold189 (.A(_00615_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold190 (.A(\soc_inst.cpu_core.csr_file.mcause[12] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold191 (.A(\soc_inst.spi_inst.tx_shift_reg[14] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold192 (.A(_00140_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold193 (.A(\soc_inst.cpu_core.ex_rs1_data[7] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold194 (.A(_01297_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold195 (.A(\soc_inst.spi_inst.tx_shift_reg[2] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold196 (.A(_00159_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold197 (.A(\soc_inst.core_instr_data[26] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold198 (.A(_00617_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold199 (.A(\soc_inst.mem_ctrl.spi_data_in[30] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold200 (.A(_00551_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold201 (.A(\soc_inst.i2c_inst.state[2] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold202 (.A(_06444_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold203 (.A(_01972_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold204 (.A(\soc_inst.mem_ctrl.next_instr_data[7] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold205 (.A(_00665_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold206 (.A(\soc_inst.cpu_core.csr_file.mscratch[20] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold207 (.A(_08522_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold208 (.A(_00743_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold209 (.A(\soc_inst.mem_ctrl.next_instr_data[14] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold210 (.A(_00672_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold211 (.A(\soc_inst.core_mem_rdata[2] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00625_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold213 (.A(\soc_inst.cpu_core.csr_file.mscratch[22] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold214 (.A(_08530_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold215 (.A(_00745_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold216 (.A(\soc_inst.core_mem_rdata[3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold217 (.A(_00626_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold218 (.A(\soc_inst.mem_ctrl.spi_data_in[24] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold219 (.A(_00545_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold220 (.A(\soc_inst.mem_ctrl.next_instr_data[25] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold221 (.A(_00683_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold222 (.A(\soc_inst.core_mem_rdata[5] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold223 (.A(\soc_inst.spi_inst.tx_shift_reg[8] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold224 (.A(_00165_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold225 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold226 (.A(_00842_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold227 (.A(\soc_inst.cpu_core.ex_rs1_data[5] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold228 (.A(_01295_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold229 (.A(\soc_inst.spi_inst.tx_shift_reg[23] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold230 (.A(_00150_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold231 (.A(\soc_inst.core_instr_data[21] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold232 (.A(_00612_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold233 (.A(\soc_inst.cpu_core.ex_rs2_data[19] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold234 (.A(_01373_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold235 (.A(\soc_inst.mem_ctrl.spi_data_in[26] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold236 (.A(_00547_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold237 (.A(\soc_inst.i2c_inst.clk_cnt[0] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold238 (.A(\soc_inst.cpu_core.ex_rs2_data[27] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold239 (.A(_01381_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold240 (.A(\soc_inst.cpu_core.csr_file.mcause[20] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold241 (.A(\soc_inst.core_instr_data[31] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold242 (.A(_00622_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold243 (.A(\soc_inst.core_instr_data[30] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold244 (.A(_00621_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold245 (.A(\soc_inst.spi_inst.tx_shift_reg[1] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold246 (.A(_00156_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold247 (.A(\soc_inst.spi_inst.tx_shift_reg[7] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold248 (.A(_00164_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold249 (.A(\soc_inst.mem_ctrl.spi_data_in[25] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold250 (.A(_00546_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold251 (.A(\soc_inst.spi_inst.tx_shift_reg[22] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold252 (.A(\soc_inst.gpio_inst.int_pend_reg[6] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold253 (.A(_05106_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold254 (.A(\soc_inst.mem_ctrl.next_instr_data[9] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold255 (.A(_00667_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold256 (.A(\soc_inst.mem_ctrl.spi_mem_inst.flash_in_cont_mode ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold257 (.A(_00845_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold258 (.A(\soc_inst.cpu_core.ex_rs2_data[0] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold259 (.A(_01354_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold260 (.A(\soc_inst.cpu_core.csr_file.mcause[30] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold261 (.A(\soc_inst.spi_inst.tx_shift_reg[28] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00155_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold263 (.A(\soc_inst.spi_inst.tx_shift_reg[24] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold264 (.A(_00151_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold265 (.A(\soc_inst.spi_inst.start_pending ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold266 (.A(_06932_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold267 (.A(\soc_inst.spi_inst.next_state[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold268 (.A(\soc_inst.mem_ctrl.spi_data_in[23] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold269 (.A(_00544_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold270 (.A(\soc_inst.spi_inst.tx_shift_reg[29] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold271 (.A(_00157_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold272 (.A(\soc_inst.cpu_core.ex_mem_we ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold273 (.A(_01418_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold274 (.A(\soc_inst.cpu_core.ex_rs1_data[6] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold275 (.A(_01296_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold276 (.A(\soc_inst.mem_ctrl.spi_data_in[31] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold277 (.A(_00552_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold278 (.A(\soc_inst.cpu_core.csr_file.mscratch[3] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold279 (.A(\soc_inst.gpio_inst.int_pend_reg[4] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold280 (.A(_05110_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold281 (.A(_01975_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold282 (.A(\soc_inst.mem_ctrl.spi_data_in[11] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold283 (.A(_00532_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold284 (.A(\soc_inst.core_instr_data[18] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00609_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold286 (.A(\soc_inst.cpu_core.ex_rs2_data[5] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold287 (.A(_01359_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold288 (.A(\soc_inst.spi_inst.tx_shift_reg[30] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold289 (.A(_00158_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold290 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold291 (.A(_00841_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold292 (.A(\soc_inst.core_instr_data[20] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold293 (.A(_00611_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold294 (.A(\soc_inst.cpu_core.ex_rs2_data[15] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold295 (.A(_01369_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold296 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[5] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold297 (.A(_05162_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold298 (.A(_02026_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold299 (.A(\soc_inst.mem_ctrl.spi_data_in[22] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold300 (.A(_00543_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold301 (.A(\soc_inst.spi_inst.tx_shift_reg[25] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold302 (.A(\soc_inst.gpio_inst.int_pend_reg[3] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold303 (.A(_05112_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold304 (.A(_01976_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold305 (.A(\soc_inst.core_mem_wdata[30] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold306 (.A(_02060_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold307 (.A(\soc_inst.spi_inst.tx_shift_reg[13] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold308 (.A(_00139_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold309 (.A(\soc_inst.cpu_core.csr_file.mtvec[5] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold310 (.A(_04974_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold311 (.A(\soc_inst.mem_ctrl.spi_data_in[2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold312 (.A(_00523_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold313 (.A(\soc_inst.core_instr_data[17] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold314 (.A(_00608_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold315 (.A(\soc_inst.spi_inst.tx_shift_reg[17] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold316 (.A(_00143_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold317 (.A(\soc_inst.core_instr_data[19] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold318 (.A(_00610_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold319 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold320 (.A(_00836_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold321 (.A(\soc_inst.cpu_core.ex_rs2_data[4] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold322 (.A(_01358_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold323 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold324 (.A(_00835_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold325 (.A(\soc_inst.mem_ctrl.next_instr_ready_reg ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold326 (.A(_07546_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00520_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold328 (.A(\soc_inst.mem_ctrl.spi_data_in[18] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold329 (.A(_00539_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold330 (.A(\soc_inst.mem_ctrl.spi_mem_inst.initialized ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold331 (.A(_06048_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold332 (.A(_06049_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold333 (.A(_00012_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold334 (.A(\soc_inst.mem_ctrl.spi_data_in[7] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold335 (.A(_00528_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold336 (.A(\soc_inst.mem_ctrl.spi_data_in[19] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold337 (.A(_00540_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold338 (.A(\soc_inst.cpu_core.csr_file.mtval[11] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold339 (.A(_01910_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold340 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold341 (.A(_00840_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold342 (.A(\soc_inst.spi_inst.tx_shift_reg[21] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold343 (.A(\soc_inst.cpu_core.csr_file.mcause[16] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold344 (.A(\soc_inst.core_mem_wdata[31] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold345 (.A(_02061_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold346 (.A(\soc_inst.cpu_core.ex_funct7[4] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold347 (.A(_01094_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold348 (.A(\soc_inst.cpu_core.csr_file.mcause[19] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold349 (.A(\soc_inst.mem_ctrl.spi_data_in[5] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold350 (.A(_00526_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold351 (.A(\soc_inst.mem_ctrl.spi_data_in[6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold352 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold353 (.A(_06133_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold354 (.A(\soc_inst.spi_inst.rx_shift_reg[31] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold355 (.A(_07118_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold356 (.A(\soc_inst.cpu_core.csr_file.mstatus[8] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold357 (.A(_00555_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold358 (.A(\soc_inst.mem_ctrl.spi_data_in[21] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00542_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold360 (.A(\soc_inst.spi_inst.tx_shift_reg[12] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold361 (.A(_00138_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold362 (.A(\soc_inst.cpu_core.csr_file.mcause[17] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold363 (.A(\soc_inst.cpu_core.csr_file.mcause[4] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold364 (.A(\soc_inst.spi_inst.tx_shift_reg[9] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold365 (.A(_00135_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold366 (.A(\soc_inst.cpu_core.ex_rs1_data[15] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold367 (.A(_01305_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold368 (.A(\soc_inst.cpu_core.csr_file.mstatus[6] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold369 (.A(_00554_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold370 (.A(\soc_inst.cpu_core.ex_funct7[5] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold371 (.A(_01095_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold372 (.A(\soc_inst.cpu_core.csr_file.mtvec[11] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold373 (.A(_04981_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold374 (.A(\soc_inst.core_instr_data[28] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold375 (.A(_00619_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold376 (.A(\soc_inst.cpu_core.register_file.registers[1][29] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold377 (.A(\soc_inst.cpu_core.csr_file.mtval[20] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold378 (.A(_01919_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold379 (.A(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold380 (.A(\soc_inst.cpu_core.csr_file.mtval[13] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold381 (.A(_01912_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold382 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold383 (.A(_00833_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold384 (.A(\soc_inst.cpu_core.csr_file.mstatus[10] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold385 (.A(_07625_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold386 (.A(_00557_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold387 (.A(\soc_inst.mem_ctrl.spi_data_in[1] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold388 (.A(_00522_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold389 (.A(\soc_inst.gpio_inst.int_pend_reg[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold390 (.A(_07129_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold391 (.A(_00400_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold392 (.A(\soc_inst.cpu_core.csr_file.mstatus[5] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold393 (.A(_00553_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold394 (.A(\soc_inst.cpu_core.csr_file.mstatus[24] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold395 (.A(_02107_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold396 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold397 (.A(_00003_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold398 (.A(\soc_inst.cpu_core.csr_file.mtval[9] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold399 (.A(_01908_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold400 (.A(\soc_inst.cpu_core.csr_file.mstatus[9] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold401 (.A(_00556_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold402 (.A(\soc_inst.core_mem_wdata[27] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold403 (.A(_02057_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold404 (.A(\soc_inst.spi_inst.tx_shift_reg[27] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold405 (.A(\soc_inst.gpio_inst.int_pend_reg[2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold406 (.A(_05114_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold407 (.A(_01977_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold408 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold409 (.A(\soc_inst.cpu_core.register_file.registers[1][14] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold410 (.A(\soc_inst.mem_ctrl.spi_data_in[15] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold411 (.A(_00536_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold412 (.A(\soc_inst.spi_inst.clk_counter[0] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold413 (.A(_00124_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold414 (.A(\soc_inst.i2c_inst.shift_reg[4] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold415 (.A(_00082_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold416 (.A(\soc_inst.spi_inst.clk_counter[1] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold417 (.A(_00125_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold418 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold419 (.A(\soc_inst.cpu_core.ex_rs2_data[24] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold420 (.A(_01378_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold421 (.A(\soc_inst.cpu_core.csr_file.mtvec[3] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold422 (.A(\soc_inst.core_mem_rdata[30] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold423 (.A(_00653_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold424 (.A(\soc_inst.spi_inst.clk_counter[7] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold425 (.A(_00131_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold426 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold427 (.A(_06123_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold428 (.A(\soc_inst.cpu_core.csr_file.mtvec[8] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold429 (.A(_04978_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold430 (.A(\soc_inst.cpu_core.ex_branch_target[15] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold431 (.A(\soc_inst.cpu_core.csr_file.mtval[17] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold432 (.A(_01916_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold433 (.A(\soc_inst.cpu_core.csr_file.mcause[13] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold434 (.A(\soc_inst.cpu_core.register_file.registers[1][4] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold435 (.A(\soc_inst.gpio_inst.int_pend_reg[1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold436 (.A(_05116_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold437 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold438 (.A(_00777_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold439 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[0] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold440 (.A(_05207_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold441 (.A(_02071_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold442 (.A(\soc_inst.spi_inst.state[1] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold443 (.A(\soc_inst.spi_inst.next_state[1] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold444 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold445 (.A(_05346_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold446 (.A(_02132_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold447 (.A(\soc_inst.cpu_core.error_flag_reg ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold448 (.A(\soc_inst.cpu_core.ex_mem_re ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold449 (.A(_00024_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold450 (.A(\soc_inst.core_instr_data[22] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold451 (.A(_00613_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold452 (.A(\soc_inst.mem_ctrl.spi_data_in[4] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold453 (.A(_00525_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold454 (.A(\soc_inst.core_mem_wdata[26] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold455 (.A(_02056_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold456 (.A(\soc_inst.mem_ctrl.spi_data_in[14] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold457 (.A(_00535_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold458 (.A(\soc_inst.i2c_inst.shift_reg[5] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold459 (.A(_00083_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold460 (.A(\soc_inst.cpu_core.csr_file.mtvec[14] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold461 (.A(_04984_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold462 (.A(_01940_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold463 (.A(\soc_inst.cpu_core.id_instr[5] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold464 (.A(_09218_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold465 (.A(\soc_inst.core_instr_data[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold466 (.A(_00592_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold467 (.A(\soc_inst.i2c_inst.shift_reg[1] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold468 (.A(_00079_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold469 (.A(\soc_inst.cpu_core.csr_file.mtvec[7] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold470 (.A(\soc_inst.cpu_core.register_file.registers[1][9] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold471 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[18] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold472 (.A(_00774_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold473 (.A(\soc_inst.core_mem_rdata[21] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold474 (.A(_00644_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold475 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold476 (.A(_00764_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold477 (.A(\soc_inst.cpu_core.register_file.registers[1][15] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold478 (.A(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold479 (.A(\soc_inst.mem_ctrl.spi_data_in[13] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00534_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold481 (.A(\soc_inst.spi_inst.tx_shift_reg[4] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold482 (.A(_00161_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold483 (.A(\soc_inst.cpu_core.register_file.registers[1][21] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold484 (.A(\soc_inst.gpio_inst.int_pend_reg[5] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold485 (.A(_05108_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold486 (.A(_01974_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold487 (.A(\soc_inst.mem_ctrl.spi_data_in[9] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold488 (.A(_00530_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold489 (.A(\soc_inst.cpu_core.id_imm12[9] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold490 (.A(\soc_inst.cpu_core.if_instr[8] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold491 (.A(_09567_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold492 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg_0 ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold493 (.A(_02147_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold494 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[7] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold495 (.A(_05206_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold496 (.A(\soc_inst.cpu_core.ex_is_ecall ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00914_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold498 (.A(\soc_inst.cpu_core.csr_file.mtval[19] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold499 (.A(_01918_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold500 (.A(\soc_inst.cpu_core.csr_file.mtval[7] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold501 (.A(_01906_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold502 (.A(\soc_inst.mem_ctrl.spi_data_in[12] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold503 (.A(_00533_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold504 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold505 (.A(\soc_inst.cpu_core.id_imm12[10] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold506 (.A(\soc_inst.spi_inst.clk_counter[2] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold507 (.A(_00126_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold508 (.A(\soc_inst.cpu_core.mem_instr[5] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold509 (.A(_01074_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold510 (.A(\soc_inst.mem_ctrl.spi_data_in[3] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold511 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold512 (.A(_00766_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold513 (.A(\soc_inst.core_mem_rdata[8] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold514 (.A(\soc_inst.i2c_inst.bit_cnt[0] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold515 (.A(\soc_inst.core_mem_rdata[12] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold516 (.A(\soc_inst.core_mem_rdata[9] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold517 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold518 (.A(_00776_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold519 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[4] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold520 (.A(_02127_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold521 (.A(\soc_inst.mem_ctrl.spi_read_enable ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold522 (.A(_00655_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold523 (.A(\soc_inst.cpu_core.csr_file.mtval[5] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold524 (.A(_01904_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold525 (.A(_00272_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold526 (.A(_01073_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold527 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[0] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold528 (.A(_02115_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold529 (.A(\soc_inst.core_mem_rdata[11] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold530 (.A(\soc_inst.spi_inst.rx_shift_reg[21] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold531 (.A(_07108_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold532 (.A(\soc_inst.core_mem_wdata[28] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold533 (.A(_02058_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold534 (.A(\soc_inst.mem_ctrl.spi_data_in[20] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold535 (.A(_00541_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold536 (.A(\soc_inst.cpu_core.csr_file.mtval[6] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold537 (.A(_01905_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold538 (.A(\soc_inst.cpu_core.ex_reg_we ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold539 (.A(_00879_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold540 (.A(\soc_inst.cpu_core.csr_file.mtvec[16] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold541 (.A(_01942_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold542 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[1] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold543 (.A(_05334_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold544 (.A(\soc_inst.spi_inst.done ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold545 (.A(_07127_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold546 (.A(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold547 (.A(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold548 (.A(\soc_inst.cpu_core.register_file.registers[1][17] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold549 (.A(\soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold550 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold551 (.A(_00772_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold552 (.A(\soc_inst.cpu_core.ex_branch_target[4] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold553 (.A(\soc_inst.cpu_core.csr_file.mtvec[19] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold554 (.A(_01945_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold555 (.A(\soc_inst.core_mem_addr[29] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold556 (.A(_01351_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold557 (.A(\soc_inst.core_mem_rdata[22] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold558 (.A(_00645_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold559 (.A(\soc_inst.cpu_core.ex_rs1_data[11] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold560 (.A(_00984_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold561 (.A(\soc_inst.core_mem_rdata[27] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold562 (.A(_00650_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold563 (.A(\soc_inst.mem_ctrl.instr_ready_reg ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold564 (.A(_00657_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold565 (.A(\soc_inst.cpu_core.csr_file.mie[11] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold566 (.A(_01869_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold567 (.A(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold568 (.A(_00170_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold569 (.A(\soc_inst.cpu_core.ex_rs1_data[22] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold570 (.A(_01312_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold571 (.A(\soc_inst.spi_inst.rx_shift_reg[24] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold572 (.A(_07111_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold573 (.A(\soc_inst.core_mem_rdata[14] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold574 (.A(\soc_inst.i2c_inst.shift_reg[3] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold575 (.A(_00081_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold576 (.A(\soc_inst.cpu_core.register_file.registers[1][28] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold577 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[3] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold578 (.A(_05337_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold579 (.A(_02126_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold580 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold581 (.A(_02116_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold582 (.A(\soc_inst.cpu_core.mem_rs1_data[4] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold583 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold584 (.A(_05326_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold585 (.A(_02118_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold586 (.A(\soc_inst.cpu_core.csr_file.mtvec[9] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold587 (.A(_04979_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold588 (.A(_01935_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold589 (.A(\soc_inst.cpu_core.if_instr[10] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00926_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold591 (.A(\soc_inst.i2c_inst.shift_reg[0] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold592 (.A(_00078_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold593 (.A(\soc_inst.mem_ctrl.spi_data_in[8] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold594 (.A(_00529_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold595 (.A(\soc_inst.cpu_core.register_file.registers[1][2] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold596 (.A(\soc_inst.core_mem_rdata[13] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold597 (.A(\soc_inst.cpu_core.i_mem_ready ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold598 (.A(_00656_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold599 (.A(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold600 (.A(\soc_inst.cpu_core.csr_file.mie[7] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold601 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold602 (.A(_02119_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold603 (.A(\soc_inst.spi_inst.rx_shift_reg[28] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold604 (.A(_07115_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold605 (.A(\soc_inst.cpu_core.register_file.registers[1][24] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold606 (.A(\soc_inst.cpu_core.register_file.registers[2][28] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold607 (.A(\soc_inst.cpu_core.register_file.registers[14][12] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold608 (.A(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold609 (.A(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold610 (.A(\soc_inst.cpu_core.register_file.registers[6][0] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold611 (.A(\soc_inst.core_instr_data[8] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold612 (.A(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold613 (.A(_06620_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold614 (.A(\soc_inst.mem_ctrl.spi_data_in[17] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold615 (.A(_00538_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold616 (.A(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold617 (.A(_00210_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold618 (.A(\soc_inst.mem_ctrl.spi_data_in[0] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold619 (.A(_00521_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold620 (.A(\soc_inst.cpu_core.register_file.registers[5][22] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold621 (.A(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold622 (.A(\soc_inst.mem_ctrl.spi_data_in[16] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold623 (.A(_00537_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold624 (.A(\soc_inst.cpu_core.register_file.registers[11][25] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold625 (.A(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold626 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold627 (.A(_00771_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold628 (.A(\soc_inst.cpu_core.if_instr[11] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold629 (.A(\soc_inst.cpu_core.ex_rs2_data[8] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold630 (.A(_01362_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold631 (.A(\soc_inst.spi_inst.rx_shift_reg[25] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold632 (.A(\soc_inst.i2c_inst.clk_cnt[2] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold633 (.A(_06475_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold634 (.A(_00072_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold635 (.A(\soc_inst.cpu_core.ex_rs2_data[29] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold636 (.A(_00911_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold637 (.A(\soc_inst.cpu_core.register_file.registers[1][13] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold638 (.A(\soc_inst.cpu_core.register_file.registers[5][27] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold639 (.A(\soc_inst.cpu_core.ex_rs2_data[10] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold640 (.A(_01364_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold641 (.A(\soc_inst.cpu_core.register_file.registers[1][26] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold642 (.A(\soc_inst.cpu_core.id_imm12[5] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold643 (.A(_01259_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold644 (.A(\soc_inst.cpu_core.register_file.registers[9][27] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold645 (.A(\soc_inst.cpu_core.register_file.registers[1][18] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold646 (.A(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold647 (.A(_00205_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold648 (.A(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold649 (.A(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold650 (.A(\soc_inst.cpu_core.register_file.registers[11][27] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold651 (.A(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold652 (.A(\soc_inst.cpu_core.ex_rs1_data[21] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold653 (.A(_01311_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold654 (.A(\soc_inst.cpu_core.register_file.registers[1][3] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold655 (.A(\soc_inst.cpu_core.csr_file.mtvec[17] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold656 (.A(_01943_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold657 (.A(\soc_inst.cpu_core.register_file.registers[2][16] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold658 (.A(\soc_inst.cpu_core.ex_alu_result[20] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold659 (.A(\soc_inst.cpu_core.ex_rs1_data[19] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold660 (.A(_01309_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold661 (.A(\soc_inst.cpu_core.register_file.registers[1][23] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold662 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold663 (.A(_00779_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold664 (.A(\soc_inst.cpu_core.ex_funct7[0] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold665 (.A(_01090_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold666 (.A(\soc_inst.cpu_core.register_file.registers[11][13] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold667 (.A(\soc_inst.core_mem_rdata[19] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold668 (.A(_00642_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold669 (.A(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold670 (.A(\soc_inst.spi_inst.tx_shift_reg[31] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold671 (.A(_07074_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold672 (.A(_00349_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold673 (.A(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold674 (.A(\soc_inst.cpu_core.csr_file.mtvec[1] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold675 (.A(\soc_inst.core_mem_rdata[20] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold676 (.A(_00643_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold677 (.A(\soc_inst.cpu_core.ex_rs1_data[23] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold678 (.A(_01313_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold679 (.A(\soc_inst.cpu_core.register_file.registers[8][30] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold680 (.A(\soc_inst.cpu_core.register_file.registers[9][0] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold681 (.A(\soc_inst.cpu_core.csr_file.mscratch[4] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold682 (.A(_00828_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold683 (.A(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold684 (.A(\soc_inst.core_mem_rdata[7] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold685 (.A(_00630_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold686 (.A(\soc_inst.cpu_core.id_rs1_data[11] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold687 (.A(\soc_inst.cpu_core.register_file.registers[6][28] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold688 (.A(\soc_inst.cpu_core.register_file.registers[8][2] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold689 (.A(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold690 (.A(\soc_inst.cpu_core.register_file.registers[1][19] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold691 (.A(\soc_inst.cpu_core.register_file.registers[1][22] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold692 (.A(\soc_inst.core_mem_wdata[15] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold693 (.A(\soc_inst.cpu_core.register_file.registers[11][21] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold694 (.A(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold695 (.A(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold696 (.A(\soc_inst.cpu_core.mem_rs1_data[3] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold697 (.A(_00976_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold698 (.A(\soc_inst.spi_inst.rx_shift_reg[20] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold699 (.A(_07107_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold700 (.A(\soc_inst.mem_ctrl.spi_data_in[10] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold701 (.A(_00531_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold702 (.A(\soc_inst.cpu_core.ex_rs1_data[13] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold703 (.A(_01303_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold704 (.A(\soc_inst.cpu_core.register_file.registers[13][1] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold705 (.A(\soc_inst.cpu_core.ex_rs2_data[3] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold706 (.A(_00885_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold707 (.A(\soc_inst.cpu_core.register_file.registers[9][4] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold708 (.A(\soc_inst.cpu_core.register_file.registers[10][14] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold709 (.A(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold710 (.A(\soc_inst.spi_inst.rx_shift_reg[22] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold711 (.A(\soc_inst.cpu_core.csr_file.mepc[13] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold712 (.A(_01958_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold713 (.A(\soc_inst.cpu_core.register_file.registers[13][6] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold714 (.A(\soc_inst.cpu_core.register_file.registers[12][28] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold715 (.A(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold716 (.A(_00200_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold717 (.A(\soc_inst.cpu_core.register_file.registers[15][28] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold718 (.A(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold719 (.A(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold720 (.A(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold721 (.A(\soc_inst.cpu_core.register_file.registers[9][3] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold722 (.A(\soc_inst.cpu_core.register_file.registers[9][5] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold723 (.A(\soc_inst.cpu_core.ex_rs1_data[2] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold724 (.A(_01292_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold725 (.A(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold726 (.A(\soc_inst.cpu_core.register_file.registers[5][25] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold727 (.A(\soc_inst.cpu_core.register_file.registers[10][27] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold728 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold729 (.A(_00767_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold730 (.A(\soc_inst.cpu_core.ex_rs1_data[1] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold731 (.A(_00974_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold732 (.A(\soc_inst.cpu_core.mem_instr[15] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold733 (.A(_01080_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold734 (.A(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold735 (.A(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold736 (.A(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold737 (.A(\soc_inst.cpu_core.register_file.registers[2][2] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold738 (.A(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold739 (.A(\soc_inst.spi_inst.bit_counter[1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold740 (.A(_07076_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold741 (.A(_00351_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold742 (.A(\soc_inst.cpu_core.register_file.registers[4][23] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold743 (.A(\soc_inst.cpu_core.mem_instr[3] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold744 (.A(_01072_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold745 (.A(\soc_inst.cpu_core.register_file.registers[3][19] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold746 (.A(\soc_inst.i2c_inst.stop_pending ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold747 (.A(_00086_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold748 (.A(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold749 (.A(_00213_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold750 (.A(\soc_inst.cpu_core.register_file.registers[9][22] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold751 (.A(\soc_inst.cpu_core.register_file.registers[5][1] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold752 (.A(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold753 (.A(\soc_inst.cpu_core.register_file.registers[6][2] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold754 (.A(\soc_inst.cpu_core.csr_file.mepc[15] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold755 (.A(_01960_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold756 (.A(\soc_inst.cpu_core.register_file.registers[9][26] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold757 (.A(\soc_inst.cpu_core.ex_rs1_data[14] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold758 (.A(_01304_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold759 (.A(\soc_inst.cpu_core.csr_file.mtvec[6] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold760 (.A(_01932_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold761 (.A(\soc_inst.cpu_core.register_file.registers[11][2] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold762 (.A(\soc_inst.cpu_core.register_file.registers[5][28] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold763 (.A(\soc_inst.cpu_core.id_instr[10] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold764 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[6] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold765 (.A(\soc_inst.cpu_core.csr_file.mscratch[2] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold766 (.A(\soc_inst.cpu_core.register_file.registers[2][10] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold767 (.A(\soc_inst.cpu_core.register_file.registers[5][2] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold768 (.A(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold769 (.A(\soc_inst.cpu_core.ex_rs1_data[29] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold770 (.A(_01319_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold771 (.A(_00270_),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold772 (.A(_01069_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold773 (.A(\soc_inst.cpu_core.register_file.registers[8][11] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold774 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold775 (.A(_00773_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold776 (.A(\soc_inst.cpu_core.alu.b[14] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold777 (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold778 (.A(_01088_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold779 (.A(\soc_inst.cpu_core.ex_rs1_data[3] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold780 (.A(_01293_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold781 (.A(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold782 (.A(_01275_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold783 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold784 (.A(_00765_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold785 (.A(\soc_inst.cpu_core.ex_rs2_data[31] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold786 (.A(_01385_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold787 (.A(\soc_inst.cpu_core.register_file.registers[2][0] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold788 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[28] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold789 (.A(_08430_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold790 (.A(\soc_inst.cpu_core.register_file.registers[9][8] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold791 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold792 (.A(_05214_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold793 (.A(_02074_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold794 (.A(\soc_inst.cpu_core.register_file.registers[1][0] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold795 (.A(\soc_inst.cpu_core.ex_rs1_data[18] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold796 (.A(_01308_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold797 (.A(\soc_inst.cpu_core.id_rs2_data[3] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold798 (.A(\soc_inst.cpu_core.register_file.registers[15][16] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold799 (.A(\soc_inst.cpu_core.ex_rs1_data[25] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold800 (.A(_01315_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold801 (.A(\soc_inst.cpu_core.register_file.registers[1][5] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold802 (.A(\soc_inst.cpu_core.register_file.registers[9][29] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold803 (.A(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold804 (.A(\soc_inst.pwm_inst.channel_duty[0][7] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold805 (.A(_00459_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold806 (.A(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold807 (.A(_00215_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold808 (.A(\soc_inst.cpu_core.register_file.registers[10][23] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold809 (.A(\soc_inst.cpu_core.ex_exception_pc[13] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold810 (.A(_01279_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold811 (.A(\soc_inst.cpu_core.register_file.registers[15][13] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold812 (.A(\soc_inst.spi_inst.rx_shift_reg[29] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold813 (.A(\soc_inst.cpu_core.register_file.registers[12][22] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold814 (.A(\soc_inst.cpu_core.register_file.registers[11][4] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold815 (.A(\soc_inst.cpu_core.register_file.registers[13][18] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold816 (.A(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold817 (.A(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold818 (.A(\soc_inst.cpu_core.ex_rs2_data[1] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold819 (.A(_00883_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold820 (.A(\soc_inst.cpu_core.ex_alu_result[19] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold821 (.A(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold822 (.A(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold823 (.A(\soc_inst.cpu_core.register_file.registers[15][9] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold824 (.A(\soc_inst.core_mem_rdata[23] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold825 (.A(_00646_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold826 (.A(\soc_inst.cpu_core.register_file.registers[12][8] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold827 (.A(\soc_inst.cpu_core.if_instr[7] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold828 (.A(_09566_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold829 (.A(\soc_inst.cpu_core.register_file.registers[4][0] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold830 (.A(\soc_inst.cpu_core.register_file.registers[4][9] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold831 (.A(\soc_inst.cpu_core.register_file.registers[2][26] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold832 (.A(\soc_inst.pwm_inst.channel_counter[1][2] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold833 (.A(_06532_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold834 (.A(_00115_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold835 (.A(\soc_inst.cpu_core.register_file.registers[9][21] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold836 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold837 (.A(_00770_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold838 (.A(\soc_inst.cpu_core.ex_rs1_data[28] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold839 (.A(_01001_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold840 (.A(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold841 (.A(_01277_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold842 (.A(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold843 (.A(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold844 (.A(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold845 (.A(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold846 (.A(\soc_inst.cpu_core.register_file.registers[13][20] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold847 (.A(\soc_inst.cpu_core.csr_file.mepc[22] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold848 (.A(_01967_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold849 (.A(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold850 (.A(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold851 (.A(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold852 (.A(\soc_inst.cpu_core.csr_file.mtvec[15] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold853 (.A(_01941_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold854 (.A(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold855 (.A(\soc_inst.i2c_inst.ctrl_reg[4] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold856 (.A(\soc_inst.cpu_core.ex_rs1_data[27] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold857 (.A(_01000_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold858 (.A(\soc_inst.cpu_core.ex_branch_target[26] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold859 (.A(_01896_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold860 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[2] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold861 (.A(_00020_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold862 (.A(\soc_inst.cpu_core.ex_rs2_data[9] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold863 (.A(_01363_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold864 (.A(\soc_inst.cpu_core.id_rs1_data[27] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold865 (.A(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold866 (.A(_01273_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold867 (.A(\soc_inst.cpu_core.csr_file.mtvec[13] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold868 (.A(_01939_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold869 (.A(\soc_inst.core_instr_data[9] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold870 (.A(_00600_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold871 (.A(\soc_inst.cpu_core.csr_file.mtvec[10] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold872 (.A(_01936_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold873 (.A(\soc_inst.cpu_core.register_file.registers[4][24] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold874 (.A(\soc_inst.i2c_inst.bit_cnt[1] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold875 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[23] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold876 (.A(_08429_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold877 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold878 (.A(_00775_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold879 (.A(\soc_inst.core_mem_wdata[4] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold880 (.A(\soc_inst.cpu_core.register_file.registers[9][12] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold881 (.A(\soc_inst.cpu_core.mem_rs1_data[2] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold882 (.A(\soc_inst.cpu_core.id_instr[7] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold883 (.A(_01241_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold884 (.A(\soc_inst.core_mem_wdata[24] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold885 (.A(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold886 (.A(\soc_inst.cpu_core.register_file.registers[9][28] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold887 (.A(\soc_inst.cpu_core.register_file.registers[3][22] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold888 (.A(\soc_inst.cpu_core.register_file.registers[3][15] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold889 (.A(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold890 (.A(_00202_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold891 (.A(\soc_inst.cpu_core.register_file.registers[13][22] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold892 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[31] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold893 (.A(_08433_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold894 (.A(\soc_inst.cpu_core.register_file.registers[10][26] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold895 (.A(\soc_inst.cpu_core.register_file.registers[9][19] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold896 (.A(\soc_inst.spi_inst.rx_shift_reg[27] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold897 (.A(_07114_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold898 (.A(\soc_inst.cpu_core.register_file.registers[14][20] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold899 (.A(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold900 (.A(\soc_inst.cpu_core.if_pc[2] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold901 (.A(_00950_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold902 (.A(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold903 (.A(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold904 (.A(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold905 (.A(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold906 (.A(\soc_inst.cpu_core.register_file.registers[13][12] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold907 (.A(\soc_inst.cpu_core.register_file.registers[8][23] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold908 (.A(\soc_inst.cpu_core.register_file.registers[1][1] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold909 (.A(\soc_inst.cpu_core.register_file.registers[3][7] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold910 (.A(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold911 (.A(\soc_inst.core_mem_rdata[10] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold912 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[2] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold913 (.A(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold914 (.A(\soc_inst.cpu_core.register_file.registers[13][27] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold915 (.A(\soc_inst.cpu_core.id_imm[31] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold916 (.A(_01160_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold917 (.A(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold918 (.A(\soc_inst.cpu_core.register_file.registers[8][19] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold919 (.A(\soc_inst.cpu_core.register_file.registers[5][24] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold920 (.A(\soc_inst.cpu_core.alu.a[2] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold921 (.A(\soc_inst.cpu_core.csr_file.mepc[9] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold922 (.A(_01954_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold923 (.A(\soc_inst.cpu_core.register_file.registers[5][7] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold924 (.A(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold925 (.A(\soc_inst.cpu_core.id_instr[17] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold926 (.A(_01251_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold927 (.A(\soc_inst.cpu_core.mem_rs1_data[25] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold928 (.A(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold929 (.A(\soc_inst.cpu_core.register_file.registers[3][12] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold930 (.A(\soc_inst.cpu_core.register_file.registers[5][30] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold931 (.A(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold932 (.A(\soc_inst.cpu_core.register_file.registers[6][30] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold933 (.A(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold934 (.A(\soc_inst.core_mem_wdata[9] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold935 (.A(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold936 (.A(\soc_inst.cpu_core.register_file.registers[10][10] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold937 (.A(\soc_inst.cpu_core.register_file.registers[5][15] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold938 (.A(\soc_inst.cpu_core.csr_file.mepc[8] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold939 (.A(_01953_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold940 (.A(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold941 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[2] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold942 (.A(_02117_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold943 (.A(\soc_inst.core_mem_wdata[19] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold944 (.A(_02049_),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold945 (.A(\soc_inst.core_mem_wdata[5] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold946 (.A(\soc_inst.spi_inst.rx_shift_reg[23] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold947 (.A(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold948 (.A(_07064_),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold949 (.A(\soc_inst.cpu_core.register_file.registers[1][16] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold950 (.A(\soc_inst.cpu_core.register_file.registers[4][5] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold951 (.A(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold952 (.A(\soc_inst.cpu_core.id_rs1_data[28] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold953 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold954 (.A(_00769_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold955 (.A(_00295_),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold956 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold957 (.A(_00014_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold958 (.A(\soc_inst.core_mem_wdata[7] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold959 (.A(\soc_inst.cpu_core.ex_branch_target[5] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold960 (.A(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold961 (.A(\soc_inst.cpu_core.register_file.registers[6][14] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold962 (.A(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold963 (.A(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold964 (.A(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold965 (.A(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold966 (.A(\soc_inst.cpu_core.register_file.registers[5][21] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold967 (.A(\soc_inst.cpu_core.register_file.registers[14][14] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold968 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[30] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold969 (.A(_08432_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold970 (.A(\soc_inst.cpu_core.id_instr[15] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold971 (.A(_01249_),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold972 (.A(\soc_inst.cpu_core.register_file.registers[5][8] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold973 (.A(\soc_inst.cpu_core.register_file.registers[4][31] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold974 (.A(\soc_inst.cpu_core.register_file.registers[2][25] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold975 (.A(\soc_inst.cpu_core.register_file.registers[10][8] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold976 (.A(_00229_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold977 (.A(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold978 (.A(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold979 (.A(\soc_inst.cpu_core.id_rs2_data[1] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold980 (.A(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold981 (.A(\soc_inst.cpu_core.register_file.registers[4][13] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold982 (.A(\soc_inst.cpu_core.register_file.registers[10][0] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold983 (.A(\soc_inst.cpu_core.id_imm[11] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold984 (.A(_02396_),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold985 (.A(_01140_),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold986 (.A(\soc_inst.cpu_core.id_instr[18] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold987 (.A(_09577_),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold988 (.A(\soc_inst.cpu_core.ex_rs2_data[16] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold989 (.A(_00898_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold990 (.A(\soc_inst.cpu_core.register_file.registers[14][10] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold991 (.A(\soc_inst.cpu_core.ex_branch_target[23] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold992 (.A(\soc_inst.cpu_core.ex_exception_pc[2] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold993 (.A(_01268_),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold994 (.A(\soc_inst.cpu_core.csr_file.mtvec[12] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold995 (.A(_01938_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold996 (.A(\soc_inst.cpu_core.mem_instr[19] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold997 (.A(_01084_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold998 (.A(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold999 (.A(\soc_inst.cpu_core.register_file.registers[3][20] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\soc_inst.spi_inst.rx_shift_reg[26] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\soc_inst.cpu_core.register_file.registers[14][1] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\soc_inst.cpu_core.register_file.registers[5][20] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\soc_inst.cpu_core.register_file.registers[5][26] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\soc_inst.cpu_core.ex_rs2_data[18] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold1008 (.A(_01372_),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\soc_inst.cpu_core.register_file.registers[6][13] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\soc_inst.cpu_core.csr_file.mepc[5] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_01950_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\soc_inst.cpu_core.register_file.registers[6][29] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold1016 (.A(_00207_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\soc_inst.cpu_core.mem_rs1_data[29] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold1019 (.A(_08419_),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\soc_inst.cpu_core.register_file.registers[12][11] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\soc_inst.cpu_core.ex_rs2_data[12] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_00894_),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\soc_inst.cpu_core.csr_file.mepc[18] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_01963_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\soc_inst.cpu_core.ex_branch_target[14] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\soc_inst.cpu_core.ex_alu_result[16] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\soc_inst.cpu_core.register_file.registers[11][11] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[0] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold1037 (.A(_05335_),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_02124_),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\soc_inst.cpu_core.register_file.registers[9][17] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\soc_inst.cpu_core.register_file.registers[9][7] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\soc_inst.i2c_inst.bit_cnt[3] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold1045 (.A(_00416_),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\soc_inst.cpu_core.register_file.registers[8][27] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\soc_inst.cpu_core.register_file.registers[6][11] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\soc_inst.cpu_core.if_instr[15] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\soc_inst.cpu_core.register_file.registers[10][2] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\soc_inst.cpu_core.ex_alu_result[18] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\soc_inst.cpu_core.register_file.registers[8][26] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\soc_inst.cpu_core.alu.a[23] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_01189_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold1054 (.A(_00309_),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_02044_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\soc_inst.cpu_core.register_file.registers[11][22] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\soc_inst.cpu_core.register_file.registers[5][12] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\soc_inst.core_instr_data[29] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\soc_inst.cpu_core.ex_rs1_data[16] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_00989_),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\soc_inst.cpu_core.register_file.registers[12][29] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\soc_inst.cpu_core.register_file.registers[10][16] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\soc_inst.cpu_core.register_file.registers[2][7] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\soc_inst.cpu_core.register_file.registers[12][21] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\soc_inst.cpu_core.ex_rs1_data[8] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold1067 (.A(_01298_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\soc_inst.cpu_core.ex_rs2_data[6] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_00888_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\soc_inst.cpu_core.register_file.registers[10][18] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\soc_inst.cpu_core.register_file.registers[6][12] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\soc_inst.cpu_core.register_file.registers[8][0] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\soc_inst.cpu_core.register_file.registers[4][12] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\soc_inst.cpu_core.register_file.registers[4][2] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[5] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\soc_inst.cpu_core.register_file.registers[8][7] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[1] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\soc_inst.cpu_core.ex_branch_target[24] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_01894_),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\soc_inst.cpu_core.alu.b[5] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold1082 (.A(_01203_),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\soc_inst.cpu_core.ex_exception_pc[15] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold1084 (.A(_01281_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\soc_inst.cpu_core.register_file.registers[10][30] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\soc_inst.cpu_core.ex_exception_pc[14] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold1089 (.A(_01280_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_00171_),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\soc_inst.core_mem_wdata[18] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\soc_inst.cpu_core.register_file.registers[1][10] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\soc_inst.cpu_core.ex_rs2_data[25] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold1095 (.A(_00907_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\soc_inst.cpu_core.ex_rs2_data[21] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_00903_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\soc_inst.cpu_core.register_file.registers[5][31] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\soc_inst.core_mem_rdata[29] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold1102 (.A(_00652_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\soc_inst.cpu_core.register_file.registers[11][1] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_00296_),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\soc_inst.i2c_inst.shift_reg[7] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold1106 (.A(_07166_),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold1107 (.A(_07168_),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\soc_inst.cpu_core.register_file.registers[6][10] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_00304_),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\soc_inst.pwm_inst.channel_duty[1][10] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold1111 (.A(_00343_),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\soc_inst.cpu_core.register_file.registers[9][24] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\soc_inst.cpu_core.register_file.registers[1][31] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\soc_inst.cpu_core.register_file.registers[14][23] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_01278_),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\soc_inst.cpu_core.csr_file.mtvec[18] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold1120 (.A(_01944_),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\soc_inst.cpu_core.csr_file.mtvec[23] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold1122 (.A(_01949_),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\soc_inst.cpu_core.ex_rs2_data[7] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\soc_inst.core_mem_wdata[0] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\soc_inst.spi_inst.rx_shift_reg[18] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold1126 (.A(_07105_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_01274_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\soc_inst.cpu_core.csr_file.mepc[10] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold1131 (.A(_01955_),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\soc_inst.cpu_core.register_file.registers[11][23] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\soc_inst.core_instr_data[7] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\soc_inst.cpu_core.register_file.registers[9][15] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\soc_inst.cpu_core.ex_rs1_data[0] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold1136 (.A(_01290_),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\soc_inst.cpu_core.register_file.registers[11][30] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_00311_),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold1140 (.A(_02046_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\soc_inst.cpu_core.register_file.registers[4][21] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\soc_inst.cpu_core.register_file.registers[4][8] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_00245_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\soc_inst.cpu_core.ex_alu_result[29] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\soc_inst.cpu_core.register_file.registers[2][15] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\soc_inst.cpu_core.register_file.registers[12][9] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\soc_inst.cpu_core.register_file.registers[13][9] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_00299_),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\soc_inst.pwm_inst.channel_counter[1][15] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_06555_),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\soc_inst.cpu_core.register_file.registers[9][6] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\soc_inst.cpu_core.if_instr[17] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\soc_inst.cpu_core.register_file.registers[11][12] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\soc_inst.cpu_core.register_file.registers[2][24] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\soc_inst.cpu_core.id_instr[19] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold1165 (.A(_01253_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold1167 (.A(_00197_),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\soc_inst.cpu_core.ex_exception_pc[18] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_01284_),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\soc_inst.cpu_core.id_rs2_data[25] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\soc_inst.spi_inst.rx_shift_reg[30] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\soc_inst.cpu_core.id_rs1_data[1] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\soc_inst.cpu_core.id_imm[19] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_01148_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\soc_inst.cpu_core.id_instr[11] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\soc_inst.cpu_core.register_file.registers[3][27] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\soc_inst.cpu_core.register_file.registers[2][27] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\soc_inst.cpu_core.ex_rs1_data[24] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold1179 (.A(_00997_),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\soc_inst.cpu_core.csr_file.mscratch[30] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_00753_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\soc_inst.cpu_core.register_file.registers[2][21] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\soc_inst.cpu_core.id_rs2_data[6] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00214_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\soc_inst.cpu_core.ex_rs2_data[2] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold1188 (.A(_00884_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\soc_inst.cpu_core.register_file.registers[1][6] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\soc_inst.cpu_core.register_file.registers[1][25] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\soc_inst.cpu_core.register_file.registers[13][3] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\soc_inst.cpu_core.register_file.registers[3][28] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\soc_inst.cpu_core.csr_file.mtval[16] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_01915_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\soc_inst.cpu_core.register_file.registers[10][25] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_02122_),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\soc_inst.cpu_core.register_file.registers[1][20] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_00251_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\soc_inst.cpu_core.id_rs2_data[21] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\soc_inst.cpu_core.id_rs2_data[16] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_00271_),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_01070_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\soc_inst.cpu_core.register_file.registers[14][2] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\soc_inst.cpu_core.register_file.registers[11][18] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\soc_inst.cpu_core.register_file.registers[14][5] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\soc_inst.cpu_core.ex_rs2_data[14] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold1216 (.A(_00896_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\soc_inst.cpu_core.ex_exception_pc[0] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_01266_),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\soc_inst.cpu_core.register_file.registers[3][8] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[6] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold1222 (.A(_02121_),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\soc_inst.cpu_core.ex_branch_target[17] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_01887_),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_00280_),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold1227 (.A(_02006_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_00230_),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\soc_inst.cpu_core.csr_file.mepc[19] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold1230 (.A(_01964_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\soc_inst.cpu_core.register_file.registers[9][11] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold1234 (.A(_05227_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_02081_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\soc_inst.cpu_core.ex_rs1_data[20] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold1237 (.A(_01310_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\soc_inst.cpu_core.register_file.registers[12][13] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\soc_inst.cpu_core.alu.b[17] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\soc_inst.cpu_core.register_file.registers[5][18] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\soc_inst.core_mem_rdata[18] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold1243 (.A(_00641_),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\soc_inst.cpu_core.ex_branch_target[12] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold1245 (.A(_01882_),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\soc_inst.cpu_core.register_file.registers[3][31] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\soc_inst.cpu_core.register_file.registers[8][17] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\soc_inst.cpu_core.register_file.registers[11][16] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\soc_inst.cpu_core.register_file.registers[4][11] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_00258_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold1253 (.A(_00448_),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\soc_inst.cpu_core.csr_file.mscratch[31] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_00754_),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\soc_inst.cpu_core.id_rs2_data[14] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\soc_inst.cpu_core.register_file.registers[1][12] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\soc_inst.cpu_core.register_file.registers[12][14] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\soc_inst.cpu_core.mem_rs1_data[0] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold1265 (.A(_00235_),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\soc_inst.cpu_core.csr_file.mscratch[24] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_00747_),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_00300_),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\soc_inst.cpu_core.register_file.registers[12][5] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\soc_inst.cpu_core.ex_exception_pc[4] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_01270_),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\soc_inst.cpu_core.register_file.registers[12][7] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\soc_inst.cpu_core.register_file.registers[3][5] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\soc_inst.cpu_core.register_file.registers[2][11] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\soc_inst.cpu_core.register_file.registers[10][7] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\soc_inst.cpu_core.register_file.registers[2][6] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_00307_),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_02042_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\soc_inst.cpu_core.register_file.registers[5][16] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_05225_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_02079_),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\soc_inst.cpu_core.register_file.registers[13][5] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\soc_inst.cpu_core.csr_file.mscratch[0] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\soc_inst.cpu_core.register_file.registers[5][29] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\soc_inst.cpu_core.id_rs2_data[12] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\soc_inst.cpu_core.register_file.registers[14][11] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold1298 (.A(_00233_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold1299 (.A(_00423_),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold1302 (.A(_06611_),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold1303 (.A(_00092_),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\soc_inst.cpu_core.csr_file.mscratch[29] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold1305 (.A(_00289_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_02015_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\soc_inst.cpu_core.register_file.registers[5][9] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\soc_inst.cpu_core.alu.b[6] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold1309 (.A(_01204_),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold1311 (.A(_00317_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_02052_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\soc_inst.cpu_core.ex_branch_target[25] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_01895_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold1318 (.A(_00768_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_00250_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[12] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold1322 (.A(_08418_),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\soc_inst.cpu_core.register_file.registers[11][28] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\soc_inst.cpu_core.register_file.registers[12][23] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\soc_inst.cpu_core.register_file.registers[14][19] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\soc_inst.cpu_core.id_rs2_data[2] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\soc_inst.cpu_core.ex_branch_target[28] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\soc_inst.cpu_core.csr_file.mscratch[1] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\soc_inst.cpu_core.csr_file.mtvec[22] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_01948_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\soc_inst.cpu_core.register_file.registers[14][27] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\soc_inst.cpu_core.alu.b[7] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold1334 (.A(_01205_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\soc_inst.cpu_core.register_file.registers[13][19] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\soc_inst.cpu_core.register_file.registers[6][18] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\soc_inst.cpu_core.alu.b[11] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_00288_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_02014_),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\soc_inst.cpu_core.register_file.registers[9][20] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\soc_inst.cpu_core.ex_exception_pc[19] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold1342 (.A(_01285_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_00287_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold1344 (.A(_02013_),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\soc_inst.cpu_core.register_file.registers[3][30] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_00283_),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold1348 (.A(_00265_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_09560_),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\soc_inst.cpu_core.register_file.registers[5][13] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\soc_inst.cpu_core.register_file.registers[6][31] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\soc_inst.cpu_core.csr_file.mtval[8] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold1354 (.A(_01907_),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_00220_),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold1356 (.A(_00393_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\soc_inst.cpu_core.csr_file.mepc[6] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\soc_inst.core_mem_rdata[16] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_00639_),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\soc_inst.cpu_core.ex_exception_pc[23] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold1362 (.A(_01289_),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\soc_inst.core_instr_data[27] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\soc_inst.cpu_core.register_file.registers[14][3] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\soc_inst.cpu_core.register_file.registers[4][14] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\soc_inst.cpu_core.register_file.registers[3][0] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\soc_inst.cpu_core.csr_file.mtval[14] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_01913_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold1371 (.A(_05221_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold1372 (.A(_02077_),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\soc_inst.cpu_core.register_file.registers[9][18] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_sample ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold1377 (.A(_00310_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\soc_inst.cpu_core.if_instr[9] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold1380 (.A(_09568_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\soc_inst.cpu_core.ex_branch_target[30] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_01900_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\soc_inst.cpu_core.ex_branch_target[8] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold1384 (.A(_01878_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold1386 (.A(_00281_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\soc_inst.core_mem_rdata[6] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\soc_inst.core_mem_rdata[28] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold1389 (.A(_00651_),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\soc_inst.cpu_core.csr_file.mscratch[26] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold1391 (.A(_00749_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\soc_inst.spi_inst.rx_shift_reg[19] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\soc_inst.cpu_core.register_file.registers[3][24] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\soc_inst.cpu_core.ex_rs2_data[11] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold1399 (.A(_01365_),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\soc_inst.cpu_core.register_file.registers[9][23] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\soc_inst.cpu_core.register_file.registers[4][25] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_00297_),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\soc_inst.cpu_core.register_file.registers[4][7] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\soc_inst.i2c_inst.bit_cnt[2] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_00242_),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold1408 (.A(_00432_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_00303_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold1410 (.A(_02038_),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\soc_inst.cpu_core.register_file.registers[14][4] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\soc_inst.cpu_core.id_imm[8] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold1413 (.A(_01137_),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold1414 (.A(_00298_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_02033_),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\soc_inst.cpu_core.alu.b[9] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold1418 (.A(_00315_),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold1419 (.A(_02050_),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold1422 (.A(_08420_),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold1423 (.A(_00231_),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\soc_inst.cpu_core.register_file.registers[10][24] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\soc_inst.cpu_core.csr_file.mtval[24] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold1426 (.A(_01923_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\soc_inst.cpu_core.register_file.registers[4][6] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\soc_inst.cpu_core.register_file.registers[8][22] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\soc_inst.cpu_core.ex_exception_pc[20] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold1432 (.A(_01286_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\soc_inst.core_mem_rdata[25] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold1434 (.A(_00648_),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold1437 (.A(_08428_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold1439 (.A(_00285_),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold1440 (.A(_02011_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\soc_inst.cpu_core.register_file.registers[3][16] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\soc_inst.cpu_core.csr_file.mtval[12] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold1443 (.A(_01911_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\soc_inst.cpu_core.register_file.registers[4][22] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\soc_inst.i2c_inst.shift_reg[2] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_00080_),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold1448 (.A(_00759_),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold1450 (.A(_00183_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\soc_inst.cpu_core.ex_instr[18] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\soc_inst.cpu_core.ex_branch_target[31] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold1453 (.A(_01901_),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\soc_inst.cpu_core.csr_file.mtvec[4] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold1456 (.A(_00562_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\soc_inst.cpu_core.register_file.registers[4][1] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\soc_inst.cpu_core.register_file.registers[9][14] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\soc_inst.core_mem_rdata[26] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold1463 (.A(_00649_),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\soc_inst.cpu_core.register_file.registers[4][4] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold1466 (.A(_00237_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\soc_inst.cpu_core.register_file.registers[2][19] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\soc_inst.cpu_core.register_file.registers[3][1] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\soc_inst.cpu_core.register_file.registers[12][12] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold1475 (.A(_07091_),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_00260_),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_00450_),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\soc_inst.i2c_inst.clk_cnt[3] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold1479 (.A(_06477_),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\soc_inst.i2c_inst.start_pending ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\soc_inst.cpu_core.csr_file.mtvec[0] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[25] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold1483 (.A(_00781_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold1485 (.A(_00241_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_00431_),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\soc_inst.cpu_core.register_file.registers[13][28] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\soc_inst.cpu_core.csr_file.mtval[10] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_01909_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\soc_inst.cpu_core.ex_exception_pc[21] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_01287_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\soc_inst.core_mem_rdata[15] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\soc_inst.cpu_core.csr_file.mscratch[28] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold1495 (.A(_00751_),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\soc_inst.core_mem_rdata[31] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold1497 (.A(_00654_),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\soc_inst.cpu_core.register_file.registers[14][15] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\soc_inst.cpu_core.csr_file.mtvec[20] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_01946_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\soc_inst.cpu_core.register_file.registers[10][6] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\soc_inst.cpu_core.id_imm[9] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_01138_),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\soc_inst.cpu_core.register_file.registers[12][16] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[3] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\soc_inst.cpu_core.register_file.registers[14][26] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\soc_inst.cpu_core.if_instr[19] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold1511 (.A(_06596_),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_00099_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\soc_inst.gpio_inst.gpio_out[5] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\soc_inst.cpu_core.id_imm[2] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\soc_inst.cpu_core.register_file.registers[5][3] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\soc_inst.cpu_core.register_file.registers[1][8] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\soc_inst.cpu_core.register_file.registers[13][25] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold1518 (.A(_00313_),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\soc_inst.cpu_core.if_funct7[1] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold1520 (.A(_00232_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\soc_inst.cpu_core.register_file.registers[9][31] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\soc_inst.cpu_core.alu.b[27] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_00254_),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold1526 (.A(_00444_),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\soc_inst.cpu_core.csr_file.mtvec[2] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\soc_inst.cpu_core.id_rs2_data[7] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\soc_inst.cpu_core.id_rs2_data[29] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold1530 (.A(_00305_),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_02040_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\soc_inst.cpu_core.register_file.registers[13][10] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_00173_),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\soc_inst.cpu_core.mem_stall ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold1536 (.A(net4951),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\soc_inst.cpu_core.register_file.registers[13][31] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\soc_inst.cpu_core.register_file.registers[14][31] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_00224_),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold1541 (.A(_00407_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\soc_inst.core_mem_wdata[11] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold1543 (.A(_00279_),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_02005_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\soc_inst.core_mem_rdata[1] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\soc_inst.cpu_core.register_file.registers[5][17] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold1551 (.A(_00758_),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\soc_inst.pwm_inst.channel_duty[0][2] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_00234_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\soc_inst.cpu_core.register_file.registers[5][10] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\soc_inst.cpu_core.csr_file.mepc[20] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold1558 (.A(_07095_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold1561 (.A(_00253_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\soc_inst.core_mem_rdata[17] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold1564 (.A(_00640_),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\soc_inst.cpu_core.register_file.registers[6][20] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_00259_),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold1567 (.A(_00449_),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\soc_inst.cpu_core.ex_exception_pc[22] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold1569 (.A(_01288_),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\soc_inst.cpu_core.id_rs2_data[20] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold1571 (.A(_01374_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\soc_inst.cpu_core.register_file.registers[15][22] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\soc_inst.cpu_core.register_file.registers[2][3] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\soc_inst.cpu_core.register_file.registers[14][6] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_00201_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\soc_inst.cpu_core.register_file.registers[11][10] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold1579 (.A(_00187_),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\soc_inst.cpu_core.ex_exception_pc[17] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_01283_),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_00211_),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\soc_inst.cpu_core.register_file.registers[3][14] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\soc_inst.spi_inst.rx_shift_reg[16] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold1587 (.A(_07103_),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\soc_inst.spi_inst.rx_shift_reg[17] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold1590 (.A(_07104_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\soc_inst.cpu_core.csr_file.mtval[28] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold1592 (.A(_04956_),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold1593 (.A(_00240_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_00430_),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\soc_inst.cpu_core.csr_file.mscratch[25] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\soc_inst.cpu_core.register_file.registers[4][26] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold1598 (.A(_00264_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_09559_),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold1601 (.A(_00782_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\soc_inst.cpu_core.register_file.registers[3][18] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold1605 (.A(_00219_),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold1606 (.A(_00392_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold1608 (.A(_00306_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\soc_inst.cpu_core.ex_instr[5] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\soc_inst.cpu_core.alu.a[7] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_01173_),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\soc_inst.i2c_inst.shift_reg[6] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold1615 (.A(_00084_),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\soc_inst.cpu_core.alu.b[30] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold1617 (.A(_00252_),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_00442_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\soc_inst.cpu_core.register_file.registers[13][26] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold1621 (.A(_02135_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\soc_inst.cpu_core.register_file.registers[9][30] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\soc_inst.i2c_inst.clk_cnt[4] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold1624 (.A(_06479_),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\soc_inst.cpu_core.register_file.registers[11][5] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\soc_inst.cpu_core.register_file.registers[13][23] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\soc_inst.cpu_core.csr_file.mscratch[27] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold1628 (.A(_00750_),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\soc_inst.pwm_inst.channel_duty[1][7] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\soc_inst.spi_inst.bit_counter[2] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold1633 (.A(_07079_),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[0] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\soc_inst.cpu_core.csr_file.mepc[21] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold1636 (.A(_01966_),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_00198_),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\soc_inst.cpu_core.register_file.registers[4][27] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold1640 (.A(_00277_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold1642 (.A(_08422_),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\soc_inst.cpu_core.if_pc[16] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold1644 (.A(_00964_),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold1646 (.A(_08431_),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_00223_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold1648 (.A(_00406_),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\soc_inst.pwm_inst.channel_duty[1][1] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold1651 (.A(_00226_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold1653 (.A(_07089_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\soc_inst.cpu_core.register_file.registers[14][25] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold1656 (.A(_07102_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\soc_inst.cpu_core.register_file.registers[2][5] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold1660 (.A(_01272_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold1661 (.A(_00312_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold1662 (.A(_02047_),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\soc_inst.cpu_core.if_pc[21] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold1664 (.A(_00969_),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold1665 (.A(_00255_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\soc_inst.pwm_inst.channel_duty[1][4] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold1667 (.A(_00249_),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold1668 (.A(_00439_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold1671 (.A(_01271_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold1673 (.A(_08408_),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\soc_inst.cpu_core.mem_stall ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\soc_inst.gpio_inst.gpio_out[0] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold1676 (.A(_00248_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\soc_inst.cpu_core.register_file.registers[11][6] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\soc_inst.pwm_inst.channel_duty[0][1] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_00292_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\soc_inst.cpu_core.register_file.registers[7][30] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold1685 (.A(_07099_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\soc_inst.cpu_core.register_file.registers[4][10] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold1687 (.A(_00243_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold1688 (.A(_00433_),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold1689 (.A(_00286_),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\soc_inst.cpu_core.register_file.registers[8][29] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold1692 (.A(_00762_),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\soc_inst.cpu_core.register_file.registers[3][25] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold1695 (.A(_00189_),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_00760_),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\soc_inst.mem_ctrl.spi_addr[22] ),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold1700 (.A(_00589_),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold1702 (.A(_00783_),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\soc_inst.cpu_core.register_file.registers[11][19] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\soc_inst.cpu_core.register_file.registers[4][16] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\soc_inst.cpu_core.ex_instr[23] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold1707 (.A(_01257_),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_00290_),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold1709 (.A(_02016_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\soc_inst.i2c_inst.data_reg[7] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_00761_),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\soc_inst.cpu_core.register_file.registers[14][18] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\soc_inst.cpu_core.register_file.registers[2][17] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\soc_inst.cpu_core.register_file.registers[3][3] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\soc_inst.core_mem_addr[7] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_01329_),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\soc_inst.cpu_core.register_file.registers[5][0] ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[1] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold1724 (.A(_02072_),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\soc_inst.cpu_core.id_imm[12] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold1726 (.A(_01141_),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\soc_inst.cpu_core.ex_branch_target[0] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\soc_inst.core_mem_addr[11] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold1730 (.A(_01333_),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold1732 (.A(_01087_),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold1735 (.A(_00778_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold1736 (.A(_00301_),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold1737 (.A(_02036_),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\soc_inst.cpu_core.if_pc[13] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold1739 (.A(_00961_),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\soc_inst.cpu_core.ex_branch_target[29] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold1744 (.A(_01899_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\soc_inst.cpu_core.register_file.registers[4][3] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\soc_inst.cpu_core.ex_branch_target[11] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold1748 (.A(_01881_),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\soc_inst.gpio_inst.gpio_out[2] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_00506_),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold1751 (.A(_00236_),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_00426_),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold1753 (.A(_00244_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold1754 (.A(_00434_),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\soc_inst.cpu_core.register_file.registers[1][27] ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\soc_inst.cpu_core.register_file.registers[11][20] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\soc_inst.cpu_core.register_file.registers[8][8] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold1760 (.A(_00282_),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\soc_inst.pwm_inst.channel_duty[0][12] ),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold1763 (.A(_05219_),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\soc_inst.cpu_core.register_file.registers[6][25] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\soc_inst.cpu_core.register_file.registers[1][11] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold1769 (.A(_08426_),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[3] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_08409_),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold1772 (.A(_00257_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\soc_inst.cpu_core.csr_file.mtval[21] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold1774 (.A(_01920_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\soc_inst.gpio_inst.gpio_out[4] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold1778 (.A(_00318_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold1779 (.A(_02053_),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\soc_inst.cpu_core.alu.b[24] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold1782 (.A(_08423_),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold1783 (.A(_00302_),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\soc_inst.cpu_core.register_file.registers[4][18] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\soc_inst.cpu_core.register_file.registers[12][15] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold1788 (.A(_00247_),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\soc_inst.pwm_inst.channel_duty[1][6] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold1790 (.A(_00339_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold1791 (.A(_00221_),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\soc_inst.cpu_core.ex_funct3[2] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\soc_inst.cpu_core.if_pc[20] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold1794 (.A(_00968_),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\soc_inst.cpu_core.ex_rs2_data[28] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold1797 (.A(_01382_),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\soc_inst.cpu_core.ex_branch_target[27] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold1799 (.A(_01897_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\soc_inst.core_mem_addr[30] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold1801 (.A(_01352_),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold1803 (.A(_00780_),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\soc_inst.cpu_core.mem_instr[17] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold1805 (.A(_01082_),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\soc_inst.core_mem_rdata[4] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\soc_inst.cpu_core.csr_file.mtvec[21] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold1809 (.A(_01947_),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\soc_inst.cpu_core.ex_branch_target[2] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold1811 (.A(_04344_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_00227_),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\soc_inst.cpu_core.register_file.registers[13][8] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold1815 (.A(_07052_),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold1816 (.A(_00195_),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\soc_inst.cpu_core.alu.b[12] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\soc_inst.cpu_core.alu.b[16] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\soc_inst.cpu_core.if_pc[11] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold1821 (.A(_00959_),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold1823 (.A(_00193_),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\soc_inst.core_mem_addr[6] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold1825 (.A(_01328_),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold1828 (.A(_00757_),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold1830 (.A(_00567_),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\soc_inst.gpio_inst.gpio_out[3] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\soc_inst.cpu_core.ex_is_ebreak ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold1834 (.A(_09247_),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\soc_inst.cpu_core.csr_file.mepc[14] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\soc_inst.cpu_core.id_imm[1] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold1838 (.A(_01130_),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold1839 (.A(_00278_),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\soc_inst.spi_inst.clk_counter[3] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold1841 (.A(_00127_),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold1843 (.A(_07098_),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\soc_inst.cpu_core.alu.a[6] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold1845 (.A(_01172_),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold1847 (.A(_00316_),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold1848 (.A(_02051_),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[0] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold1850 (.A(_08406_),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold1852 (.A(_08412_),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\soc_inst.cpu_core.csr_file.mtval[31] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold1856 (.A(_04973_),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\soc_inst.spi_inst.clk_counter[4] ),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold1858 (.A(_00128_),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\soc_inst.cpu_core.csr_file.mstatus[29] ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold1860 (.A(_02112_),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\soc_inst.pwm_inst.channel_duty[1][2] ),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\soc_inst.cpu_core.csr_file.mtval[23] ),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold1863 (.A(_01922_),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold1864 (.A(_00246_),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\soc_inst.gpio_bidir_out [0]),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\soc_inst.cpu_core.register_file.registers[3][23] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\soc_inst.cpu_core.if_pc[15] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold1869 (.A(_00963_),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\soc_inst.cpu_core.csr_file.mepc[23] ),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold1873 (.A(_00763_),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold1874 (.A(_00225_),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold1875 (.A(_00408_),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[1] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold1877 (.A(_08407_),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\soc_inst.cpu_core.ex_exception_pc[16] ),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold1880 (.A(_01282_),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\soc_inst.cpu_core.id_imm[3] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\soc_inst.cpu_core.alu.b[10] ),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold1883 (.A(_01208_),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[3] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold1885 (.A(_02025_),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold1886 (.A(_00284_),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\soc_inst.cpu_core.register_file.registers[6][19] ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\soc_inst.pwm_inst.channel_duty[1][5] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\soc_inst.core_mem_wdata[8] ),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\soc_inst.gpio_inst.int_en_reg[4] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold1892 (.A(_00261_),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\soc_inst.cpu_core.ex_rs2_data[23] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold1895 (.A(_01377_),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\soc_inst.cpu_core.ex_alu_result[23] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\soc_inst.cpu_core.if_pc[14] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold1898 (.A(_00962_),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold1900 (.A(_07101_),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[2] ),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold1902 (.A(_02024_),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\soc_inst.cpu_core.id_instr[9] ),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold1904 (.A(_01243_),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\soc_inst.spi_inst.bit_counter[3] ),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold1906 (.A(_07080_),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold1907 (.A(_00353_),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\soc_inst.cpu_core.if_funct3[0] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold1909 (.A(_09571_),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\soc_inst.cpu_core.if_pc[12] ),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold1911 (.A(_00960_),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold1914 (.A(_02120_),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\soc_inst.spi_inst.clk_counter[6] ),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold1916 (.A(_06406_),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold1917 (.A(_00130_),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\soc_inst.cpu_core.ex_alu_result[17] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\soc_inst.cpu_core.register_file.registers[8][3] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\soc_inst.gpio_bidir_oe [0]),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold1923 (.A(_00876_),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\soc_inst.cpu_core.csr_file.mstatus[17] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold1925 (.A(_02100_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\soc_inst.cpu_core.if_pc[22] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold1929 (.A(_00970_),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold1930 (.A(_00308_),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold1931 (.A(_02043_),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\soc_inst.cpu_core.register_file.registers[4][17] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\soc_inst.cpu_core.csr_file.mstatus[2] ),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\soc_inst.cpu_core.csr_file.mstatus[19] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold1935 (.A(_02102_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\soc_inst.cpu_core.ex_instr[2] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold1937 (.A(_01236_),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\soc_inst.cpu_core.register_file.registers[1][7] ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\soc_inst.core_mem_addr[5] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold1940 (.A(_01327_),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\soc_inst.cpu_core.id_imm[4] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold1942 (.A(_01133_),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\soc_inst.cpu_core.register_file.registers[3][11] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\soc_inst.cpu_core.csr_file.mtval[18] ),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold1945 (.A(_01917_),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold1946 (.A(_00256_),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold1947 (.A(_00446_),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\soc_inst.cpu_core.if_pc[19] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold1949 (.A(_00967_),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\soc_inst.cpu_core.alu.b[25] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\soc_inst.cpu_core.if_is_compressed ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\soc_inst.cpu_core.if_pc[8] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold1953 (.A(_00956_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\soc_inst.cpu_core.if_pc[10] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold1955 (.A(_00958_),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\soc_inst.cpu_core.if_pc[3] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold1957 (.A(_00951_),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\soc_inst.cpu_core.id_imm[7] ),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold1959 (.A(_01136_),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\soc_inst.cpu_core.csr_file.mtval[15] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold1961 (.A(_01914_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\soc_inst.cpu_core.ex_instr[20] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold1964 (.A(_01254_),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\soc_inst.cpu_core.mem_instr[18] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\soc_inst.cpu_core.register_file.registers[13][4] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold1968 (.A(_01096_),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\soc_inst.cpu_core.csr_file.mstatus[14] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold1970 (.A(_02097_),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold1972 (.A(_00192_),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold1974 (.A(_01276_),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\soc_inst.cpu_core.register_file.registers[6][26] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\soc_inst.i2c_inst.data_reg[3] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold1977 (.A(_06993_),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\soc_inst.cpu_core.csr_file.mstatus[25] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold1980 (.A(_02108_),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold1982 (.A(_02073_),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\soc_inst.cpu_core.csr_file.mepc[16] ),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\soc_inst.cpu_core.ex_branch_target[19] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\soc_inst.cpu_core.csr_file.mstatus[27] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold1986 (.A(_02110_),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold1987 (.A(_00222_),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\soc_inst.cpu_core.ex_instr[11] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\soc_inst.cpu_core.ex_funct7[1] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold1990 (.A(_01091_),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\soc_inst.cpu_core.register_file.registers[8][1] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\soc_inst.cpu_core.csr_file.mstatus[18] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold1993 (.A(_02101_),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\soc_inst.mem_ctrl.spi_data_out[26] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold1995 (.A(_00872_),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold1996 (.A(_00294_),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold1997 (.A(_02021_),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\soc_inst.cpu_core.csr_file.mtval[22] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\soc_inst.cpu_core.if_funct7[3] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\soc_inst.cpu_core.ex_funct7[2] ),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold2001 (.A(_01261_),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold2003 (.A(_00462_),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\soc_inst.cpu_core.ex_funct7[3] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold2005 (.A(_01262_),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\soc_inst.cpu_core.csr_file.mstatus[7] ),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold2007 (.A(_02019_),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\soc_inst.cpu_core.ex_instr[10] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold2010 (.A(_00218_),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\soc_inst.cpu_core.id_imm[18] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold2012 (.A(_01147_),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\soc_inst.cpu_core.id_imm[6] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\soc_inst.cpu_core.ex_rs1_data[30] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold2015 (.A(_01320_),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold2017 (.A(_00466_),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\soc_inst.core_instr_data[25] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\soc_inst.mem_ctrl.spi_data_out[31] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold2020 (.A(_00877_),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\soc_inst.cpu_core.csr_file.mstatus[16] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold2022 (.A(_02099_),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\soc_inst.gpio_inst.int_en_reg[2] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold2024 (.A(_00512_),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold2026 (.A(_02091_),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\soc_inst.cpu_core.ex_instr[7] ),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold2028 (.A(_01230_),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\soc_inst.cpu_core.ex_rs1_data[12] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold2030 (.A(_01302_),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\soc_inst.cpu_core.csr_file.mstatus[26] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold2032 (.A(_02109_),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\soc_inst.cpu_core.register_file.registers[2][23] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold2035 (.A(_05358_),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold2036 (.A(_05361_),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\soc_inst.cpu_core.csr_file.mepc[17] ),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold2038 (.A(_00291_),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold2039 (.A(_02017_),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\soc_inst.pwm_inst.channel_duty[1][0] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold2041 (.A(_00239_),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\soc_inst.cpu_core.csr_file.mstatus[23] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold2043 (.A(_02106_),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\soc_inst.cpu_core.if_funct7[5] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold2047 (.A(_06114_),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold2049 (.A(_00178_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold2051 (.A(_00238_),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\soc_inst.cpu_core.mem_instr[16] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold2053 (.A(_01081_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold2055 (.A(_05365_),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold2056 (.A(_02142_),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\soc_inst.cpu_core.if_pc[1] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold2058 (.A(_00949_),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\soc_inst.i2c_inst.prescale_reg[6] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold2060 (.A(_00411_),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\soc_inst.cpu_core.id_imm12[6] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold2063 (.A(_07094_),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold2065 (.A(_05229_),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\soc_inst.cpu_core.alu.b[15] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\soc_inst.i2c_inst.data_reg[1] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold2069 (.A(_06988_),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold2070 (.A(_02149_),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\soc_inst.i2c_inst.ack_enable ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\soc_inst.gpio_inst.int_en_reg[0] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\soc_inst.cpu_core.id_instr[16] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold2074 (.A(_01250_),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\soc_inst.core_mem_addr[26] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold2076 (.A(_01348_),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\soc_inst.i2c_inst.data_reg[5] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold2078 (.A(_06997_),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold2079 (.A(_02153_),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\soc_inst.cpu_core.id_is_compressed ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\soc_inst.cpu_core.ex_rs2_data[13] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold2085 (.A(_00895_),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\soc_inst.cpu_core.if_pc[23] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold2087 (.A(_00971_),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\soc_inst.cpu_core.id_imm[10] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold2090 (.A(_05231_),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\soc_inst.gpio_inst.int_en_reg[5] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold2092 (.A(_00266_),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold2093 (.A(_09563_),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\soc_inst.cpu_core.id_imm[17] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold2095 (.A(\soc_inst.core_instr_addr[0] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold2096 (.A(_00794_),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\soc_inst.i2c_inst.state[0] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold2098 (.A(_00563_),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\soc_inst.i2c_inst.clk_cnt[5] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\soc_inst.gpio_inst.int_en_reg[1] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\soc_inst.pwm_inst.channel_duty[1][12] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold2103 (.A(_05355_),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold2104 (.A(_02137_),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\soc_inst.cpu_core.id_instr[8] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold2106 (.A(_01242_),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\soc_inst.cpu_core.ex_exception_pc[1] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold2108 (.A(_01267_),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\soc_inst.cpu_core.mem_instr[6] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold2110 (.A(_01075_),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\soc_inst.cpu_core.id_imm[16] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold2112 (.A(_01145_),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold2115 (.A(_07029_),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\soc_inst.core_mem_wdata[10] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\soc_inst.core_mem_addr[10] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold2118 (.A(_01332_),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\soc_inst.pwm_inst.channel_duty[1][15] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\soc_inst.cpu_core.if_pc[0] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\soc_inst.pwm_inst.channel_duty[1][11] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold2125 (.A(_00263_),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold2126 (.A(_05951_),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold2127 (.A(_00331_),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\soc_inst.core_instr_data[13] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\soc_inst.cpu_core.ex_branch_target[9] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold2131 (.A(_01879_),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\soc_inst.pwm_inst.channel_duty[1][8] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\soc_inst.gpio_inst.int_en_reg[6] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\soc_inst.cpu_core.csr_file.mstatus[20] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\soc_inst.cpu_core.ex_alu_result[22] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold2138 (.A(_06044_),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold2141 (.A(_07044_),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold2142 (.A(_00186_),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold2143 (.A(_00319_),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\soc_inst.cpu_core.if_funct3[2] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\soc_inst.cpu_core.ex_rs1_data[17] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold2146 (.A(_00990_),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\soc_inst.cpu_core.ex_branch_target[20] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_01890_),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold2150 (.A(_00185_),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\soc_inst.cpu_core.if_pc[7] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold2152 (.A(_00955_),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\soc_inst.cpu_core.csr_file.mstatus[22] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold2154 (.A(_02105_),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\soc_inst.cpu_core.csr_file.mstatus[31] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold2156 (.A(_02114_),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\soc_inst.cpu_core.id_rs2_data[22] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold2158 (.A(_01376_),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\soc_inst.spi_inst.clock_divider[7] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\soc_inst.cpu_core.id_imm[5] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold2161 (.A(_01134_),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold2163 (.A(_02023_),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\soc_inst.pwm_inst.channel_counter[1][3] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold2165 (.A(_06533_),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\soc_inst.cpu_core.alu.a[25] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\soc_inst.cpu_core.ex_exception_pc[3] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold2168 (.A(_01269_),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\soc_inst.cpu_core.csr_file.mcause[31] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold2170 (.A(_05099_),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold2171 (.A(_01969_),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\soc_inst.cpu_core.if_funct7[0] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\soc_inst.cpu_core.ex_funct3[1] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\soc_inst.core_mem_addr[31] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold2177 (.A(_01353_),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\soc_inst.cpu_core.id_rs2_data[0] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\soc_inst.cpu_core.id_rs2_data[13] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold2180 (.A(\soc_inst.cpu_core.csr_file.mret_trigger ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\soc_inst.core_mem_addr[28] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold2182 (.A(_01350_),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\soc_inst.cpu_core.ex_funct7[1] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\soc_inst.pwm_inst.channel_duty[0][4] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\soc_inst.cpu_core.ex_branch_target[10] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\soc_inst.cpu_core.ex_rs1_data[26] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold2187 (.A(_01316_),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\soc_inst.core_mem_addr[24] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold2190 (.A(_01346_),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\soc_inst.cpu_core.ex_funct7[6] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold2192 (.A(_01265_),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\soc_inst.pwm_inst.channel_counter[1][10] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold2194 (.A(_06546_),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold2195 (.A(_00108_),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\soc_inst.i2c_inst.clk_cnt[6] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\soc_inst.cpu_core.id_rs2_data[4] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\soc_inst.cpu_core.if_funct3[1] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\soc_inst.spi_inst.spi_sclk ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold2200 (.A(_06408_),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold2201 (.A(_00132_),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\soc_inst.cpu_core.id_imm[14] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold2203 (.A(_00268_),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold2204 (.A(_01235_),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\soc_inst.cpu_core.alu.b[31] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold2206 (.A(_01229_),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\soc_inst.cpu_core.if_pc[9] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold2208 (.A(_00957_),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\soc_inst.cpu_core.if_pc[5] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold2210 (.A(_00953_),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold2211 (.A(_00267_),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold2212 (.A(_01234_),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\soc_inst.cpu_core.ex_alu_result[31] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\soc_inst.pwm_inst.channel_duty[1][3] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold2216 (.A(_00465_),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold2218 (.A(_06602_),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold2219 (.A(_00102_),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\soc_inst.spi_inst.state[0] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\soc_inst.cpu_core.id_rs2_data[5] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\soc_inst.pwm_inst.channel_counter[1][13] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold2223 (.A(_06553_),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold2224 (.A(_00111_),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\soc_inst.spi_inst.clock_divider[6] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold2226 (.A(_00320_),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold2227 (.A(_02055_),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\soc_inst.cpu_core.csr_file.mcause[0] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\soc_inst.cpu_core.id_imm12[8] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\soc_inst.i2c_inst.data_reg[4] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold2231 (.A(_06995_),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold2232 (.A(_02152_),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold2233 (.A(_00324_),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold2234 (.A(_02059_),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\soc_inst.pwm_inst.channel_duty[1][13] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold2236 (.A(_00346_),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\soc_inst.cpu_core.if_pc[6] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold2238 (.A(_00954_),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold2240 (.A(_06605_),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold2241 (.A(_00103_),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\soc_inst.spi_inst.bit_counter[0] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\soc_inst.pwm_inst.channel_counter[1][4] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold2245 (.A(_00458_),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\soc_inst.cpu_core.if_funct7[4] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\soc_inst.mem_ctrl.spi_addr[10] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold2249 (.A(_00577_),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\soc_inst.cpu_core.csr_file.mstatus[21] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\soc_inst.cpu_core.id_imm12[2] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold2253 (.A(_01256_),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\soc_inst.cpu_core.id_imm[15] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\soc_inst.cpu_core.alu.a[5] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\soc_inst.cpu_core.csr_file.mstatus[0] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\soc_inst.mem_ctrl.spi_addr[5] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold2258 (.A(_00572_),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold2260 (.A(_07088_),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\soc_inst.cpu_core.register_file.registers[2][30] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold2263 (.A(_00269_),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold2264 (.A(_01238_),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\soc_inst.cpu_core.if_pc[18] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold2266 (.A(_00966_),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\soc_inst.cpu_core.alu.a[0] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\soc_inst.core_mem_addr[25] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold2269 (.A(_01347_),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold2270 (.A(\soc_inst.cpu_core.csr_file.mtval[25] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\soc_inst.cpu_core.alu.op[1] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\soc_inst.cpu_core.ex_branch_target[21] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold2273 (.A(_01891_),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\soc_inst.cpu_core.ex_branch_target[13] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\soc_inst.cpu_core.id_imm12[4] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold2277 (.A(_09583_),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\soc_inst.pwm_inst.channel_counter[1][1] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\soc_inst.i2c_inst.prescale_reg[5] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\soc_inst.cpu_core.id_imm12[7] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold2281 (.A(_09586_),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold2282 (.A(\soc_inst.cpu_core.id_imm[30] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold2283 (.A(_02463_),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\soc_inst.cpu_core.ex_instr[24] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold2285 (.A(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\soc_inst.cpu_core.if_instr[16] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\soc_inst.cpu_core.if_pc[17] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold2291 (.A(_00965_),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\soc_inst.cpu_core.csr_file.mstatus[15] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\soc_inst.core_mem_addr[9] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold2294 (.A(_01331_),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold2296 (.A(_00832_),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\soc_inst.spi_inst.bit_counter[4] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\soc_inst.cpu_core.id_rs2_data[8] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\soc_inst.spi_inst.clk_counter[5] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold2301 (.A(_00129_),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\soc_inst.cpu_core.alu.a[8] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold2304 (.A(_00293_),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold2305 (.A(_02020_),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\soc_inst.cpu_core.ex_branch_target[3] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\soc_inst.cpu_core.register_file.registers[1][30] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold2310 (.A(_00576_),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\soc_inst.cpu_core.alu.b[22] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\soc_inst.pwm_inst.channel_counter[1][8] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold2313 (.A(_06543_),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\soc_inst.pwm_inst.channel_counter[1][12] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold2315 (.A(_06550_),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold2316 (.A(_00110_),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\soc_inst.cpu_core.csr_file.mstatus[1] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\soc_inst.cpu_core.alu.a[1] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\soc_inst.cpu_core.ex_rs2_data[26] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\soc_inst.cpu_core.csr_file.mtval[27] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold2321 (.A(_04949_),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold2322 (.A(_01926_),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\soc_inst.cpu_core.csr_file.mstatus[4] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\soc_inst.cpu_core.if_pc[4] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold2325 (.A(_00952_),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\soc_inst.i2c_inst.restart_pending ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[0] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold2328 (.A(_02022_),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\soc_inst.pwm_inst.channel_duty[1][14] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold2330 (.A(_00347_),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\soc_inst.gpio_inst.int_en_reg[3] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\soc_inst.cpu_core.csr_file.mstatus[30] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold2333 (.A(_02113_),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\soc_inst.core_mem_addr[27] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold2335 (.A(_01349_),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\soc_inst.cpu_core.csr_file.mstatus[13] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\soc_inst.pwm_inst.channel_duty[1][9] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\soc_inst.core_mem_rdata[24] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\soc_inst.cpu_core.alu.a[9] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\soc_inst.cpu_core.csr_file.mtval[29] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold2342 (.A(_00181_),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\soc_inst.mem_ctrl.spi_addr[14] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold2344 (.A(_00581_),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\soc_inst.cpu_core.alu.op[2] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold2347 (.A(_00176_),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\soc_inst.cpu_core.ex_alu_result[10] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\soc_inst.mem_ctrl.spi_addr[23] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold2350 (.A(_00590_),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\soc_inst.cpu_core.alu.b[28] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold2354 (.A(_06614_),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\soc_inst.core_mem_addr[22] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\soc_inst.cpu_core.if_imm12[2] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\soc_inst.cpu_core.id_rs2_data[23] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\soc_inst.cpu_core.csr_file.mstatus[28] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold2359 (.A(_02111_),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold2361 (.A(_00177_),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\soc_inst.cpu_core.register_file.registers[12][31] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\soc_inst.cpu_core.ex_branch_target[1] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\soc_inst.cpu_core.ex_instr[3] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold2365 (.A(_01237_),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\soc_inst.cpu_core.id_rs2_data[17] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold2367 (.A(_01371_),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold2368 (.A(\soc_inst.pwm_inst.channel_counter[1][6] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold2369 (.A(_06540_),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold2370 (.A(_00119_),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\soc_inst.cpu_core.csr_file.mcause[1] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold2373 (.A(_00038_),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\soc_inst.cpu_core.csr_file.mcause[2] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\soc_inst.cpu_core.alu.a[31] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\soc_inst.cpu_core.alu.a[26] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\soc_inst.cpu_core.alu.a[3] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\soc_inst.cpu_core.ex_rs1_data[10] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold2379 (.A(_00983_),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\soc_inst.mem_ctrl.spi_addr[17] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold2381 (.A(_00584_),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold2382 (.A(\soc_inst.core_instr_data[12] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\soc_inst.i2c_inst.clk_cnt[1] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold2385 (.A(_09188_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold2386 (.A(_00875_),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\soc_inst.cpu_core.alu.a[14] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold2388 (.A(\soc_inst.cpu_core.ex_rs2_data[30] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\soc_inst.pwm_inst.channel_counter[1][11] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold2390 (.A(_06549_),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\soc_inst.pwm_ena[1] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\soc_inst.cpu_core.alu.b[23] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold2394 (.A(_06601_),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold2395 (.A(_00101_),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\soc_inst.cpu_core.alu.b[8] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\soc_inst.cpu_core.csr_file.mtval[3] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\soc_inst.cpu_core.ex_alu_result[27] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\soc_inst.spi_inst.clock_divider[5] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold2400 (.A(\soc_inst.cpu_core.csr_file.mtval[1] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold2401 (.A(_00065_),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\soc_inst.cpu_core.alu.b[18] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold2403 (.A(\soc_inst.pwm_inst.channel_counter[1][5] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\soc_inst.spi_inst.len_sel[0] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold2405 (.A(_00468_),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\soc_inst.cpu_core.csr_file.mepc[11] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold2407 (.A(_01956_),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold2409 (.A(_00588_),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\soc_inst.pwm_ena[0] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\soc_inst.core_mem_addr[14] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold2412 (.A(_01336_),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold2413 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold2415 (.A(\soc_inst.cpu_core.id_imm[13] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\soc_inst.mem_ctrl.spi_addr[8] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold2417 (.A(_00575_),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold2418 (.A(\soc_inst.core_instr_addr[3] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold2419 (.A(_00797_),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\soc_inst.cpu_core.id_funct3[1] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\soc_inst.core_instr_data[0] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\soc_inst.cpu_core.id_rs2_data[24] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold2424 (.A(\soc_inst.core_mem_rdata[0] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\soc_inst.mem_ctrl.spi_addr[4] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold2426 (.A(_00571_),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold2427 (.A(\soc_inst.cpu_core.id_imm12[11] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold2428 (.A(_09591_),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold2430 (.A(_00582_),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\soc_inst.mem_ctrl.spi_is_instr ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold2432 (.A(_00004_),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\soc_inst.mem_ctrl.spi_addr[7] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold2434 (.A(_00574_),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\soc_inst.mem_ctrl.spi_addr[20] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold2436 (.A(_00587_),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\soc_inst.core_mem_addr[16] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold2438 (.A(\soc_inst.cpu_core.ex_branch_target[7] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\soc_inst.cpu_core.id_imm[0] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold2440 (.A(\soc_inst.cpu_core.alu.a[4] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\soc_inst.cpu_core.alu.a[11] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold2442 (.A(\soc_inst.cpu_core.ex_branch_target[18] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold2443 (.A(_00217_),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold2444 (.A(\soc_inst.mem_ctrl.spi_addr[19] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold2445 (.A(_00586_),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold2446 (.A(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold2447 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold2448 (.A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold2449 (.A(_00580_),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[6] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold2451 (.A(_05169_),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold2452 (.A(_05171_),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\soc_inst.cpu_core.csr_file.mcause[3] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold2454 (.A(_00051_),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold2455 (.A(\soc_inst.core_instr_addr[1] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold2456 (.A(_00795_),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\soc_inst.cpu_core.ex_instr[21] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold2458 (.A(_01255_),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\soc_inst.core_instr_addr[4] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold2460 (.A(_00798_),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold2461 (.A(\soc_inst.spi_inst.bit_counter[5] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold2463 (.A(_07041_),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold2464 (.A(_00184_),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold2465 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold2466 (.A(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold2467 (.A(_06618_),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold2468 (.A(\soc_inst.cpu_core.csr_file.mtval[30] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold2469 (.A(_01929_),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold2470 (.A(\soc_inst.core_mem_addr[20] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold2471 (.A(\soc_inst.pwm_inst.channel_counter[1][14] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\soc_inst.cpu_core.id_rs1_data[10] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold2473 (.A(\soc_inst.cpu_core.id_rs1_data[14] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold2474 (.A(\soc_inst.core_instr_data[2] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold2475 (.A(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold2476 (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold2477 (.A(\soc_inst.cpu_core.id_rs2_data[28] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\soc_inst.cpu_core.csr_file.mtval[2] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold2479 (.A(\soc_inst.cpu_core.ex_instr[9] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold2480 (.A(_01232_),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold2481 (.A(\soc_inst.cpu_core.csr_file.mepc[12] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\soc_inst.cpu_core.id_pc[23] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold2484 (.A(_00573_),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold2485 (.A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\soc_inst.mem_ctrl.spi_data_out[21] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold2487 (.A(\soc_inst.mem_ctrl.spi_data_out[22] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\soc_inst.mem_ctrl.access_state[3] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold2489 (.A(_00008_),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold2490 (.A(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold2491 (.A(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold2492 (.A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold2493 (.A(_00579_),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold2495 (.A(_00570_),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\soc_inst.mem_ctrl.spi_addr[11] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold2497 (.A(_00578_),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\soc_inst.cpu_core.id_rs2_data[10] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold2500 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold2501 (.A(_00000_),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold2502 (.A(\soc_inst.cpu_core.if_instr[2] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold2503 (.A(_09561_),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold2504 (.A(\soc_inst.cpu_core.id_pc[4] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\soc_inst.core_mem_addr[8] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold2506 (.A(_01330_),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\soc_inst.cpu_core.id_imm12[3] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold2508 (.A(_09582_),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold2509 (.A(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold2510 (.A(_00196_),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold2511 (.A(\soc_inst.cpu_core.ex_rs1_data[9] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold2512 (.A(_01299_),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold2513 (.A(\soc_inst.cpu_core.alu.b[21] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold2514 (.A(\soc_inst.gpio_inst.gpio_out[1] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold2515 (.A(_00505_),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold2516 (.A(\soc_inst.cpu_core.csr_file.mtval[26] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold2517 (.A(_04943_),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold2518 (.A(_01925_),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold2519 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[3] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold2520 (.A(_05350_),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold2521 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\soc_inst.cpu_core.alu.a[16] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold2524 (.A(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\soc_inst.core_instr_data[14] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\soc_inst.i2c_inst.clk_cnt[7] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\soc_inst.cpu_core.id_imm[29] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold2528 (.A(_02459_),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold2529 (.A(\soc_inst.core_instr_addr[13] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold2530 (.A(\soc_inst.cpu_core.if_instr[5] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold2531 (.A(\soc_inst.cpu_core.ex_funct3[0] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold2532 (.A(_01246_),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold2533 (.A(\soc_inst.mem_ctrl.spi_data_out[17] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold2534 (.A(\soc_inst.cpu_core.id_rs2_data[27] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold2535 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\soc_inst.pwm_inst.channel_counter[1][9] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold2538 (.A(_00874_),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold2539 (.A(\soc_inst.cpu_core.alu.b[19] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold2540 (.A(_01217_),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\soc_inst.cpu_core.ex_alu_result[24] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold2542 (.A(uio_out[4]),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\soc_inst.cpu_core.alu.b[13] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold2544 (.A(\soc_inst.cpu_core.id_pc[8] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\soc_inst.cpu_core.id_imm[25] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold2546 (.A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold2547 (.A(_00585_),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold2548 (.A(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold2549 (.A(\soc_inst.cpu_core.alu.b[20] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold2550 (.A(\soc_inst.cpu_core.id_pc[19] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\soc_inst.core_instr_addr[5] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold2552 (.A(\soc_inst.spi_inst.cpol ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold2553 (.A(\soc_inst.cpu_core.id_imm12[1] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold2554 (.A(_09580_),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\soc_inst.cpu_core.ex_rs1_data[31] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold2556 (.A(_01321_),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold2558 (.A(\soc_inst.cpu_core.id_rs2_data[15] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold2559 (.A(_01112_),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold2560 (.A(\soc_inst.core_mem_flag[0] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold2561 (.A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold2563 (.A(\soc_inst.mem_ctrl.spi_data_out[25] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold2564 (.A(_00871_),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold2565 (.A(\soc_inst.cpu_core.ex_alu_result[21] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold2566 (.A(\soc_inst.pwm_inst.channel_counter[1][7] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold2567 (.A(\soc_inst.i2c_inst.data_reg[6] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold2570 (.A(\soc_inst.cpu_core.ex_alu_result[26] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\soc_inst.cpu_core.ex_alu_result[13] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold2572 (.A(\soc_inst.cpu_core.id_imm[27] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold2573 (.A(_02451_),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold2574 (.A(_00327_),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold2575 (.A(_02087_),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold2576 (.A(_00329_),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold2577 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold2578 (.A(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold2579 (.A(_00857_),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold2581 (.A(\soc_inst.cpu_core.id_pc[10] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\soc_inst.cpu_core.id_pc[11] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold2583 (.A(\soc_inst.i2c_inst.start_pending ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\soc_inst.i2c_inst.state[1] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold2585 (.A(_00564_),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold2586 (.A(\soc_inst.cpu_core.csr_file.mepc[0] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold2587 (.A(_00058_),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold2588 (.A(\soc_inst.mem_ctrl.spi_data_out[23] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold2589 (.A(_00869_),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold2590 (.A(\soc_inst.cpu_core.id_pc[14] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold2591 (.A(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold2592 (.A(_00856_),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\soc_inst.cpu_core.id_pc[18] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold2594 (.A(\soc_inst.core_mem_addr[18] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold2595 (.A(\soc_inst.cpu_core.ex_alu_result[15] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\soc_inst.cpu_core.csr_file.mtval[0] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold2597 (.A(_00064_),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold2598 (.A(\soc_inst.cpu_core.if_imm12[0] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\soc_inst.mem_ctrl.spi_data_out[16] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold2600 (.A(_00862_),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold2601 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold2602 (.A(\soc_inst.cpu_core.ex_instr[8] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold2603 (.A(_01231_),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold2604 (.A(\soc_inst.spi_inst.cpha ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold2605 (.A(\soc_inst.cpu_core.csr_file.mepc[7] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold2606 (.A(_01952_),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold2607 (.A(\soc_inst.mem_ctrl.spi_addr[16] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold2608 (.A(_00583_),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold2609 (.A(\soc_inst.spi_ena ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\soc_inst.cpu_core.alu.a[21] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold2611 (.A(\soc_inst.cpu_core.id_pc[12] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold2613 (.A(_00569_),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold2614 (.A(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold2616 (.A(_00861_),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold2618 (.A(\soc_inst.cpu_core.csr_file.mtval[4] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold2619 (.A(_00068_),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold2620 (.A(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold2622 (.A(_00568_),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold2623 (.A(\soc_inst.cpu_core.id_imm[28] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold2624 (.A(\soc_inst.cpu_core.id_imm12[0] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\soc_inst.cpu_core.id_imm[23] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold2626 (.A(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold2627 (.A(\soc_inst.core_instr_data[10] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold2628 (.A(uio_out[1]),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\soc_inst.core_instr_addr[8] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold2630 (.A(\soc_inst.cpu_core.id_imm[22] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold2631 (.A(\soc_inst.cpu_core.ex_instr[6] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold2632 (.A(_01240_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold2633 (.A(\soc_inst.cpu_core.alu.a[17] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold2634 (.A(\soc_inst.i2c_inst.data_reg[2] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\soc_inst.cpu_core.id_imm[26] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold2636 (.A(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold2637 (.A(_00853_),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold2639 (.A(\soc_inst.cpu_core.if_imm12[4] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\soc_inst.cpu_core.alu.b[26] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold2641 (.A(\soc_inst.cpu_core.alu.a[10] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\soc_inst.cpu_core.if_funct7[6] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold2643 (.A(\soc_inst.cpu_core.csr_file.mepc[2] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold2644 (.A(_00060_),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\soc_inst.mem_ctrl.spi_data_len[5] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold2646 (.A(_00519_),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\soc_inst.core_mem_addr[19] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold2648 (.A(\soc_inst.core_instr_addr[2] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\soc_inst.cpu_core.ex_branch_target[6] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold2651 (.A(_04406_),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold2652 (.A(\soc_inst.core_mem_addr[23] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold2653 (.A(\soc_inst.cpu_core.id_imm[21] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold2654 (.A(_00262_),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold2655 (.A(_08452_),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\soc_inst.cpu_core.id_rs1_data[6] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold2657 (.A(\soc_inst.mem_ctrl.spi_done ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold2658 (.A(_00725_),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold2659 (.A(\soc_inst.core_instr_addr[7] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold2660 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold2661 (.A(_05147_),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold2662 (.A(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold2663 (.A(\soc_inst.mem_ctrl.spi_data_len[4] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold2664 (.A(_00518_),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold2665 (.A(\soc_inst.cpu_core.ex_alu_result[4] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold2666 (.A(_01326_),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold2667 (.A(\soc_inst.cpu_core.alu.op[0] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold2668 (.A(\soc_inst.cpu_core.ex_branch_target[16] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\soc_inst.cpu_core.alu.op[3] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold2670 (.A(\soc_inst.mem_ctrl.access_state[4] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\soc_inst.cpu_core.if_funct7[2] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold2672 (.A(\soc_inst.cpu_core.id_pc[6] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\soc_inst.cpu_core.ex_alu_result[2] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold2674 (.A(_01324_),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold2675 (.A(\soc_inst.cpu_core.id_rs1_data[23] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold2676 (.A(\soc_inst.core_mem_wdata[22] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold2677 (.A(_00904_),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold2678 (.A(\soc_inst.cpu_core.id_rs2_data[30] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold2679 (.A(\soc_inst.cpu_core.id_pc[20] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\soc_inst.core_mem_wdata[23] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold2681 (.A(\soc_inst.mem_ctrl.spi_data_len[3] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold2682 (.A(\soc_inst.core_mem_addr[0] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold2683 (.A(_01322_),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold2684 (.A(\soc_inst.core_instr_addr[14] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold2685 (.A(\soc_inst.cpu_core.id_pc[9] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\soc_inst.cpu_core.mem_reg_we ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold2687 (.A(\soc_inst.cpu_core.id_pc[21] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold2688 (.A(_00328_),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold2689 (.A(_02088_),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\soc_inst.cpu_core.ex_branch_target[22] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold2691 (.A(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold2692 (.A(\soc_inst.core_instr_addr[17] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold2693 (.A(\soc_inst.core_instr_addr[10] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold2694 (.A(\soc_inst.cpu_core.id_pc[17] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\soc_inst.cpu_core.ex_alu_result[11] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold2696 (.A(uio_out[2]),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold2697 (.A(\soc_inst.cpu_core.csr_file.mepc[4] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold2699 (.A(\soc_inst.cpu_core.ex_alu_result[3] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold2700 (.A(_01325_),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold2701 (.A(uio_out[5]),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold2702 (.A(_00791_),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold2703 (.A(\soc_inst.core_instr_addr[9] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\soc_inst.core_instr_addr[6] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold2705 (.A(\soc_inst.cpu_core.if_instr[18] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold2706 (.A(\soc_inst.core_instr_data[3] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold2707 (.A(_00594_),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\soc_inst.cpu_core.id_int_is_interrupt ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold2709 (.A(\soc_inst.cpu_core.id_rs2_data[26] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold2711 (.A(\soc_inst.core_instr_addr[11] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold2712 (.A(\soc_inst.cpu_core.id_pc[15] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold2713 (.A(\soc_inst.core_mem_addr[21] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold2714 (.A(\soc_inst.cpu_core.alu.a[15] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold2715 (.A(\soc_inst.cpu_core.ex_alu_result[28] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold2716 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold2717 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold2718 (.A(_05369_),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold2719 (.A(\soc_inst.cpu_core.id_rs1_data[18] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold2720 (.A(\soc_inst.cpu_core.if_instr[3] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold2721 (.A(_09562_),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold2722 (.A(\soc_inst.cpu_core.id_rs1_data[30] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold2723 (.A(\soc_inst.cpu_core.if_instr[2] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold2724 (.A(\soc_inst.cpu_core.ex_alu_result[9] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold2725 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold2726 (.A(\soc_inst.cpu_core.ex_alu_result[1] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold2727 (.A(\soc_inst.cpu_core.id_pc[5] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\soc_inst.cpu_core.id_pc[13] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold2729 (.A(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold2730 (.A(_00276_),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold2731 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold2732 (.A(\soc_inst.cpu_core.id_pc[2] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold2734 (.A(_00860_),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\soc_inst.core_mem_addr[17] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold2736 (.A(\soc_inst.cpu_core.id_imm[24] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold2737 (.A(\soc_inst.cpu_core.ex_alu_result[14] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold2738 (.A(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold2739 (.A(\soc_inst.cpu_core.ex_alu_result[8] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold2740 (.A(_01394_),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold2741 (.A(\soc_inst.core_instr_data[4] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold2742 (.A(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold2743 (.A(_00852_),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold2744 (.A(\soc_inst.cpu_core.id_rs1_data[9] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold2745 (.A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold2746 (.A(\soc_inst.cpu_core.id_rs1_data[22] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold2747 (.A(\soc_inst.mem_ctrl.access_state[2] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold2748 (.A(\soc_inst.cpu_core.alu.a[22] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold2749 (.A(\soc_inst.core_mem_addr[1] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold2750 (.A(\soc_inst.i2c_inst.data_reg[0] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\soc_inst.cpu_core.id_rs1_data[4] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold2752 (.A(\soc_inst.cpu_core.id_pc[16] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold2753 (.A(\soc_inst.core_instr_addr[23] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold2754 (.A(\soc_inst.core_instr_addr[15] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold2755 (.A(\soc_inst.cpu_core.ex_alu_result[12] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold2756 (.A(_01398_),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold2757 (.A(\soc_inst.cpu_core.id_imm[20] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold2758 (.A(\soc_inst.cpu_core.id_rs2_data[19] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\soc_inst.cpu_core.alu.a[27] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\soc_inst.cpu_core.id_pc[1] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold2761 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold2763 (.A(_09178_),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold2764 (.A(_00873_),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold2765 (.A(\soc_inst.cpu_core.csr_file.mepc[1] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold2766 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\soc_inst.cpu_core.ex_alu_result[0] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\soc_inst.cpu_core.id_rs2_data[11] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold2769 (.A(\soc_inst.core_instr_data[15] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\soc_inst.mem_ctrl.spi_data_out[20] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold2771 (.A(_00866_),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold2772 (.A(\soc_inst.cpu_core.id_rs1_data[8] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold2773 (.A(\soc_inst.cpu_core.ex_rs2_data[20] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold2774 (.A(_00902_),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold2775 (.A(\soc_inst.core_instr_addr[16] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold2776 (.A(\soc_inst.core_instr_addr[22] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold2777 (.A(\soc_inst.core_instr_addr[19] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold2778 (.A(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold2779 (.A(\soc_inst.cpu_core.alu.b[4] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold2780 (.A(uio_oe[5]),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold2781 (.A(_08575_),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold2782 (.A(_00755_),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold2783 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold2784 (.A(\soc_inst.mem_ctrl.spi_mem_inst.is_write_op ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold2785 (.A(_00723_),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold2786 (.A(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold2787 (.A(\soc_inst.cpu_core.id_rs1_data[15] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold2788 (.A(\soc_inst.cpu_core.id_rs1_data[7] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold2789 (.A(\soc_inst.cpu_core.ex_alu_result[7] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold2790 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold2791 (.A(_00830_),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold2792 (.A(\soc_inst.cpu_core.ex_rs2_data[17] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold2793 (.A(_00899_),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold2794 (.A(\soc_inst.cpu_core.id_pc[22] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold2795 (.A(\soc_inst.cpu_core.id_pc[0] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold2796 (.A(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold2797 (.A(\soc_inst.cpu_core.alu.a[2] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold2798 (.A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold2799 (.A(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold2800 (.A(\soc_inst.cpu_core.id_pc[3] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold2801 (.A(\soc_inst.mem_ctrl.spi_data_out[24] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold2802 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold2803 (.A(\soc_inst.mem_ctrl.spi_data_out[19] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold2804 (.A(_00865_),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold2805 (.A(\soc_inst.core_instr_addr[18] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold2806 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold2807 (.A(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold2808 (.A(_07026_),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold2809 (.A(_00216_),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold2810 (.A(\soc_inst.cpu_core.alu.a[24] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\soc_inst.cpu_core.if_imm12[1] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold2812 (.A(\soc_inst.core_instr_data[5] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold2813 (.A(_00596_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold2814 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold2815 (.A(\soc_inst.cpu_core.alu.a[29] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold2816 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold2817 (.A(\soc_inst.cpu_core.alu.a[12] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold2818 (.A(\soc_inst.cpu_core.id_rs1_data[31] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold2819 (.A(\soc_inst.cpu_core.id_rs2_data[9] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold2820 (.A(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold2821 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold2822 (.A(_00829_),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold2823 (.A(\soc_inst.core_instr_addr[20] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold2824 (.A(\soc_inst.cpu_core.csr_file.mepc[3] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold2825 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold2826 (.A(_09164_),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold2827 (.A(\soc_inst.cpu_core.id_rs1_data[3] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold2828 (.A(\soc_inst.core_instr_data[11] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold2829 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold2830 (.A(\soc_inst.cpu_core.ex_alu_result[6] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold2831 (.A(\soc_inst.core_instr_addr[21] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold2832 (.A(\soc_inst.cpu_core.id_pc[7] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold2833 (.A(\soc_inst.cpu_core.alu.b[29] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold2834 (.A(_01227_),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold2835 (.A(\soc_inst.spi_inst.busy ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold2836 (.A(\soc_inst.cpu_core.id_rs1_data[5] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold2837 (.A(\soc_inst.cpu_core.id_rs1_data[13] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold2838 (.A(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold2839 (.A(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold2840 (.A(\soc_inst.cpu_core.id_rs1_data[2] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold2841 (.A(\soc_inst.cpu_core.ex_alu_result[25] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold2842 (.A(\soc_inst.cpu_core.id_rs1_data[0] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold2843 (.A(\soc_inst.cpu_core.id_rs2_data[18] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold2844 (.A(\soc_inst.cpu_core.alu.a[30] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold2845 (.A(\soc_inst.cpu_core.ex_alu_result[5] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold2846 (.A(_01391_),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold2847 (.A(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold2848 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold2849 (.A(_01903_),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold2850 (.A(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold2851 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold2852 (.A(\soc_inst.cpu_core.alu.a[18] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold2853 (.A(\soc_inst.core_instr_addr[12] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold2854 (.A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold2855 (.A(\soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold2856 (.A(\soc_inst.cpu_core.id_rs2_data[31] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold2857 (.A(\soc_inst.core_mem_addr[13] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold2858 (.A(\soc_inst.i2c_inst.state[3] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold2859 (.A(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold2860 (.A(\soc_inst.cpu_core.alu.b[2] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold2861 (.A(\soc_inst.core_mem_we ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold2862 (.A(\soc_inst.cpu_core.ex_alu_result[30] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold2863 (.A(\soc_inst.core_instr_data[6] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold2864 (.A(\soc_inst.cpu_core.id_instr[6] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold2865 (.A(_09565_),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold2866 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold2867 (.A(_06130_),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold2868 (.A(_06150_),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold2869 (.A(_00015_),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold2870 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold2871 (.A(_00831_),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold2872 (.A(\soc_inst.i2c_inst.ctrl_reg[2] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold2873 (.A(\soc_inst.core_mem_addr[15] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold2874 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold2875 (.A(_06128_),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold2876 (.A(_00010_),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold2877 (.A(_00330_),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold2878 (.A(\soc_inst.cpu_core.if_imm12[3] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold2879 (.A(\soc_inst.cpu_core.alu.a[28] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold2880 (.A(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold2881 (.A(_06281_),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold2882 (.A(_00023_),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold2883 (.A(\soc_inst.cpu_core.alu.a[20] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold2884 (.A(\soc_inst.cpu_core.id_rs1_data[29] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold2885 (.A(\soc_inst.spi_inst.len_sel[1] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold2886 (.A(_00469_),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold2887 (.A(\soc_inst.cpu_core.alu.b[1] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold2888 (.A(\soc_inst.cpu_core.alu.a[13] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold2889 (.A(\soc_inst.cpu_core.alu.a[19] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold2890 (.A(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold2891 (.A(_00690_),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold2892 (.A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold2893 (.A(\soc_inst.core_mem_addr[12] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold2894 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold2895 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold2896 (.A(\soc_inst.cpu_core.if_instr[6] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold2897 (.A(\soc_inst.cpu_core.alu.b[0] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold2898 (.A(\soc_inst.cpu_core.if_funct7[4] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold2899 (.A(\soc_inst.cpu_core.if_instr[6] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold2900 (.A(\soc_inst.cpu_core.ex_alu_result[2] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold2901 (.A(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold2902 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold2903 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold2904 (.A(\soc_inst.cpu_core.if_funct3[0] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold2905 (.A(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold2906 (.A(\soc_inst.pwm_ena[0] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold2907 (.A(\soc_inst.cpu_core.id_pc[19] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold2908 (.A(_01889_),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold2909 (.A(\soc_inst.cpu_core.id_pc[3] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold2910 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ),
    .X(net2988));
 sg13g2_antennanp ANTENNA_1 (.A(\soc_inst.mem_ctrl.spi_data_out[27] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_4 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_104 ();
 sg13g2_decap_8 FILLER_0_111 ();
 sg13g2_fill_2 FILLER_0_118 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_fill_1 FILLER_0_131 ();
 sg13g2_decap_4 FILLER_0_145 ();
 sg13g2_fill_1 FILLER_0_149 ();
 sg13g2_decap_4 FILLER_0_163 ();
 sg13g2_fill_2 FILLER_0_167 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_4 FILLER_0_219 ();
 sg13g2_fill_1 FILLER_0_223 ();
 sg13g2_fill_2 FILLER_0_242 ();
 sg13g2_fill_2 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_4 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_fill_2 FILLER_0_285 ();
 sg13g2_decap_4 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_4 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_fill_1 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_4 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_decap_8 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_505 ();
 sg13g2_fill_2 FILLER_0_512 ();
 sg13g2_fill_1 FILLER_0_514 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_fill_1 FILLER_0_547 ();
 sg13g2_decap_4 FILLER_0_569 ();
 sg13g2_fill_2 FILLER_0_576 ();
 sg13g2_fill_1 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_603 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_4 FILLER_0_624 ();
 sg13g2_fill_1 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_632 ();
 sg13g2_fill_2 FILLER_0_639 ();
 sg13g2_fill_1 FILLER_0_641 ();
 sg13g2_decap_8 FILLER_0_647 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_4 FILLER_0_661 ();
 sg13g2_fill_2 FILLER_0_711 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_4 FILLER_0_729 ();
 sg13g2_decap_8 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_fill_2 FILLER_0_778 ();
 sg13g2_fill_1 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_788 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_decap_8 FILLER_0_802 ();
 sg13g2_fill_1 FILLER_0_809 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_fill_2 FILLER_0_896 ();
 sg13g2_fill_1 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_4 FILLER_0_997 ();
 sg13g2_fill_1 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1019 ();
 sg13g2_decap_8 FILLER_0_1026 ();
 sg13g2_decap_8 FILLER_0_1033 ();
 sg13g2_decap_8 FILLER_0_1040 ();
 sg13g2_decap_8 FILLER_0_1047 ();
 sg13g2_decap_8 FILLER_0_1054 ();
 sg13g2_decap_8 FILLER_0_1061 ();
 sg13g2_decap_8 FILLER_0_1068 ();
 sg13g2_decap_8 FILLER_0_1075 ();
 sg13g2_decap_4 FILLER_0_1082 ();
 sg13g2_fill_1 FILLER_0_1086 ();
 sg13g2_fill_2 FILLER_0_1141 ();
 sg13g2_fill_1 FILLER_0_1143 ();
 sg13g2_fill_2 FILLER_0_1162 ();
 sg13g2_fill_1 FILLER_0_1164 ();
 sg13g2_fill_2 FILLER_0_1171 ();
 sg13g2_fill_1 FILLER_0_1173 ();
 sg13g2_fill_2 FILLER_0_1183 ();
 sg13g2_fill_1 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1241 ();
 sg13g2_decap_8 FILLER_0_1248 ();
 sg13g2_fill_2 FILLER_0_1255 ();
 sg13g2_fill_1 FILLER_0_1284 ();
 sg13g2_fill_2 FILLER_0_1291 ();
 sg13g2_fill_1 FILLER_0_1293 ();
 sg13g2_decap_4 FILLER_0_1297 ();
 sg13g2_fill_1 FILLER_0_1310 ();
 sg13g2_decap_8 FILLER_0_1348 ();
 sg13g2_decap_8 FILLER_0_1355 ();
 sg13g2_decap_8 FILLER_0_1362 ();
 sg13g2_fill_2 FILLER_0_1369 ();
 sg13g2_fill_2 FILLER_0_1381 ();
 sg13g2_fill_1 FILLER_0_1425 ();
 sg13g2_decap_8 FILLER_0_1440 ();
 sg13g2_decap_8 FILLER_0_1447 ();
 sg13g2_decap_8 FILLER_0_1454 ();
 sg13g2_fill_1 FILLER_0_1461 ();
 sg13g2_fill_2 FILLER_0_1501 ();
 sg13g2_fill_1 FILLER_0_1503 ();
 sg13g2_fill_1 FILLER_0_1533 ();
 sg13g2_fill_2 FILLER_0_1562 ();
 sg13g2_fill_1 FILLER_0_1574 ();
 sg13g2_fill_1 FILLER_0_1588 ();
 sg13g2_fill_1 FILLER_0_1599 ();
 sg13g2_decap_8 FILLER_0_1637 ();
 sg13g2_fill_1 FILLER_0_1644 ();
 sg13g2_fill_2 FILLER_0_1658 ();
 sg13g2_fill_1 FILLER_0_1660 ();
 sg13g2_decap_8 FILLER_0_1681 ();
 sg13g2_decap_8 FILLER_0_1688 ();
 sg13g2_decap_8 FILLER_0_1695 ();
 sg13g2_decap_8 FILLER_0_1702 ();
 sg13g2_decap_8 FILLER_0_1709 ();
 sg13g2_decap_8 FILLER_0_1716 ();
 sg13g2_decap_4 FILLER_0_1723 ();
 sg13g2_fill_1 FILLER_0_1727 ();
 sg13g2_fill_1 FILLER_0_1768 ();
 sg13g2_fill_2 FILLER_0_1774 ();
 sg13g2_fill_1 FILLER_0_1794 ();
 sg13g2_decap_4 FILLER_0_1804 ();
 sg13g2_fill_2 FILLER_0_1808 ();
 sg13g2_fill_2 FILLER_0_1819 ();
 sg13g2_decap_8 FILLER_0_1831 ();
 sg13g2_fill_2 FILLER_0_1838 ();
 sg13g2_fill_1 FILLER_0_1840 ();
 sg13g2_fill_2 FILLER_0_1860 ();
 sg13g2_decap_4 FILLER_0_1890 ();
 sg13g2_fill_1 FILLER_0_1894 ();
 sg13g2_decap_8 FILLER_0_1904 ();
 sg13g2_decap_8 FILLER_0_1911 ();
 sg13g2_decap_8 FILLER_0_1918 ();
 sg13g2_decap_8 FILLER_0_1925 ();
 sg13g2_decap_8 FILLER_0_1932 ();
 sg13g2_decap_8 FILLER_0_1939 ();
 sg13g2_decap_8 FILLER_0_1946 ();
 sg13g2_decap_8 FILLER_0_1953 ();
 sg13g2_decap_8 FILLER_0_1960 ();
 sg13g2_decap_8 FILLER_0_1967 ();
 sg13g2_decap_8 FILLER_0_1974 ();
 sg13g2_decap_8 FILLER_0_1981 ();
 sg13g2_decap_8 FILLER_0_1988 ();
 sg13g2_decap_8 FILLER_0_1995 ();
 sg13g2_decap_8 FILLER_0_2002 ();
 sg13g2_decap_8 FILLER_0_2009 ();
 sg13g2_decap_8 FILLER_0_2016 ();
 sg13g2_decap_8 FILLER_0_2023 ();
 sg13g2_decap_8 FILLER_0_2030 ();
 sg13g2_decap_8 FILLER_0_2037 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2051 ();
 sg13g2_decap_8 FILLER_0_2058 ();
 sg13g2_decap_8 FILLER_0_2065 ();
 sg13g2_decap_8 FILLER_0_2072 ();
 sg13g2_decap_8 FILLER_0_2079 ();
 sg13g2_decap_8 FILLER_0_2086 ();
 sg13g2_decap_8 FILLER_0_2093 ();
 sg13g2_decap_8 FILLER_0_2100 ();
 sg13g2_decap_8 FILLER_0_2107 ();
 sg13g2_decap_8 FILLER_0_2114 ();
 sg13g2_decap_8 FILLER_0_2121 ();
 sg13g2_decap_8 FILLER_0_2128 ();
 sg13g2_decap_8 FILLER_0_2135 ();
 sg13g2_decap_8 FILLER_0_2142 ();
 sg13g2_decap_8 FILLER_0_2149 ();
 sg13g2_decap_8 FILLER_0_2156 ();
 sg13g2_decap_8 FILLER_0_2163 ();
 sg13g2_decap_8 FILLER_0_2170 ();
 sg13g2_decap_8 FILLER_0_2177 ();
 sg13g2_decap_8 FILLER_0_2184 ();
 sg13g2_decap_8 FILLER_0_2191 ();
 sg13g2_decap_8 FILLER_0_2198 ();
 sg13g2_decap_8 FILLER_0_2205 ();
 sg13g2_decap_8 FILLER_0_2212 ();
 sg13g2_decap_8 FILLER_0_2219 ();
 sg13g2_decap_8 FILLER_0_2226 ();
 sg13g2_decap_8 FILLER_0_2233 ();
 sg13g2_decap_8 FILLER_0_2240 ();
 sg13g2_decap_8 FILLER_0_2247 ();
 sg13g2_decap_8 FILLER_0_2254 ();
 sg13g2_decap_8 FILLER_0_2261 ();
 sg13g2_decap_8 FILLER_0_2268 ();
 sg13g2_decap_8 FILLER_0_2275 ();
 sg13g2_decap_8 FILLER_0_2282 ();
 sg13g2_decap_8 FILLER_0_2289 ();
 sg13g2_decap_8 FILLER_0_2296 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_8 FILLER_0_2310 ();
 sg13g2_decap_8 FILLER_0_2317 ();
 sg13g2_decap_8 FILLER_0_2324 ();
 sg13g2_decap_8 FILLER_0_2331 ();
 sg13g2_decap_8 FILLER_0_2338 ();
 sg13g2_decap_8 FILLER_0_2345 ();
 sg13g2_decap_8 FILLER_0_2352 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_8 FILLER_0_2366 ();
 sg13g2_decap_8 FILLER_0_2373 ();
 sg13g2_decap_8 FILLER_0_2380 ();
 sg13g2_decap_8 FILLER_0_2387 ();
 sg13g2_decap_8 FILLER_0_2394 ();
 sg13g2_decap_8 FILLER_0_2401 ();
 sg13g2_decap_8 FILLER_0_2408 ();
 sg13g2_decap_8 FILLER_0_2415 ();
 sg13g2_decap_8 FILLER_0_2422 ();
 sg13g2_decap_8 FILLER_0_2429 ();
 sg13g2_decap_8 FILLER_0_2436 ();
 sg13g2_decap_8 FILLER_0_2443 ();
 sg13g2_decap_8 FILLER_0_2450 ();
 sg13g2_decap_8 FILLER_0_2457 ();
 sg13g2_decap_8 FILLER_0_2464 ();
 sg13g2_decap_8 FILLER_0_2471 ();
 sg13g2_decap_8 FILLER_0_2478 ();
 sg13g2_decap_8 FILLER_0_2485 ();
 sg13g2_decap_8 FILLER_0_2492 ();
 sg13g2_decap_8 FILLER_0_2499 ();
 sg13g2_decap_8 FILLER_0_2506 ();
 sg13g2_decap_8 FILLER_0_2513 ();
 sg13g2_decap_8 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2527 ();
 sg13g2_decap_8 FILLER_0_2534 ();
 sg13g2_decap_8 FILLER_0_2541 ();
 sg13g2_decap_8 FILLER_0_2548 ();
 sg13g2_decap_8 FILLER_0_2555 ();
 sg13g2_decap_8 FILLER_0_2562 ();
 sg13g2_decap_8 FILLER_0_2569 ();
 sg13g2_decap_8 FILLER_0_2576 ();
 sg13g2_decap_8 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_decap_8 FILLER_0_2597 ();
 sg13g2_decap_8 FILLER_0_2604 ();
 sg13g2_decap_8 FILLER_0_2611 ();
 sg13g2_decap_8 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2625 ();
 sg13g2_decap_8 FILLER_0_2632 ();
 sg13g2_decap_8 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2646 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_decap_8 FILLER_0_2667 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_169 ();
 sg13g2_fill_2 FILLER_1_175 ();
 sg13g2_fill_2 FILLER_1_217 ();
 sg13g2_fill_2 FILLER_1_246 ();
 sg13g2_fill_1 FILLER_1_248 ();
 sg13g2_decap_4 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_4 FILLER_1_322 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_decap_4 FILLER_1_364 ();
 sg13g2_fill_2 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_381 ();
 sg13g2_fill_1 FILLER_1_409 ();
 sg13g2_fill_1 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_452 ();
 sg13g2_decap_8 FILLER_1_486 ();
 sg13g2_decap_8 FILLER_1_493 ();
 sg13g2_decap_4 FILLER_1_500 ();
 sg13g2_decap_8 FILLER_1_527 ();
 sg13g2_fill_1 FILLER_1_534 ();
 sg13g2_fill_2 FILLER_1_548 ();
 sg13g2_fill_2 FILLER_1_568 ();
 sg13g2_fill_1 FILLER_1_641 ();
 sg13g2_fill_2 FILLER_1_676 ();
 sg13g2_fill_2 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_744 ();
 sg13g2_fill_1 FILLER_1_751 ();
 sg13g2_fill_2 FILLER_1_780 ();
 sg13g2_decap_4 FILLER_1_810 ();
 sg13g2_fill_1 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_843 ();
 sg13g2_fill_1 FILLER_1_850 ();
 sg13g2_decap_8 FILLER_1_886 ();
 sg13g2_decap_4 FILLER_1_893 ();
 sg13g2_fill_1 FILLER_1_897 ();
 sg13g2_decap_8 FILLER_1_982 ();
 sg13g2_fill_1 FILLER_1_989 ();
 sg13g2_fill_1 FILLER_1_994 ();
 sg13g2_decap_4 FILLER_1_1026 ();
 sg13g2_fill_1 FILLER_1_1030 ();
 sg13g2_fill_1 FILLER_1_1034 ();
 sg13g2_fill_2 FILLER_1_1110 ();
 sg13g2_fill_1 FILLER_1_1112 ();
 sg13g2_fill_1 FILLER_1_1122 ();
 sg13g2_fill_2 FILLER_1_1248 ();
 sg13g2_fill_1 FILLER_1_1250 ();
 sg13g2_fill_1 FILLER_1_1287 ();
 sg13g2_decap_8 FILLER_1_1363 ();
 sg13g2_fill_1 FILLER_1_1370 ();
 sg13g2_fill_1 FILLER_1_1399 ();
 sg13g2_decap_4 FILLER_1_1443 ();
 sg13g2_fill_1 FILLER_1_1447 ();
 sg13g2_fill_1 FILLER_1_1476 ();
 sg13g2_fill_2 FILLER_1_1486 ();
 sg13g2_fill_2 FILLER_1_1521 ();
 sg13g2_fill_2 FILLER_1_1528 ();
 sg13g2_decap_4 FILLER_1_1641 ();
 sg13g2_fill_2 FILLER_1_1678 ();
 sg13g2_fill_1 FILLER_1_1680 ();
 sg13g2_decap_4 FILLER_1_1708 ();
 sg13g2_fill_1 FILLER_1_1712 ();
 sg13g2_fill_2 FILLER_1_1750 ();
 sg13g2_fill_1 FILLER_1_1752 ();
 sg13g2_fill_2 FILLER_1_1762 ();
 sg13g2_fill_1 FILLER_1_1764 ();
 sg13g2_decap_4 FILLER_1_1793 ();
 sg13g2_decap_4 FILLER_1_1807 ();
 sg13g2_fill_1 FILLER_1_1811 ();
 sg13g2_fill_2 FILLER_1_1840 ();
 sg13g2_decap_4 FILLER_1_1879 ();
 sg13g2_fill_2 FILLER_1_1883 ();
 sg13g2_decap_8 FILLER_1_1904 ();
 sg13g2_decap_8 FILLER_1_1911 ();
 sg13g2_decap_8 FILLER_1_1918 ();
 sg13g2_decap_8 FILLER_1_1925 ();
 sg13g2_decap_8 FILLER_1_1932 ();
 sg13g2_decap_8 FILLER_1_1939 ();
 sg13g2_decap_8 FILLER_1_1946 ();
 sg13g2_decap_8 FILLER_1_1953 ();
 sg13g2_decap_8 FILLER_1_1960 ();
 sg13g2_decap_8 FILLER_1_1967 ();
 sg13g2_decap_8 FILLER_1_1974 ();
 sg13g2_decap_8 FILLER_1_1981 ();
 sg13g2_decap_8 FILLER_1_1988 ();
 sg13g2_decap_8 FILLER_1_1995 ();
 sg13g2_decap_8 FILLER_1_2002 ();
 sg13g2_decap_8 FILLER_1_2009 ();
 sg13g2_decap_8 FILLER_1_2016 ();
 sg13g2_decap_8 FILLER_1_2023 ();
 sg13g2_decap_8 FILLER_1_2030 ();
 sg13g2_decap_8 FILLER_1_2037 ();
 sg13g2_decap_8 FILLER_1_2044 ();
 sg13g2_decap_8 FILLER_1_2051 ();
 sg13g2_decap_8 FILLER_1_2058 ();
 sg13g2_decap_8 FILLER_1_2065 ();
 sg13g2_decap_8 FILLER_1_2072 ();
 sg13g2_decap_8 FILLER_1_2079 ();
 sg13g2_decap_8 FILLER_1_2086 ();
 sg13g2_decap_8 FILLER_1_2093 ();
 sg13g2_decap_8 FILLER_1_2100 ();
 sg13g2_decap_8 FILLER_1_2107 ();
 sg13g2_decap_8 FILLER_1_2114 ();
 sg13g2_decap_8 FILLER_1_2121 ();
 sg13g2_decap_8 FILLER_1_2128 ();
 sg13g2_decap_8 FILLER_1_2135 ();
 sg13g2_decap_8 FILLER_1_2142 ();
 sg13g2_decap_8 FILLER_1_2149 ();
 sg13g2_decap_8 FILLER_1_2156 ();
 sg13g2_decap_8 FILLER_1_2163 ();
 sg13g2_decap_8 FILLER_1_2170 ();
 sg13g2_decap_8 FILLER_1_2177 ();
 sg13g2_decap_8 FILLER_1_2184 ();
 sg13g2_decap_8 FILLER_1_2191 ();
 sg13g2_decap_8 FILLER_1_2198 ();
 sg13g2_decap_8 FILLER_1_2205 ();
 sg13g2_decap_8 FILLER_1_2212 ();
 sg13g2_decap_8 FILLER_1_2219 ();
 sg13g2_decap_8 FILLER_1_2226 ();
 sg13g2_decap_8 FILLER_1_2233 ();
 sg13g2_decap_8 FILLER_1_2240 ();
 sg13g2_decap_8 FILLER_1_2247 ();
 sg13g2_decap_8 FILLER_1_2254 ();
 sg13g2_decap_8 FILLER_1_2261 ();
 sg13g2_decap_8 FILLER_1_2268 ();
 sg13g2_decap_8 FILLER_1_2275 ();
 sg13g2_decap_8 FILLER_1_2282 ();
 sg13g2_decap_8 FILLER_1_2289 ();
 sg13g2_decap_8 FILLER_1_2296 ();
 sg13g2_decap_8 FILLER_1_2303 ();
 sg13g2_decap_8 FILLER_1_2310 ();
 sg13g2_decap_8 FILLER_1_2317 ();
 sg13g2_decap_8 FILLER_1_2324 ();
 sg13g2_decap_8 FILLER_1_2331 ();
 sg13g2_decap_8 FILLER_1_2338 ();
 sg13g2_decap_8 FILLER_1_2345 ();
 sg13g2_decap_8 FILLER_1_2352 ();
 sg13g2_decap_8 FILLER_1_2359 ();
 sg13g2_decap_8 FILLER_1_2366 ();
 sg13g2_decap_8 FILLER_1_2373 ();
 sg13g2_decap_8 FILLER_1_2380 ();
 sg13g2_decap_8 FILLER_1_2387 ();
 sg13g2_decap_8 FILLER_1_2394 ();
 sg13g2_decap_8 FILLER_1_2401 ();
 sg13g2_decap_8 FILLER_1_2408 ();
 sg13g2_decap_8 FILLER_1_2415 ();
 sg13g2_decap_8 FILLER_1_2422 ();
 sg13g2_decap_8 FILLER_1_2429 ();
 sg13g2_decap_8 FILLER_1_2436 ();
 sg13g2_decap_8 FILLER_1_2443 ();
 sg13g2_decap_8 FILLER_1_2450 ();
 sg13g2_decap_8 FILLER_1_2457 ();
 sg13g2_decap_8 FILLER_1_2464 ();
 sg13g2_decap_8 FILLER_1_2471 ();
 sg13g2_decap_8 FILLER_1_2478 ();
 sg13g2_decap_8 FILLER_1_2485 ();
 sg13g2_decap_8 FILLER_1_2492 ();
 sg13g2_decap_8 FILLER_1_2499 ();
 sg13g2_decap_8 FILLER_1_2506 ();
 sg13g2_decap_8 FILLER_1_2513 ();
 sg13g2_decap_8 FILLER_1_2520 ();
 sg13g2_decap_8 FILLER_1_2527 ();
 sg13g2_decap_8 FILLER_1_2534 ();
 sg13g2_decap_8 FILLER_1_2541 ();
 sg13g2_decap_8 FILLER_1_2548 ();
 sg13g2_decap_8 FILLER_1_2555 ();
 sg13g2_decap_8 FILLER_1_2562 ();
 sg13g2_decap_8 FILLER_1_2569 ();
 sg13g2_decap_8 FILLER_1_2576 ();
 sg13g2_decap_8 FILLER_1_2583 ();
 sg13g2_decap_8 FILLER_1_2590 ();
 sg13g2_decap_8 FILLER_1_2597 ();
 sg13g2_decap_8 FILLER_1_2604 ();
 sg13g2_decap_8 FILLER_1_2611 ();
 sg13g2_decap_8 FILLER_1_2618 ();
 sg13g2_decap_8 FILLER_1_2625 ();
 sg13g2_decap_8 FILLER_1_2632 ();
 sg13g2_decap_8 FILLER_1_2639 ();
 sg13g2_decap_8 FILLER_1_2646 ();
 sg13g2_decap_8 FILLER_1_2653 ();
 sg13g2_decap_8 FILLER_1_2660 ();
 sg13g2_decap_8 FILLER_1_2667 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_18 ();
 sg13g2_fill_1 FILLER_2_47 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_2 FILLER_2_147 ();
 sg13g2_fill_1 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_204 ();
 sg13g2_decap_4 FILLER_2_211 ();
 sg13g2_fill_1 FILLER_2_215 ();
 sg13g2_fill_2 FILLER_2_315 ();
 sg13g2_fill_1 FILLER_2_317 ();
 sg13g2_fill_2 FILLER_2_424 ();
 sg13g2_fill_1 FILLER_2_426 ();
 sg13g2_fill_2 FILLER_2_459 ();
 sg13g2_fill_1 FILLER_2_461 ();
 sg13g2_decap_8 FILLER_2_489 ();
 sg13g2_decap_4 FILLER_2_496 ();
 sg13g2_fill_1 FILLER_2_500 ();
 sg13g2_fill_2 FILLER_2_527 ();
 sg13g2_fill_1 FILLER_2_533 ();
 sg13g2_fill_1 FILLER_2_570 ();
 sg13g2_fill_1 FILLER_2_624 ();
 sg13g2_fill_1 FILLER_2_631 ();
 sg13g2_decap_4 FILLER_2_689 ();
 sg13g2_fill_1 FILLER_2_693 ();
 sg13g2_fill_2 FILLER_2_781 ();
 sg13g2_fill_1 FILLER_2_783 ();
 sg13g2_decap_4 FILLER_2_856 ();
 sg13g2_fill_1 FILLER_2_860 ();
 sg13g2_fill_2 FILLER_2_917 ();
 sg13g2_fill_1 FILLER_2_919 ();
 sg13g2_fill_1 FILLER_2_983 ();
 sg13g2_fill_1 FILLER_2_1031 ();
 sg13g2_fill_1 FILLER_2_1111 ();
 sg13g2_fill_1 FILLER_2_1236 ();
 sg13g2_fill_1 FILLER_2_1275 ();
 sg13g2_fill_1 FILLER_2_1405 ();
 sg13g2_fill_2 FILLER_2_1448 ();
 sg13g2_fill_1 FILLER_2_1450 ();
 sg13g2_fill_1 FILLER_2_1513 ();
 sg13g2_fill_1 FILLER_2_1569 ();
 sg13g2_fill_2 FILLER_2_1597 ();
 sg13g2_fill_2 FILLER_2_1648 ();
 sg13g2_fill_1 FILLER_2_1650 ();
 sg13g2_fill_1 FILLER_2_1661 ();
 sg13g2_fill_2 FILLER_2_1727 ();
 sg13g2_fill_1 FILLER_2_1748 ();
 sg13g2_fill_2 FILLER_2_1754 ();
 sg13g2_fill_1 FILLER_2_1774 ();
 sg13g2_decap_8 FILLER_2_1931 ();
 sg13g2_decap_8 FILLER_2_1938 ();
 sg13g2_decap_8 FILLER_2_1945 ();
 sg13g2_decap_8 FILLER_2_1952 ();
 sg13g2_decap_8 FILLER_2_1959 ();
 sg13g2_decap_8 FILLER_2_1966 ();
 sg13g2_decap_8 FILLER_2_1973 ();
 sg13g2_decap_8 FILLER_2_1980 ();
 sg13g2_decap_8 FILLER_2_1987 ();
 sg13g2_fill_2 FILLER_2_1994 ();
 sg13g2_decap_8 FILLER_2_2000 ();
 sg13g2_decap_8 FILLER_2_2007 ();
 sg13g2_decap_8 FILLER_2_2014 ();
 sg13g2_fill_2 FILLER_2_2021 ();
 sg13g2_fill_1 FILLER_2_2023 ();
 sg13g2_decap_8 FILLER_2_2052 ();
 sg13g2_decap_8 FILLER_2_2059 ();
 sg13g2_decap_8 FILLER_2_2066 ();
 sg13g2_decap_8 FILLER_2_2073 ();
 sg13g2_decap_8 FILLER_2_2080 ();
 sg13g2_decap_4 FILLER_2_2087 ();
 sg13g2_fill_1 FILLER_2_2091 ();
 sg13g2_decap_4 FILLER_2_2096 ();
 sg13g2_fill_2 FILLER_2_2100 ();
 sg13g2_decap_8 FILLER_2_2106 ();
 sg13g2_decap_8 FILLER_2_2113 ();
 sg13g2_decap_8 FILLER_2_2120 ();
 sg13g2_decap_8 FILLER_2_2127 ();
 sg13g2_decap_8 FILLER_2_2134 ();
 sg13g2_decap_8 FILLER_2_2141 ();
 sg13g2_decap_8 FILLER_2_2148 ();
 sg13g2_decap_8 FILLER_2_2155 ();
 sg13g2_decap_8 FILLER_2_2162 ();
 sg13g2_decap_8 FILLER_2_2169 ();
 sg13g2_decap_8 FILLER_2_2176 ();
 sg13g2_decap_8 FILLER_2_2183 ();
 sg13g2_decap_8 FILLER_2_2190 ();
 sg13g2_decap_8 FILLER_2_2197 ();
 sg13g2_decap_8 FILLER_2_2204 ();
 sg13g2_decap_8 FILLER_2_2211 ();
 sg13g2_decap_8 FILLER_2_2218 ();
 sg13g2_decap_8 FILLER_2_2225 ();
 sg13g2_decap_8 FILLER_2_2232 ();
 sg13g2_decap_8 FILLER_2_2239 ();
 sg13g2_decap_8 FILLER_2_2246 ();
 sg13g2_decap_8 FILLER_2_2253 ();
 sg13g2_decap_8 FILLER_2_2260 ();
 sg13g2_decap_8 FILLER_2_2267 ();
 sg13g2_decap_8 FILLER_2_2274 ();
 sg13g2_decap_8 FILLER_2_2281 ();
 sg13g2_decap_8 FILLER_2_2288 ();
 sg13g2_decap_8 FILLER_2_2295 ();
 sg13g2_decap_8 FILLER_2_2302 ();
 sg13g2_decap_8 FILLER_2_2309 ();
 sg13g2_decap_8 FILLER_2_2316 ();
 sg13g2_decap_8 FILLER_2_2323 ();
 sg13g2_decap_8 FILLER_2_2330 ();
 sg13g2_decap_8 FILLER_2_2337 ();
 sg13g2_decap_8 FILLER_2_2344 ();
 sg13g2_decap_8 FILLER_2_2351 ();
 sg13g2_decap_8 FILLER_2_2358 ();
 sg13g2_decap_8 FILLER_2_2365 ();
 sg13g2_decap_8 FILLER_2_2372 ();
 sg13g2_decap_8 FILLER_2_2379 ();
 sg13g2_decap_8 FILLER_2_2386 ();
 sg13g2_decap_8 FILLER_2_2393 ();
 sg13g2_decap_8 FILLER_2_2400 ();
 sg13g2_decap_8 FILLER_2_2407 ();
 sg13g2_decap_8 FILLER_2_2414 ();
 sg13g2_decap_8 FILLER_2_2421 ();
 sg13g2_decap_8 FILLER_2_2428 ();
 sg13g2_decap_8 FILLER_2_2435 ();
 sg13g2_decap_8 FILLER_2_2442 ();
 sg13g2_decap_8 FILLER_2_2449 ();
 sg13g2_decap_8 FILLER_2_2456 ();
 sg13g2_decap_8 FILLER_2_2463 ();
 sg13g2_decap_8 FILLER_2_2470 ();
 sg13g2_decap_8 FILLER_2_2477 ();
 sg13g2_decap_8 FILLER_2_2484 ();
 sg13g2_decap_8 FILLER_2_2491 ();
 sg13g2_decap_8 FILLER_2_2498 ();
 sg13g2_decap_8 FILLER_2_2505 ();
 sg13g2_decap_8 FILLER_2_2512 ();
 sg13g2_decap_8 FILLER_2_2519 ();
 sg13g2_decap_8 FILLER_2_2526 ();
 sg13g2_decap_8 FILLER_2_2533 ();
 sg13g2_decap_8 FILLER_2_2540 ();
 sg13g2_decap_8 FILLER_2_2547 ();
 sg13g2_decap_8 FILLER_2_2554 ();
 sg13g2_decap_8 FILLER_2_2561 ();
 sg13g2_decap_8 FILLER_2_2568 ();
 sg13g2_decap_8 FILLER_2_2575 ();
 sg13g2_decap_8 FILLER_2_2582 ();
 sg13g2_decap_8 FILLER_2_2589 ();
 sg13g2_decap_8 FILLER_2_2596 ();
 sg13g2_decap_8 FILLER_2_2603 ();
 sg13g2_decap_8 FILLER_2_2610 ();
 sg13g2_decap_8 FILLER_2_2617 ();
 sg13g2_decap_8 FILLER_2_2624 ();
 sg13g2_decap_8 FILLER_2_2631 ();
 sg13g2_decap_8 FILLER_2_2638 ();
 sg13g2_decap_8 FILLER_2_2645 ();
 sg13g2_decap_8 FILLER_2_2652 ();
 sg13g2_decap_8 FILLER_2_2659 ();
 sg13g2_decap_8 FILLER_2_2666 ();
 sg13g2_fill_1 FILLER_2_2673 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_67 ();
 sg13g2_fill_2 FILLER_3_109 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_208 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_fill_2 FILLER_3_266 ();
 sg13g2_fill_2 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_310 ();
 sg13g2_fill_2 FILLER_3_320 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_decap_4 FILLER_3_449 ();
 sg13g2_decap_4 FILLER_3_488 ();
 sg13g2_fill_2 FILLER_3_535 ();
 sg13g2_fill_1 FILLER_3_537 ();
 sg13g2_fill_1 FILLER_3_617 ();
 sg13g2_fill_2 FILLER_3_653 ();
 sg13g2_fill_1 FILLER_3_655 ();
 sg13g2_fill_1 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_692 ();
 sg13g2_fill_1 FILLER_3_699 ();
 sg13g2_fill_2 FILLER_3_740 ();
 sg13g2_fill_2 FILLER_3_784 ();
 sg13g2_fill_1 FILLER_3_786 ();
 sg13g2_decap_4 FILLER_3_814 ();
 sg13g2_fill_2 FILLER_3_818 ();
 sg13g2_fill_1 FILLER_3_954 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_fill_2 FILLER_3_1028 ();
 sg13g2_fill_1 FILLER_3_1030 ();
 sg13g2_decap_4 FILLER_3_1068 ();
 sg13g2_fill_2 FILLER_3_1081 ();
 sg13g2_fill_2 FILLER_3_1203 ();
 sg13g2_fill_2 FILLER_3_1250 ();
 sg13g2_fill_2 FILLER_3_1262 ();
 sg13g2_fill_1 FILLER_3_1264 ();
 sg13g2_fill_1 FILLER_3_1278 ();
 sg13g2_decap_4 FILLER_3_1338 ();
 sg13g2_fill_1 FILLER_3_1411 ();
 sg13g2_decap_4 FILLER_3_1452 ();
 sg13g2_fill_1 FILLER_3_1456 ();
 sg13g2_fill_2 FILLER_3_1529 ();
 sg13g2_fill_1 FILLER_3_1531 ();
 sg13g2_fill_1 FILLER_3_1601 ();
 sg13g2_fill_1 FILLER_3_1612 ();
 sg13g2_fill_2 FILLER_3_1742 ();
 sg13g2_fill_2 FILLER_3_1749 ();
 sg13g2_fill_2 FILLER_3_1771 ();
 sg13g2_fill_1 FILLER_3_1773 ();
 sg13g2_decap_4 FILLER_3_1830 ();
 sg13g2_decap_8 FILLER_3_1847 ();
 sg13g2_fill_1 FILLER_3_1854 ();
 sg13g2_decap_8 FILLER_3_1932 ();
 sg13g2_decap_8 FILLER_3_1939 ();
 sg13g2_decap_8 FILLER_3_1946 ();
 sg13g2_decap_8 FILLER_3_1953 ();
 sg13g2_decap_8 FILLER_3_1960 ();
 sg13g2_decap_8 FILLER_3_1967 ();
 sg13g2_fill_1 FILLER_3_1974 ();
 sg13g2_decap_8 FILLER_3_2007 ();
 sg13g2_decap_8 FILLER_3_2014 ();
 sg13g2_decap_4 FILLER_3_2021 ();
 sg13g2_fill_1 FILLER_3_2025 ();
 sg13g2_decap_8 FILLER_3_2063 ();
 sg13g2_fill_2 FILLER_3_2070 ();
 sg13g2_fill_2 FILLER_3_2100 ();
 sg13g2_fill_1 FILLER_3_2102 ();
 sg13g2_decap_4 FILLER_3_2112 ();
 sg13g2_fill_1 FILLER_3_2116 ();
 sg13g2_decap_8 FILLER_3_2126 ();
 sg13g2_decap_8 FILLER_3_2133 ();
 sg13g2_decap_8 FILLER_3_2140 ();
 sg13g2_decap_8 FILLER_3_2147 ();
 sg13g2_decap_8 FILLER_3_2154 ();
 sg13g2_decap_8 FILLER_3_2161 ();
 sg13g2_decap_8 FILLER_3_2168 ();
 sg13g2_decap_8 FILLER_3_2175 ();
 sg13g2_decap_8 FILLER_3_2182 ();
 sg13g2_decap_8 FILLER_3_2189 ();
 sg13g2_decap_8 FILLER_3_2196 ();
 sg13g2_decap_8 FILLER_3_2203 ();
 sg13g2_decap_8 FILLER_3_2210 ();
 sg13g2_decap_8 FILLER_3_2217 ();
 sg13g2_decap_8 FILLER_3_2224 ();
 sg13g2_decap_8 FILLER_3_2231 ();
 sg13g2_decap_8 FILLER_3_2238 ();
 sg13g2_decap_8 FILLER_3_2245 ();
 sg13g2_decap_8 FILLER_3_2252 ();
 sg13g2_decap_8 FILLER_3_2259 ();
 sg13g2_decap_8 FILLER_3_2266 ();
 sg13g2_decap_8 FILLER_3_2273 ();
 sg13g2_decap_8 FILLER_3_2280 ();
 sg13g2_decap_8 FILLER_3_2287 ();
 sg13g2_decap_8 FILLER_3_2294 ();
 sg13g2_decap_8 FILLER_3_2301 ();
 sg13g2_decap_8 FILLER_3_2308 ();
 sg13g2_decap_8 FILLER_3_2315 ();
 sg13g2_decap_8 FILLER_3_2322 ();
 sg13g2_decap_8 FILLER_3_2329 ();
 sg13g2_decap_8 FILLER_3_2336 ();
 sg13g2_decap_8 FILLER_3_2343 ();
 sg13g2_decap_8 FILLER_3_2350 ();
 sg13g2_decap_8 FILLER_3_2357 ();
 sg13g2_decap_8 FILLER_3_2364 ();
 sg13g2_decap_8 FILLER_3_2371 ();
 sg13g2_decap_8 FILLER_3_2378 ();
 sg13g2_decap_8 FILLER_3_2385 ();
 sg13g2_decap_8 FILLER_3_2392 ();
 sg13g2_decap_8 FILLER_3_2399 ();
 sg13g2_decap_8 FILLER_3_2406 ();
 sg13g2_decap_8 FILLER_3_2413 ();
 sg13g2_decap_8 FILLER_3_2420 ();
 sg13g2_decap_8 FILLER_3_2427 ();
 sg13g2_decap_8 FILLER_3_2434 ();
 sg13g2_decap_8 FILLER_3_2441 ();
 sg13g2_decap_8 FILLER_3_2448 ();
 sg13g2_decap_8 FILLER_3_2455 ();
 sg13g2_decap_8 FILLER_3_2462 ();
 sg13g2_decap_8 FILLER_3_2469 ();
 sg13g2_decap_8 FILLER_3_2476 ();
 sg13g2_decap_8 FILLER_3_2483 ();
 sg13g2_decap_8 FILLER_3_2490 ();
 sg13g2_decap_8 FILLER_3_2497 ();
 sg13g2_decap_8 FILLER_3_2504 ();
 sg13g2_decap_8 FILLER_3_2511 ();
 sg13g2_decap_8 FILLER_3_2518 ();
 sg13g2_decap_8 FILLER_3_2525 ();
 sg13g2_decap_8 FILLER_3_2532 ();
 sg13g2_decap_8 FILLER_3_2539 ();
 sg13g2_decap_8 FILLER_3_2546 ();
 sg13g2_decap_8 FILLER_3_2553 ();
 sg13g2_decap_8 FILLER_3_2560 ();
 sg13g2_decap_8 FILLER_3_2567 ();
 sg13g2_decap_8 FILLER_3_2574 ();
 sg13g2_decap_8 FILLER_3_2581 ();
 sg13g2_decap_8 FILLER_3_2588 ();
 sg13g2_decap_8 FILLER_3_2595 ();
 sg13g2_decap_8 FILLER_3_2602 ();
 sg13g2_decap_8 FILLER_3_2609 ();
 sg13g2_decap_8 FILLER_3_2616 ();
 sg13g2_decap_8 FILLER_3_2623 ();
 sg13g2_decap_8 FILLER_3_2630 ();
 sg13g2_decap_8 FILLER_3_2637 ();
 sg13g2_decap_8 FILLER_3_2644 ();
 sg13g2_decap_8 FILLER_3_2651 ();
 sg13g2_decap_8 FILLER_3_2658 ();
 sg13g2_decap_8 FILLER_3_2665 ();
 sg13g2_fill_2 FILLER_3_2672 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_35 ();
 sg13g2_fill_2 FILLER_4_40 ();
 sg13g2_fill_2 FILLER_4_51 ();
 sg13g2_fill_2 FILLER_4_58 ();
 sg13g2_fill_2 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_fill_1 FILLER_4_169 ();
 sg13g2_fill_2 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_204 ();
 sg13g2_decap_4 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_222 ();
 sg13g2_fill_2 FILLER_4_241 ();
 sg13g2_fill_2 FILLER_4_248 ();
 sg13g2_fill_2 FILLER_4_264 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_296 ();
 sg13g2_fill_2 FILLER_4_316 ();
 sg13g2_fill_1 FILLER_4_318 ();
 sg13g2_fill_2 FILLER_4_396 ();
 sg13g2_fill_2 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_fill_2 FILLER_4_434 ();
 sg13g2_fill_1 FILLER_4_436 ();
 sg13g2_fill_1 FILLER_4_444 ();
 sg13g2_fill_1 FILLER_4_478 ();
 sg13g2_decap_8 FILLER_4_484 ();
 sg13g2_decap_4 FILLER_4_491 ();
 sg13g2_fill_2 FILLER_4_531 ();
 sg13g2_fill_1 FILLER_4_561 ();
 sg13g2_fill_1 FILLER_4_577 ();
 sg13g2_decap_4 FILLER_4_619 ();
 sg13g2_fill_2 FILLER_4_623 ();
 sg13g2_fill_2 FILLER_4_641 ();
 sg13g2_fill_1 FILLER_4_643 ();
 sg13g2_decap_4 FILLER_4_653 ();
 sg13g2_fill_1 FILLER_4_657 ();
 sg13g2_fill_2 FILLER_4_667 ();
 sg13g2_fill_1 FILLER_4_681 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_fill_2 FILLER_4_704 ();
 sg13g2_fill_2 FILLER_4_709 ();
 sg13g2_fill_1 FILLER_4_711 ();
 sg13g2_fill_1 FILLER_4_720 ();
 sg13g2_fill_1 FILLER_4_739 ();
 sg13g2_fill_2 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_958 ();
 sg13g2_fill_1 FILLER_4_995 ();
 sg13g2_decap_8 FILLER_4_1018 ();
 sg13g2_decap_8 FILLER_4_1025 ();
 sg13g2_decap_8 FILLER_4_1032 ();
 sg13g2_decap_4 FILLER_4_1039 ();
 sg13g2_decap_4 FILLER_4_1070 ();
 sg13g2_fill_2 FILLER_4_1074 ();
 sg13g2_fill_2 FILLER_4_1083 ();
 sg13g2_fill_1 FILLER_4_1085 ();
 sg13g2_fill_2 FILLER_4_1102 ();
 sg13g2_fill_1 FILLER_4_1191 ();
 sg13g2_fill_2 FILLER_4_1205 ();
 sg13g2_fill_1 FILLER_4_1225 ();
 sg13g2_fill_2 FILLER_4_1266 ();
 sg13g2_fill_2 FILLER_4_1297 ();
 sg13g2_decap_8 FILLER_4_1326 ();
 sg13g2_decap_4 FILLER_4_1333 ();
 sg13g2_fill_2 FILLER_4_1344 ();
 sg13g2_decap_8 FILLER_4_1355 ();
 sg13g2_decap_4 FILLER_4_1362 ();
 sg13g2_fill_2 FILLER_4_1366 ();
 sg13g2_fill_2 FILLER_4_1458 ();
 sg13g2_fill_1 FILLER_4_1460 ();
 sg13g2_fill_1 FILLER_4_1475 ();
 sg13g2_fill_2 FILLER_4_1495 ();
 sg13g2_fill_2 FILLER_4_1552 ();
 sg13g2_fill_1 FILLER_4_1554 ();
 sg13g2_fill_1 FILLER_4_1622 ();
 sg13g2_fill_1 FILLER_4_1665 ();
 sg13g2_fill_2 FILLER_4_1716 ();
 sg13g2_fill_1 FILLER_4_1718 ();
 sg13g2_fill_2 FILLER_4_1732 ();
 sg13g2_fill_1 FILLER_4_1753 ();
 sg13g2_fill_2 FILLER_4_1759 ();
 sg13g2_fill_2 FILLER_4_1771 ();
 sg13g2_decap_4 FILLER_4_1833 ();
 sg13g2_fill_1 FILLER_4_1837 ();
 sg13g2_decap_8 FILLER_4_1944 ();
 sg13g2_decap_4 FILLER_4_1951 ();
 sg13g2_decap_4 FILLER_4_2013 ();
 sg13g2_fill_1 FILLER_4_2057 ();
 sg13g2_fill_2 FILLER_4_2077 ();
 sg13g2_fill_2 FILLER_4_2092 ();
 sg13g2_decap_8 FILLER_4_2131 ();
 sg13g2_decap_8 FILLER_4_2138 ();
 sg13g2_decap_8 FILLER_4_2145 ();
 sg13g2_decap_8 FILLER_4_2152 ();
 sg13g2_decap_8 FILLER_4_2159 ();
 sg13g2_decap_8 FILLER_4_2166 ();
 sg13g2_decap_8 FILLER_4_2173 ();
 sg13g2_decap_8 FILLER_4_2180 ();
 sg13g2_decap_8 FILLER_4_2187 ();
 sg13g2_decap_8 FILLER_4_2194 ();
 sg13g2_decap_8 FILLER_4_2201 ();
 sg13g2_decap_8 FILLER_4_2208 ();
 sg13g2_decap_8 FILLER_4_2215 ();
 sg13g2_decap_8 FILLER_4_2222 ();
 sg13g2_decap_8 FILLER_4_2229 ();
 sg13g2_decap_8 FILLER_4_2236 ();
 sg13g2_decap_8 FILLER_4_2243 ();
 sg13g2_decap_8 FILLER_4_2250 ();
 sg13g2_decap_8 FILLER_4_2257 ();
 sg13g2_decap_8 FILLER_4_2264 ();
 sg13g2_decap_8 FILLER_4_2271 ();
 sg13g2_decap_8 FILLER_4_2278 ();
 sg13g2_decap_8 FILLER_4_2285 ();
 sg13g2_decap_8 FILLER_4_2292 ();
 sg13g2_decap_8 FILLER_4_2299 ();
 sg13g2_decap_8 FILLER_4_2306 ();
 sg13g2_decap_8 FILLER_4_2313 ();
 sg13g2_decap_8 FILLER_4_2320 ();
 sg13g2_decap_8 FILLER_4_2327 ();
 sg13g2_decap_8 FILLER_4_2334 ();
 sg13g2_decap_8 FILLER_4_2341 ();
 sg13g2_decap_8 FILLER_4_2348 ();
 sg13g2_decap_8 FILLER_4_2355 ();
 sg13g2_decap_8 FILLER_4_2362 ();
 sg13g2_decap_8 FILLER_4_2369 ();
 sg13g2_decap_8 FILLER_4_2376 ();
 sg13g2_decap_8 FILLER_4_2383 ();
 sg13g2_decap_8 FILLER_4_2390 ();
 sg13g2_decap_8 FILLER_4_2397 ();
 sg13g2_decap_8 FILLER_4_2404 ();
 sg13g2_decap_8 FILLER_4_2411 ();
 sg13g2_decap_8 FILLER_4_2418 ();
 sg13g2_decap_8 FILLER_4_2425 ();
 sg13g2_decap_8 FILLER_4_2432 ();
 sg13g2_decap_8 FILLER_4_2439 ();
 sg13g2_decap_8 FILLER_4_2446 ();
 sg13g2_decap_8 FILLER_4_2453 ();
 sg13g2_decap_8 FILLER_4_2460 ();
 sg13g2_decap_8 FILLER_4_2467 ();
 sg13g2_decap_8 FILLER_4_2474 ();
 sg13g2_decap_8 FILLER_4_2481 ();
 sg13g2_decap_8 FILLER_4_2488 ();
 sg13g2_decap_8 FILLER_4_2495 ();
 sg13g2_decap_8 FILLER_4_2502 ();
 sg13g2_decap_8 FILLER_4_2509 ();
 sg13g2_decap_8 FILLER_4_2516 ();
 sg13g2_decap_8 FILLER_4_2523 ();
 sg13g2_decap_8 FILLER_4_2530 ();
 sg13g2_decap_8 FILLER_4_2537 ();
 sg13g2_decap_8 FILLER_4_2544 ();
 sg13g2_decap_8 FILLER_4_2551 ();
 sg13g2_decap_8 FILLER_4_2558 ();
 sg13g2_decap_8 FILLER_4_2565 ();
 sg13g2_decap_8 FILLER_4_2572 ();
 sg13g2_decap_8 FILLER_4_2579 ();
 sg13g2_decap_8 FILLER_4_2586 ();
 sg13g2_decap_8 FILLER_4_2593 ();
 sg13g2_decap_8 FILLER_4_2600 ();
 sg13g2_decap_8 FILLER_4_2607 ();
 sg13g2_decap_8 FILLER_4_2614 ();
 sg13g2_decap_8 FILLER_4_2621 ();
 sg13g2_decap_8 FILLER_4_2628 ();
 sg13g2_decap_8 FILLER_4_2635 ();
 sg13g2_decap_8 FILLER_4_2642 ();
 sg13g2_decap_8 FILLER_4_2649 ();
 sg13g2_decap_8 FILLER_4_2656 ();
 sg13g2_decap_8 FILLER_4_2663 ();
 sg13g2_decap_4 FILLER_4_2670 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_44 ();
 sg13g2_fill_1 FILLER_5_100 ();
 sg13g2_fill_1 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_fill_2 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_fill_2 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_270 ();
 sg13g2_fill_1 FILLER_5_272 ();
 sg13g2_fill_2 FILLER_5_300 ();
 sg13g2_fill_1 FILLER_5_302 ();
 sg13g2_fill_2 FILLER_5_356 ();
 sg13g2_fill_1 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_430 ();
 sg13g2_decap_8 FILLER_5_437 ();
 sg13g2_decap_4 FILLER_5_444 ();
 sg13g2_fill_2 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_477 ();
 sg13g2_decap_8 FILLER_5_484 ();
 sg13g2_decap_8 FILLER_5_491 ();
 sg13g2_decap_8 FILLER_5_498 ();
 sg13g2_fill_1 FILLER_5_505 ();
 sg13g2_fill_1 FILLER_5_511 ();
 sg13g2_decap_4 FILLER_5_537 ();
 sg13g2_fill_2 FILLER_5_546 ();
 sg13g2_fill_1 FILLER_5_548 ();
 sg13g2_fill_2 FILLER_5_559 ();
 sg13g2_fill_1 FILLER_5_561 ();
 sg13g2_decap_4 FILLER_5_567 ();
 sg13g2_fill_2 FILLER_5_571 ();
 sg13g2_fill_1 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_600 ();
 sg13g2_fill_2 FILLER_5_607 ();
 sg13g2_fill_1 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_fill_1 FILLER_5_637 ();
 sg13g2_decap_4 FILLER_5_654 ();
 sg13g2_fill_1 FILLER_5_658 ();
 sg13g2_fill_2 FILLER_5_699 ();
 sg13g2_fill_2 FILLER_5_704 ();
 sg13g2_fill_2 FILLER_5_734 ();
 sg13g2_fill_1 FILLER_5_767 ();
 sg13g2_fill_1 FILLER_5_781 ();
 sg13g2_fill_2 FILLER_5_797 ();
 sg13g2_fill_1 FILLER_5_860 ();
 sg13g2_fill_2 FILLER_5_896 ();
 sg13g2_decap_8 FILLER_5_911 ();
 sg13g2_decap_4 FILLER_5_918 ();
 sg13g2_decap_8 FILLER_5_957 ();
 sg13g2_fill_1 FILLER_5_964 ();
 sg13g2_fill_1 FILLER_5_981 ();
 sg13g2_fill_1 FILLER_5_1003 ();
 sg13g2_decap_8 FILLER_5_1009 ();
 sg13g2_fill_2 FILLER_5_1016 ();
 sg13g2_fill_2 FILLER_5_1024 ();
 sg13g2_decap_8 FILLER_5_1031 ();
 sg13g2_fill_2 FILLER_5_1121 ();
 sg13g2_fill_2 FILLER_5_1138 ();
 sg13g2_fill_1 FILLER_5_1191 ();
 sg13g2_fill_1 FILLER_5_1243 ();
 sg13g2_fill_2 FILLER_5_1315 ();
 sg13g2_decap_4 FILLER_5_1326 ();
 sg13g2_fill_2 FILLER_5_1330 ();
 sg13g2_decap_4 FILLER_5_1341 ();
 sg13g2_fill_2 FILLER_5_1345 ();
 sg13g2_decap_8 FILLER_5_1356 ();
 sg13g2_decap_4 FILLER_5_1363 ();
 sg13g2_fill_2 FILLER_5_1367 ();
 sg13g2_fill_2 FILLER_5_1378 ();
 sg13g2_fill_2 FILLER_5_1394 ();
 sg13g2_fill_2 FILLER_5_1405 ();
 sg13g2_fill_1 FILLER_5_1407 ();
 sg13g2_fill_1 FILLER_5_1450 ();
 sg13g2_fill_1 FILLER_5_1480 ();
 sg13g2_fill_1 FILLER_5_1612 ();
 sg13g2_fill_2 FILLER_5_1668 ();
 sg13g2_fill_1 FILLER_5_1685 ();
 sg13g2_fill_1 FILLER_5_1699 ();
 sg13g2_fill_2 FILLER_5_1709 ();
 sg13g2_fill_2 FILLER_5_1746 ();
 sg13g2_fill_1 FILLER_5_1748 ();
 sg13g2_fill_1 FILLER_5_1786 ();
 sg13g2_decap_4 FILLER_5_1817 ();
 sg13g2_fill_1 FILLER_5_1840 ();
 sg13g2_fill_2 FILLER_5_1845 ();
 sg13g2_decap_4 FILLER_5_1866 ();
 sg13g2_fill_1 FILLER_5_1870 ();
 sg13g2_fill_2 FILLER_5_1881 ();
 sg13g2_fill_1 FILLER_5_1883 ();
 sg13g2_decap_8 FILLER_5_1929 ();
 sg13g2_decap_8 FILLER_5_1936 ();
 sg13g2_decap_8 FILLER_5_1943 ();
 sg13g2_decap_8 FILLER_5_1950 ();
 sg13g2_decap_4 FILLER_5_1957 ();
 sg13g2_fill_2 FILLER_5_1961 ();
 sg13g2_fill_1 FILLER_5_2018 ();
 sg13g2_decap_4 FILLER_5_2023 ();
 sg13g2_fill_1 FILLER_5_2027 ();
 sg13g2_fill_2 FILLER_5_2042 ();
 sg13g2_fill_1 FILLER_5_2044 ();
 sg13g2_fill_2 FILLER_5_2095 ();
 sg13g2_fill_1 FILLER_5_2097 ();
 sg13g2_decap_8 FILLER_5_2107 ();
 sg13g2_decap_8 FILLER_5_2114 ();
 sg13g2_decap_8 FILLER_5_2121 ();
 sg13g2_decap_8 FILLER_5_2128 ();
 sg13g2_decap_8 FILLER_5_2135 ();
 sg13g2_decap_8 FILLER_5_2142 ();
 sg13g2_decap_8 FILLER_5_2149 ();
 sg13g2_decap_8 FILLER_5_2156 ();
 sg13g2_decap_8 FILLER_5_2163 ();
 sg13g2_decap_8 FILLER_5_2170 ();
 sg13g2_decap_8 FILLER_5_2177 ();
 sg13g2_decap_8 FILLER_5_2184 ();
 sg13g2_decap_8 FILLER_5_2191 ();
 sg13g2_decap_8 FILLER_5_2198 ();
 sg13g2_decap_8 FILLER_5_2205 ();
 sg13g2_decap_8 FILLER_5_2212 ();
 sg13g2_decap_8 FILLER_5_2219 ();
 sg13g2_decap_8 FILLER_5_2226 ();
 sg13g2_decap_8 FILLER_5_2233 ();
 sg13g2_decap_8 FILLER_5_2240 ();
 sg13g2_decap_8 FILLER_5_2247 ();
 sg13g2_decap_8 FILLER_5_2254 ();
 sg13g2_decap_8 FILLER_5_2261 ();
 sg13g2_decap_8 FILLER_5_2268 ();
 sg13g2_decap_8 FILLER_5_2275 ();
 sg13g2_decap_8 FILLER_5_2282 ();
 sg13g2_decap_8 FILLER_5_2289 ();
 sg13g2_decap_8 FILLER_5_2296 ();
 sg13g2_decap_8 FILLER_5_2303 ();
 sg13g2_decap_8 FILLER_5_2310 ();
 sg13g2_decap_8 FILLER_5_2317 ();
 sg13g2_decap_8 FILLER_5_2324 ();
 sg13g2_decap_8 FILLER_5_2331 ();
 sg13g2_decap_8 FILLER_5_2338 ();
 sg13g2_decap_8 FILLER_5_2345 ();
 sg13g2_decap_8 FILLER_5_2352 ();
 sg13g2_decap_8 FILLER_5_2359 ();
 sg13g2_decap_8 FILLER_5_2366 ();
 sg13g2_decap_8 FILLER_5_2373 ();
 sg13g2_decap_8 FILLER_5_2380 ();
 sg13g2_decap_8 FILLER_5_2387 ();
 sg13g2_decap_8 FILLER_5_2394 ();
 sg13g2_decap_8 FILLER_5_2401 ();
 sg13g2_decap_8 FILLER_5_2408 ();
 sg13g2_decap_8 FILLER_5_2415 ();
 sg13g2_decap_8 FILLER_5_2422 ();
 sg13g2_decap_8 FILLER_5_2429 ();
 sg13g2_decap_8 FILLER_5_2436 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2450 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_decap_8 FILLER_5_2464 ();
 sg13g2_decap_8 FILLER_5_2471 ();
 sg13g2_decap_8 FILLER_5_2478 ();
 sg13g2_decap_8 FILLER_5_2485 ();
 sg13g2_decap_8 FILLER_5_2492 ();
 sg13g2_decap_8 FILLER_5_2499 ();
 sg13g2_decap_8 FILLER_5_2506 ();
 sg13g2_decap_8 FILLER_5_2513 ();
 sg13g2_decap_8 FILLER_5_2520 ();
 sg13g2_decap_8 FILLER_5_2527 ();
 sg13g2_decap_8 FILLER_5_2534 ();
 sg13g2_decap_8 FILLER_5_2541 ();
 sg13g2_decap_8 FILLER_5_2548 ();
 sg13g2_decap_8 FILLER_5_2555 ();
 sg13g2_decap_8 FILLER_5_2562 ();
 sg13g2_decap_8 FILLER_5_2569 ();
 sg13g2_decap_8 FILLER_5_2576 ();
 sg13g2_decap_8 FILLER_5_2583 ();
 sg13g2_decap_8 FILLER_5_2590 ();
 sg13g2_decap_8 FILLER_5_2597 ();
 sg13g2_decap_8 FILLER_5_2604 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_decap_8 FILLER_5_2667 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_37 ();
 sg13g2_decap_4 FILLER_6_102 ();
 sg13g2_fill_2 FILLER_6_106 ();
 sg13g2_fill_2 FILLER_6_168 ();
 sg13g2_fill_1 FILLER_6_170 ();
 sg13g2_fill_2 FILLER_6_239 ();
 sg13g2_fill_2 FILLER_6_282 ();
 sg13g2_fill_1 FILLER_6_302 ();
 sg13g2_fill_1 FILLER_6_380 ();
 sg13g2_fill_1 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_425 ();
 sg13g2_fill_2 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_488 ();
 sg13g2_decap_4 FILLER_6_495 ();
 sg13g2_fill_1 FILLER_6_499 ();
 sg13g2_fill_1 FILLER_6_517 ();
 sg13g2_fill_2 FILLER_6_528 ();
 sg13g2_fill_2 FILLER_6_540 ();
 sg13g2_fill_1 FILLER_6_542 ();
 sg13g2_decap_4 FILLER_6_553 ();
 sg13g2_fill_1 FILLER_6_557 ();
 sg13g2_decap_4 FILLER_6_562 ();
 sg13g2_fill_1 FILLER_6_566 ();
 sg13g2_fill_2 FILLER_6_582 ();
 sg13g2_fill_1 FILLER_6_584 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_4 FILLER_6_623 ();
 sg13g2_fill_1 FILLER_6_627 ();
 sg13g2_fill_2 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_654 ();
 sg13g2_decap_4 FILLER_6_661 ();
 sg13g2_fill_1 FILLER_6_665 ();
 sg13g2_fill_2 FILLER_6_674 ();
 sg13g2_fill_1 FILLER_6_676 ();
 sg13g2_fill_2 FILLER_6_683 ();
 sg13g2_fill_1 FILLER_6_685 ();
 sg13g2_fill_1 FILLER_6_691 ();
 sg13g2_fill_2 FILLER_6_701 ();
 sg13g2_fill_2 FILLER_6_728 ();
 sg13g2_fill_1 FILLER_6_730 ();
 sg13g2_fill_1 FILLER_6_759 ();
 sg13g2_fill_1 FILLER_6_805 ();
 sg13g2_fill_1 FILLER_6_875 ();
 sg13g2_decap_4 FILLER_6_917 ();
 sg13g2_fill_1 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_926 ();
 sg13g2_fill_2 FILLER_6_933 ();
 sg13g2_decap_8 FILLER_6_948 ();
 sg13g2_decap_4 FILLER_6_955 ();
 sg13g2_decap_4 FILLER_6_1000 ();
 sg13g2_fill_2 FILLER_6_1004 ();
 sg13g2_fill_1 FILLER_6_1021 ();
 sg13g2_fill_1 FILLER_6_1030 ();
 sg13g2_fill_1 FILLER_6_1044 ();
 sg13g2_decap_4 FILLER_6_1050 ();
 sg13g2_fill_1 FILLER_6_1054 ();
 sg13g2_fill_1 FILLER_6_1068 ();
 sg13g2_decap_8 FILLER_6_1077 ();
 sg13g2_fill_2 FILLER_6_1084 ();
 sg13g2_decap_4 FILLER_6_1123 ();
 sg13g2_fill_2 FILLER_6_1206 ();
 sg13g2_fill_1 FILLER_6_1241 ();
 sg13g2_fill_2 FILLER_6_1307 ();
 sg13g2_decap_4 FILLER_6_1321 ();
 sg13g2_fill_1 FILLER_6_1381 ();
 sg13g2_fill_2 FILLER_6_1404 ();
 sg13g2_fill_1 FILLER_6_1445 ();
 sg13g2_fill_2 FILLER_6_1460 ();
 sg13g2_fill_1 FILLER_6_1462 ();
 sg13g2_fill_2 FILLER_6_1478 ();
 sg13g2_fill_2 FILLER_6_1530 ();
 sg13g2_fill_1 FILLER_6_1575 ();
 sg13g2_fill_2 FILLER_6_1613 ();
 sg13g2_fill_2 FILLER_6_1630 ();
 sg13g2_fill_1 FILLER_6_1632 ();
 sg13g2_fill_1 FILLER_6_1661 ();
 sg13g2_fill_2 FILLER_6_1675 ();
 sg13g2_fill_2 FILLER_6_1690 ();
 sg13g2_fill_2 FILLER_6_1730 ();
 sg13g2_fill_2 FILLER_6_1754 ();
 sg13g2_fill_1 FILLER_6_1756 ();
 sg13g2_fill_1 FILLER_6_1811 ();
 sg13g2_fill_1 FILLER_6_1864 ();
 sg13g2_decap_4 FILLER_6_1901 ();
 sg13g2_fill_1 FILLER_6_1905 ();
 sg13g2_decap_8 FILLER_6_1914 ();
 sg13g2_decap_4 FILLER_6_1949 ();
 sg13g2_fill_2 FILLER_6_1953 ();
 sg13g2_fill_2 FILLER_6_2006 ();
 sg13g2_fill_1 FILLER_6_2017 ();
 sg13g2_fill_1 FILLER_6_2055 ();
 sg13g2_fill_2 FILLER_6_2092 ();
 sg13g2_decap_8 FILLER_6_2130 ();
 sg13g2_decap_8 FILLER_6_2137 ();
 sg13g2_decap_8 FILLER_6_2144 ();
 sg13g2_fill_2 FILLER_6_2151 ();
 sg13g2_fill_1 FILLER_6_2153 ();
 sg13g2_decap_8 FILLER_6_2157 ();
 sg13g2_decap_8 FILLER_6_2164 ();
 sg13g2_decap_8 FILLER_6_2171 ();
 sg13g2_decap_8 FILLER_6_2178 ();
 sg13g2_decap_8 FILLER_6_2185 ();
 sg13g2_decap_8 FILLER_6_2192 ();
 sg13g2_decap_8 FILLER_6_2199 ();
 sg13g2_decap_8 FILLER_6_2206 ();
 sg13g2_decap_8 FILLER_6_2213 ();
 sg13g2_decap_8 FILLER_6_2220 ();
 sg13g2_decap_8 FILLER_6_2227 ();
 sg13g2_decap_8 FILLER_6_2234 ();
 sg13g2_decap_8 FILLER_6_2241 ();
 sg13g2_decap_8 FILLER_6_2248 ();
 sg13g2_decap_8 FILLER_6_2255 ();
 sg13g2_decap_8 FILLER_6_2262 ();
 sg13g2_decap_8 FILLER_6_2269 ();
 sg13g2_decap_8 FILLER_6_2276 ();
 sg13g2_decap_8 FILLER_6_2283 ();
 sg13g2_decap_8 FILLER_6_2290 ();
 sg13g2_decap_8 FILLER_6_2297 ();
 sg13g2_decap_8 FILLER_6_2304 ();
 sg13g2_decap_8 FILLER_6_2311 ();
 sg13g2_decap_8 FILLER_6_2318 ();
 sg13g2_decap_8 FILLER_6_2325 ();
 sg13g2_decap_8 FILLER_6_2332 ();
 sg13g2_decap_8 FILLER_6_2339 ();
 sg13g2_decap_8 FILLER_6_2346 ();
 sg13g2_decap_8 FILLER_6_2353 ();
 sg13g2_decap_8 FILLER_6_2360 ();
 sg13g2_decap_8 FILLER_6_2367 ();
 sg13g2_decap_8 FILLER_6_2374 ();
 sg13g2_decap_8 FILLER_6_2381 ();
 sg13g2_decap_8 FILLER_6_2388 ();
 sg13g2_decap_8 FILLER_6_2395 ();
 sg13g2_decap_8 FILLER_6_2402 ();
 sg13g2_decap_8 FILLER_6_2409 ();
 sg13g2_decap_8 FILLER_6_2416 ();
 sg13g2_decap_8 FILLER_6_2423 ();
 sg13g2_decap_8 FILLER_6_2430 ();
 sg13g2_decap_8 FILLER_6_2437 ();
 sg13g2_decap_8 FILLER_6_2444 ();
 sg13g2_decap_8 FILLER_6_2451 ();
 sg13g2_decap_8 FILLER_6_2458 ();
 sg13g2_decap_8 FILLER_6_2465 ();
 sg13g2_decap_8 FILLER_6_2472 ();
 sg13g2_decap_8 FILLER_6_2479 ();
 sg13g2_decap_8 FILLER_6_2486 ();
 sg13g2_decap_8 FILLER_6_2493 ();
 sg13g2_decap_8 FILLER_6_2500 ();
 sg13g2_decap_8 FILLER_6_2507 ();
 sg13g2_decap_8 FILLER_6_2514 ();
 sg13g2_decap_8 FILLER_6_2521 ();
 sg13g2_decap_8 FILLER_6_2528 ();
 sg13g2_decap_8 FILLER_6_2535 ();
 sg13g2_decap_8 FILLER_6_2542 ();
 sg13g2_decap_8 FILLER_6_2549 ();
 sg13g2_decap_8 FILLER_6_2556 ();
 sg13g2_decap_8 FILLER_6_2563 ();
 sg13g2_decap_8 FILLER_6_2570 ();
 sg13g2_decap_8 FILLER_6_2577 ();
 sg13g2_decap_8 FILLER_6_2584 ();
 sg13g2_decap_8 FILLER_6_2591 ();
 sg13g2_decap_8 FILLER_6_2598 ();
 sg13g2_decap_8 FILLER_6_2605 ();
 sg13g2_decap_8 FILLER_6_2612 ();
 sg13g2_decap_8 FILLER_6_2619 ();
 sg13g2_decap_8 FILLER_6_2626 ();
 sg13g2_decap_8 FILLER_6_2633 ();
 sg13g2_decap_8 FILLER_6_2640 ();
 sg13g2_decap_8 FILLER_6_2647 ();
 sg13g2_decap_8 FILLER_6_2654 ();
 sg13g2_decap_8 FILLER_6_2661 ();
 sg13g2_decap_4 FILLER_6_2668 ();
 sg13g2_fill_2 FILLER_6_2672 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_36 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_decap_8 FILLER_7_92 ();
 sg13g2_decap_8 FILLER_7_99 ();
 sg13g2_fill_2 FILLER_7_106 ();
 sg13g2_fill_2 FILLER_7_161 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_fill_1 FILLER_7_313 ();
 sg13g2_decap_4 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_430 ();
 sg13g2_fill_1 FILLER_7_432 ();
 sg13g2_fill_1 FILLER_7_451 ();
 sg13g2_fill_2 FILLER_7_488 ();
 sg13g2_fill_1 FILLER_7_490 ();
 sg13g2_fill_1 FILLER_7_541 ();
 sg13g2_decap_8 FILLER_7_547 ();
 sg13g2_decap_8 FILLER_7_554 ();
 sg13g2_decap_8 FILLER_7_561 ();
 sg13g2_fill_1 FILLER_7_568 ();
 sg13g2_fill_1 FILLER_7_587 ();
 sg13g2_decap_8 FILLER_7_607 ();
 sg13g2_decap_8 FILLER_7_614 ();
 sg13g2_fill_2 FILLER_7_651 ();
 sg13g2_fill_1 FILLER_7_653 ();
 sg13g2_decap_8 FILLER_7_663 ();
 sg13g2_fill_2 FILLER_7_681 ();
 sg13g2_fill_1 FILLER_7_683 ();
 sg13g2_fill_1 FILLER_7_694 ();
 sg13g2_fill_2 FILLER_7_710 ();
 sg13g2_fill_1 FILLER_7_722 ();
 sg13g2_fill_1 FILLER_7_805 ();
 sg13g2_fill_1 FILLER_7_837 ();
 sg13g2_fill_1 FILLER_7_925 ();
 sg13g2_decap_8 FILLER_7_954 ();
 sg13g2_decap_8 FILLER_7_961 ();
 sg13g2_decap_8 FILLER_7_999 ();
 sg13g2_decap_8 FILLER_7_1006 ();
 sg13g2_decap_4 FILLER_7_1013 ();
 sg13g2_fill_2 FILLER_7_1017 ();
 sg13g2_fill_1 FILLER_7_1043 ();
 sg13g2_decap_8 FILLER_7_1048 ();
 sg13g2_decap_4 FILLER_7_1055 ();
 sg13g2_fill_1 FILLER_7_1059 ();
 sg13g2_decap_8 FILLER_7_1072 ();
 sg13g2_fill_1 FILLER_7_1079 ();
 sg13g2_fill_1 FILLER_7_1103 ();
 sg13g2_fill_2 FILLER_7_1120 ();
 sg13g2_fill_2 FILLER_7_1128 ();
 sg13g2_fill_1 FILLER_7_1130 ();
 sg13g2_fill_1 FILLER_7_1159 ();
 sg13g2_decap_4 FILLER_7_1214 ();
 sg13g2_fill_1 FILLER_7_1218 ();
 sg13g2_fill_2 FILLER_7_1228 ();
 sg13g2_decap_4 FILLER_7_1311 ();
 sg13g2_fill_1 FILLER_7_1324 ();
 sg13g2_fill_1 FILLER_7_1381 ();
 sg13g2_fill_1 FILLER_7_1433 ();
 sg13g2_fill_1 FILLER_7_1482 ();
 sg13g2_fill_2 FILLER_7_1695 ();
 sg13g2_fill_1 FILLER_7_1762 ();
 sg13g2_fill_1 FILLER_7_1785 ();
 sg13g2_fill_2 FILLER_7_1820 ();
 sg13g2_fill_2 FILLER_7_1849 ();
 sg13g2_fill_2 FILLER_7_1887 ();
 sg13g2_fill_1 FILLER_7_1982 ();
 sg13g2_fill_1 FILLER_7_2017 ();
 sg13g2_fill_2 FILLER_7_2050 ();
 sg13g2_decap_8 FILLER_7_2166 ();
 sg13g2_decap_8 FILLER_7_2173 ();
 sg13g2_decap_8 FILLER_7_2180 ();
 sg13g2_decap_8 FILLER_7_2187 ();
 sg13g2_decap_8 FILLER_7_2194 ();
 sg13g2_decap_8 FILLER_7_2201 ();
 sg13g2_decap_8 FILLER_7_2208 ();
 sg13g2_decap_8 FILLER_7_2215 ();
 sg13g2_decap_8 FILLER_7_2222 ();
 sg13g2_decap_8 FILLER_7_2229 ();
 sg13g2_decap_8 FILLER_7_2236 ();
 sg13g2_decap_8 FILLER_7_2243 ();
 sg13g2_decap_8 FILLER_7_2250 ();
 sg13g2_decap_8 FILLER_7_2257 ();
 sg13g2_decap_8 FILLER_7_2264 ();
 sg13g2_decap_8 FILLER_7_2271 ();
 sg13g2_decap_8 FILLER_7_2278 ();
 sg13g2_decap_8 FILLER_7_2285 ();
 sg13g2_decap_8 FILLER_7_2292 ();
 sg13g2_decap_8 FILLER_7_2299 ();
 sg13g2_decap_8 FILLER_7_2306 ();
 sg13g2_decap_8 FILLER_7_2313 ();
 sg13g2_decap_8 FILLER_7_2320 ();
 sg13g2_decap_8 FILLER_7_2327 ();
 sg13g2_decap_8 FILLER_7_2334 ();
 sg13g2_decap_8 FILLER_7_2341 ();
 sg13g2_decap_8 FILLER_7_2348 ();
 sg13g2_decap_8 FILLER_7_2355 ();
 sg13g2_decap_8 FILLER_7_2362 ();
 sg13g2_decap_8 FILLER_7_2369 ();
 sg13g2_decap_8 FILLER_7_2376 ();
 sg13g2_decap_8 FILLER_7_2383 ();
 sg13g2_decap_8 FILLER_7_2390 ();
 sg13g2_decap_8 FILLER_7_2397 ();
 sg13g2_decap_8 FILLER_7_2404 ();
 sg13g2_decap_8 FILLER_7_2411 ();
 sg13g2_decap_8 FILLER_7_2418 ();
 sg13g2_decap_8 FILLER_7_2425 ();
 sg13g2_decap_8 FILLER_7_2432 ();
 sg13g2_decap_8 FILLER_7_2439 ();
 sg13g2_decap_8 FILLER_7_2446 ();
 sg13g2_decap_8 FILLER_7_2453 ();
 sg13g2_decap_8 FILLER_7_2460 ();
 sg13g2_decap_8 FILLER_7_2467 ();
 sg13g2_decap_8 FILLER_7_2474 ();
 sg13g2_decap_8 FILLER_7_2481 ();
 sg13g2_decap_8 FILLER_7_2488 ();
 sg13g2_decap_8 FILLER_7_2495 ();
 sg13g2_decap_8 FILLER_7_2502 ();
 sg13g2_decap_8 FILLER_7_2509 ();
 sg13g2_decap_8 FILLER_7_2516 ();
 sg13g2_decap_8 FILLER_7_2523 ();
 sg13g2_decap_8 FILLER_7_2530 ();
 sg13g2_decap_8 FILLER_7_2537 ();
 sg13g2_decap_8 FILLER_7_2544 ();
 sg13g2_decap_8 FILLER_7_2551 ();
 sg13g2_decap_8 FILLER_7_2558 ();
 sg13g2_decap_8 FILLER_7_2565 ();
 sg13g2_decap_8 FILLER_7_2572 ();
 sg13g2_decap_8 FILLER_7_2579 ();
 sg13g2_decap_8 FILLER_7_2586 ();
 sg13g2_decap_8 FILLER_7_2593 ();
 sg13g2_decap_8 FILLER_7_2600 ();
 sg13g2_decap_8 FILLER_7_2607 ();
 sg13g2_decap_8 FILLER_7_2614 ();
 sg13g2_decap_8 FILLER_7_2621 ();
 sg13g2_decap_8 FILLER_7_2628 ();
 sg13g2_decap_8 FILLER_7_2635 ();
 sg13g2_decap_8 FILLER_7_2642 ();
 sg13g2_decap_8 FILLER_7_2649 ();
 sg13g2_decap_8 FILLER_7_2656 ();
 sg13g2_decap_8 FILLER_7_2663 ();
 sg13g2_decap_4 FILLER_7_2670 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_32 ();
 sg13g2_fill_2 FILLER_8_51 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_fill_1 FILLER_8_69 ();
 sg13g2_decap_8 FILLER_8_101 ();
 sg13g2_fill_2 FILLER_8_108 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_125 ();
 sg13g2_decap_8 FILLER_8_187 ();
 sg13g2_decap_4 FILLER_8_194 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_decap_4 FILLER_8_204 ();
 sg13g2_decap_4 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_269 ();
 sg13g2_fill_1 FILLER_8_271 ();
 sg13g2_fill_2 FILLER_8_281 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_2 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_432 ();
 sg13g2_fill_1 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_478 ();
 sg13g2_decap_8 FILLER_8_485 ();
 sg13g2_fill_1 FILLER_8_492 ();
 sg13g2_decap_8 FILLER_8_568 ();
 sg13g2_fill_1 FILLER_8_575 ();
 sg13g2_fill_1 FILLER_8_594 ();
 sg13g2_decap_8 FILLER_8_605 ();
 sg13g2_decap_8 FILLER_8_612 ();
 sg13g2_fill_2 FILLER_8_619 ();
 sg13g2_fill_1 FILLER_8_621 ();
 sg13g2_fill_2 FILLER_8_653 ();
 sg13g2_decap_4 FILLER_8_670 ();
 sg13g2_fill_1 FILLER_8_684 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_4 FILLER_8_712 ();
 sg13g2_fill_2 FILLER_8_775 ();
 sg13g2_decap_4 FILLER_8_781 ();
 sg13g2_fill_1 FILLER_8_807 ();
 sg13g2_fill_2 FILLER_8_836 ();
 sg13g2_fill_2 FILLER_8_887 ();
 sg13g2_fill_2 FILLER_8_935 ();
 sg13g2_decap_8 FILLER_8_965 ();
 sg13g2_fill_2 FILLER_8_972 ();
 sg13g2_fill_2 FILLER_8_984 ();
 sg13g2_fill_2 FILLER_8_995 ();
 sg13g2_fill_1 FILLER_8_997 ();
 sg13g2_decap_8 FILLER_8_1002 ();
 sg13g2_decap_8 FILLER_8_1009 ();
 sg13g2_decap_8 FILLER_8_1016 ();
 sg13g2_decap_8 FILLER_8_1033 ();
 sg13g2_decap_8 FILLER_8_1040 ();
 sg13g2_decap_8 FILLER_8_1047 ();
 sg13g2_fill_1 FILLER_8_1054 ();
 sg13g2_decap_8 FILLER_8_1059 ();
 sg13g2_decap_8 FILLER_8_1066 ();
 sg13g2_decap_8 FILLER_8_1073 ();
 sg13g2_decap_4 FILLER_8_1080 ();
 sg13g2_fill_1 FILLER_8_1138 ();
 sg13g2_fill_1 FILLER_8_1270 ();
 sg13g2_fill_2 FILLER_8_1307 ();
 sg13g2_fill_1 FILLER_8_1309 ();
 sg13g2_decap_8 FILLER_8_1315 ();
 sg13g2_fill_2 FILLER_8_1322 ();
 sg13g2_fill_2 FILLER_8_1397 ();
 sg13g2_fill_1 FILLER_8_1399 ();
 sg13g2_fill_2 FILLER_8_1408 ();
 sg13g2_fill_1 FILLER_8_1410 ();
 sg13g2_decap_8 FILLER_8_1429 ();
 sg13g2_fill_2 FILLER_8_1436 ();
 sg13g2_fill_1 FILLER_8_1438 ();
 sg13g2_fill_1 FILLER_8_1460 ();
 sg13g2_fill_2 FILLER_8_1470 ();
 sg13g2_fill_2 FILLER_8_1507 ();
 sg13g2_fill_1 FILLER_8_1523 ();
 sg13g2_fill_1 FILLER_8_1577 ();
 sg13g2_decap_4 FILLER_8_1676 ();
 sg13g2_fill_2 FILLER_8_1763 ();
 sg13g2_fill_2 FILLER_8_1792 ();
 sg13g2_fill_1 FILLER_8_1794 ();
 sg13g2_decap_4 FILLER_8_1804 ();
 sg13g2_fill_2 FILLER_8_1817 ();
 sg13g2_fill_1 FILLER_8_1846 ();
 sg13g2_fill_2 FILLER_8_1875 ();
 sg13g2_fill_2 FILLER_8_1910 ();
 sg13g2_fill_2 FILLER_8_1953 ();
 sg13g2_fill_1 FILLER_8_1955 ();
 sg13g2_fill_2 FILLER_8_1988 ();
 sg13g2_fill_1 FILLER_8_1990 ();
 sg13g2_fill_2 FILLER_8_2019 ();
 sg13g2_fill_2 FILLER_8_2064 ();
 sg13g2_fill_2 FILLER_8_2085 ();
 sg13g2_fill_2 FILLER_8_2101 ();
 sg13g2_fill_1 FILLER_8_2143 ();
 sg13g2_decap_8 FILLER_8_2172 ();
 sg13g2_decap_8 FILLER_8_2179 ();
 sg13g2_decap_8 FILLER_8_2186 ();
 sg13g2_decap_8 FILLER_8_2193 ();
 sg13g2_decap_8 FILLER_8_2200 ();
 sg13g2_decap_8 FILLER_8_2207 ();
 sg13g2_decap_8 FILLER_8_2214 ();
 sg13g2_decap_8 FILLER_8_2221 ();
 sg13g2_decap_8 FILLER_8_2228 ();
 sg13g2_decap_8 FILLER_8_2235 ();
 sg13g2_decap_8 FILLER_8_2242 ();
 sg13g2_decap_8 FILLER_8_2249 ();
 sg13g2_decap_8 FILLER_8_2256 ();
 sg13g2_decap_8 FILLER_8_2263 ();
 sg13g2_decap_8 FILLER_8_2270 ();
 sg13g2_decap_8 FILLER_8_2277 ();
 sg13g2_decap_8 FILLER_8_2284 ();
 sg13g2_decap_8 FILLER_8_2291 ();
 sg13g2_decap_8 FILLER_8_2298 ();
 sg13g2_decap_8 FILLER_8_2305 ();
 sg13g2_decap_8 FILLER_8_2312 ();
 sg13g2_decap_8 FILLER_8_2319 ();
 sg13g2_decap_8 FILLER_8_2326 ();
 sg13g2_decap_8 FILLER_8_2333 ();
 sg13g2_decap_8 FILLER_8_2340 ();
 sg13g2_decap_8 FILLER_8_2347 ();
 sg13g2_decap_8 FILLER_8_2354 ();
 sg13g2_decap_8 FILLER_8_2361 ();
 sg13g2_decap_8 FILLER_8_2368 ();
 sg13g2_decap_8 FILLER_8_2375 ();
 sg13g2_decap_8 FILLER_8_2382 ();
 sg13g2_decap_8 FILLER_8_2389 ();
 sg13g2_decap_8 FILLER_8_2396 ();
 sg13g2_decap_8 FILLER_8_2403 ();
 sg13g2_decap_8 FILLER_8_2410 ();
 sg13g2_decap_8 FILLER_8_2417 ();
 sg13g2_decap_8 FILLER_8_2424 ();
 sg13g2_decap_8 FILLER_8_2431 ();
 sg13g2_decap_8 FILLER_8_2438 ();
 sg13g2_decap_8 FILLER_8_2445 ();
 sg13g2_decap_8 FILLER_8_2452 ();
 sg13g2_decap_8 FILLER_8_2459 ();
 sg13g2_decap_8 FILLER_8_2466 ();
 sg13g2_decap_8 FILLER_8_2473 ();
 sg13g2_decap_8 FILLER_8_2480 ();
 sg13g2_decap_8 FILLER_8_2487 ();
 sg13g2_decap_8 FILLER_8_2494 ();
 sg13g2_decap_8 FILLER_8_2501 ();
 sg13g2_decap_8 FILLER_8_2508 ();
 sg13g2_decap_8 FILLER_8_2515 ();
 sg13g2_decap_8 FILLER_8_2522 ();
 sg13g2_decap_8 FILLER_8_2529 ();
 sg13g2_decap_8 FILLER_8_2536 ();
 sg13g2_decap_8 FILLER_8_2543 ();
 sg13g2_decap_8 FILLER_8_2550 ();
 sg13g2_decap_8 FILLER_8_2557 ();
 sg13g2_decap_8 FILLER_8_2564 ();
 sg13g2_decap_8 FILLER_8_2571 ();
 sg13g2_decap_8 FILLER_8_2578 ();
 sg13g2_decap_8 FILLER_8_2585 ();
 sg13g2_decap_8 FILLER_8_2592 ();
 sg13g2_decap_8 FILLER_8_2599 ();
 sg13g2_decap_8 FILLER_8_2606 ();
 sg13g2_decap_8 FILLER_8_2613 ();
 sg13g2_decap_8 FILLER_8_2620 ();
 sg13g2_decap_8 FILLER_8_2627 ();
 sg13g2_decap_8 FILLER_8_2634 ();
 sg13g2_decap_8 FILLER_8_2641 ();
 sg13g2_decap_8 FILLER_8_2648 ();
 sg13g2_decap_8 FILLER_8_2655 ();
 sg13g2_decap_8 FILLER_8_2662 ();
 sg13g2_decap_4 FILLER_8_2669 ();
 sg13g2_fill_1 FILLER_8_2673 ();
 sg13g2_fill_2 FILLER_9_41 ();
 sg13g2_fill_1 FILLER_9_43 ();
 sg13g2_fill_1 FILLER_9_71 ();
 sg13g2_fill_2 FILLER_9_94 ();
 sg13g2_fill_1 FILLER_9_96 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_decap_4 FILLER_9_197 ();
 sg13g2_fill_1 FILLER_9_201 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_fill_2 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_4 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_298 ();
 sg13g2_fill_2 FILLER_9_309 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_365 ();
 sg13g2_fill_1 FILLER_9_367 ();
 sg13g2_fill_2 FILLER_9_424 ();
 sg13g2_fill_1 FILLER_9_426 ();
 sg13g2_fill_2 FILLER_9_454 ();
 sg13g2_fill_1 FILLER_9_456 ();
 sg13g2_decap_8 FILLER_9_474 ();
 sg13g2_decap_8 FILLER_9_481 ();
 sg13g2_decap_8 FILLER_9_488 ();
 sg13g2_fill_1 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_526 ();
 sg13g2_decap_8 FILLER_9_533 ();
 sg13g2_decap_8 FILLER_9_540 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_4 FILLER_9_574 ();
 sg13g2_fill_1 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_608 ();
 sg13g2_decap_8 FILLER_9_615 ();
 sg13g2_decap_4 FILLER_9_622 ();
 sg13g2_fill_1 FILLER_9_626 ();
 sg13g2_fill_1 FILLER_9_677 ();
 sg13g2_fill_1 FILLER_9_690 ();
 sg13g2_decap_8 FILLER_9_708 ();
 sg13g2_decap_8 FILLER_9_715 ();
 sg13g2_fill_2 FILLER_9_722 ();
 sg13g2_fill_1 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_768 ();
 sg13g2_decap_8 FILLER_9_775 ();
 sg13g2_fill_2 FILLER_9_782 ();
 sg13g2_fill_1 FILLER_9_858 ();
 sg13g2_fill_2 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_888 ();
 sg13g2_fill_2 FILLER_9_904 ();
 sg13g2_fill_1 FILLER_9_906 ();
 sg13g2_fill_2 FILLER_9_921 ();
 sg13g2_decap_8 FILLER_9_967 ();
 sg13g2_decap_4 FILLER_9_974 ();
 sg13g2_fill_1 FILLER_9_978 ();
 sg13g2_decap_8 FILLER_9_1012 ();
 sg13g2_decap_8 FILLER_9_1019 ();
 sg13g2_decap_8 FILLER_9_1026 ();
 sg13g2_decap_8 FILLER_9_1033 ();
 sg13g2_decap_8 FILLER_9_1040 ();
 sg13g2_decap_4 FILLER_9_1047 ();
 sg13g2_decap_8 FILLER_9_1069 ();
 sg13g2_decap_8 FILLER_9_1076 ();
 sg13g2_decap_4 FILLER_9_1083 ();
 sg13g2_fill_1 FILLER_9_1134 ();
 sg13g2_fill_2 FILLER_9_1298 ();
 sg13g2_fill_1 FILLER_9_1300 ();
 sg13g2_fill_1 FILLER_9_1313 ();
 sg13g2_fill_2 FILLER_9_1319 ();
 sg13g2_decap_4 FILLER_9_1325 ();
 sg13g2_fill_2 FILLER_9_1329 ();
 sg13g2_fill_1 FILLER_9_1348 ();
 sg13g2_fill_1 FILLER_9_1433 ();
 sg13g2_fill_2 FILLER_9_1444 ();
 sg13g2_decap_8 FILLER_9_1463 ();
 sg13g2_decap_4 FILLER_9_1470 ();
 sg13g2_fill_2 FILLER_9_1474 ();
 sg13g2_fill_2 FILLER_9_1535 ();
 sg13g2_fill_2 FILLER_9_1602 ();
 sg13g2_fill_2 FILLER_9_1631 ();
 sg13g2_fill_1 FILLER_9_1633 ();
 sg13g2_fill_2 FILLER_9_1701 ();
 sg13g2_fill_1 FILLER_9_1703 ();
 sg13g2_fill_2 FILLER_9_1760 ();
 sg13g2_fill_1 FILLER_9_1762 ();
 sg13g2_fill_2 FILLER_9_1790 ();
 sg13g2_fill_1 FILLER_9_1947 ();
 sg13g2_fill_1 FILLER_9_1970 ();
 sg13g2_fill_1 FILLER_9_2045 ();
 sg13g2_fill_2 FILLER_9_2122 ();
 sg13g2_fill_1 FILLER_9_2124 ();
 sg13g2_decap_8 FILLER_9_2183 ();
 sg13g2_decap_8 FILLER_9_2190 ();
 sg13g2_decap_8 FILLER_9_2197 ();
 sg13g2_decap_8 FILLER_9_2204 ();
 sg13g2_decap_8 FILLER_9_2211 ();
 sg13g2_decap_8 FILLER_9_2218 ();
 sg13g2_decap_8 FILLER_9_2225 ();
 sg13g2_decap_8 FILLER_9_2232 ();
 sg13g2_decap_8 FILLER_9_2239 ();
 sg13g2_decap_8 FILLER_9_2246 ();
 sg13g2_decap_8 FILLER_9_2253 ();
 sg13g2_decap_8 FILLER_9_2260 ();
 sg13g2_decap_8 FILLER_9_2267 ();
 sg13g2_decap_8 FILLER_9_2274 ();
 sg13g2_decap_8 FILLER_9_2281 ();
 sg13g2_decap_8 FILLER_9_2288 ();
 sg13g2_decap_8 FILLER_9_2295 ();
 sg13g2_decap_8 FILLER_9_2302 ();
 sg13g2_decap_8 FILLER_9_2309 ();
 sg13g2_decap_8 FILLER_9_2316 ();
 sg13g2_decap_8 FILLER_9_2323 ();
 sg13g2_decap_8 FILLER_9_2330 ();
 sg13g2_decap_8 FILLER_9_2337 ();
 sg13g2_decap_8 FILLER_9_2344 ();
 sg13g2_decap_8 FILLER_9_2351 ();
 sg13g2_decap_8 FILLER_9_2358 ();
 sg13g2_decap_8 FILLER_9_2365 ();
 sg13g2_decap_8 FILLER_9_2372 ();
 sg13g2_decap_8 FILLER_9_2379 ();
 sg13g2_decap_8 FILLER_9_2386 ();
 sg13g2_decap_8 FILLER_9_2393 ();
 sg13g2_decap_8 FILLER_9_2400 ();
 sg13g2_decap_8 FILLER_9_2407 ();
 sg13g2_decap_8 FILLER_9_2414 ();
 sg13g2_decap_8 FILLER_9_2421 ();
 sg13g2_decap_8 FILLER_9_2428 ();
 sg13g2_decap_8 FILLER_9_2435 ();
 sg13g2_decap_8 FILLER_9_2442 ();
 sg13g2_decap_8 FILLER_9_2449 ();
 sg13g2_decap_8 FILLER_9_2456 ();
 sg13g2_decap_8 FILLER_9_2463 ();
 sg13g2_decap_8 FILLER_9_2470 ();
 sg13g2_decap_8 FILLER_9_2477 ();
 sg13g2_decap_8 FILLER_9_2484 ();
 sg13g2_decap_8 FILLER_9_2491 ();
 sg13g2_decap_8 FILLER_9_2498 ();
 sg13g2_decap_8 FILLER_9_2505 ();
 sg13g2_decap_8 FILLER_9_2512 ();
 sg13g2_decap_8 FILLER_9_2519 ();
 sg13g2_decap_8 FILLER_9_2526 ();
 sg13g2_decap_8 FILLER_9_2533 ();
 sg13g2_decap_8 FILLER_9_2540 ();
 sg13g2_decap_8 FILLER_9_2547 ();
 sg13g2_decap_8 FILLER_9_2554 ();
 sg13g2_decap_8 FILLER_9_2561 ();
 sg13g2_decap_8 FILLER_9_2568 ();
 sg13g2_decap_8 FILLER_9_2575 ();
 sg13g2_decap_8 FILLER_9_2582 ();
 sg13g2_decap_8 FILLER_9_2589 ();
 sg13g2_decap_8 FILLER_9_2596 ();
 sg13g2_decap_8 FILLER_9_2603 ();
 sg13g2_decap_8 FILLER_9_2610 ();
 sg13g2_decap_8 FILLER_9_2617 ();
 sg13g2_decap_8 FILLER_9_2624 ();
 sg13g2_decap_8 FILLER_9_2631 ();
 sg13g2_decap_8 FILLER_9_2638 ();
 sg13g2_decap_8 FILLER_9_2645 ();
 sg13g2_decap_8 FILLER_9_2652 ();
 sg13g2_decap_8 FILLER_9_2659 ();
 sg13g2_decap_8 FILLER_9_2666 ();
 sg13g2_fill_1 FILLER_9_2673 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_66 ();
 sg13g2_fill_2 FILLER_10_79 ();
 sg13g2_decap_4 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_177 ();
 sg13g2_fill_2 FILLER_10_192 ();
 sg13g2_fill_1 FILLER_10_194 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_fill_2 FILLER_10_267 ();
 sg13g2_fill_2 FILLER_10_283 ();
 sg13g2_decap_4 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_313 ();
 sg13g2_fill_2 FILLER_10_354 ();
 sg13g2_decap_4 FILLER_10_456 ();
 sg13g2_fill_1 FILLER_10_460 ();
 sg13g2_decap_8 FILLER_10_470 ();
 sg13g2_decap_8 FILLER_10_477 ();
 sg13g2_decap_8 FILLER_10_484 ();
 sg13g2_fill_1 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_fill_2 FILLER_10_539 ();
 sg13g2_fill_1 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_fill_1 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_612 ();
 sg13g2_decap_8 FILLER_10_619 ();
 sg13g2_decap_8 FILLER_10_626 ();
 sg13g2_fill_2 FILLER_10_633 ();
 sg13g2_fill_1 FILLER_10_635 ();
 sg13g2_fill_2 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_655 ();
 sg13g2_fill_1 FILLER_10_657 ();
 sg13g2_decap_4 FILLER_10_663 ();
 sg13g2_decap_4 FILLER_10_682 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_fill_2 FILLER_10_728 ();
 sg13g2_fill_1 FILLER_10_730 ();
 sg13g2_fill_2 FILLER_10_748 ();
 sg13g2_fill_1 FILLER_10_750 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_776 ();
 sg13g2_decap_4 FILLER_10_783 ();
 sg13g2_fill_1 FILLER_10_787 ();
 sg13g2_decap_4 FILLER_10_865 ();
 sg13g2_fill_2 FILLER_10_869 ();
 sg13g2_fill_2 FILLER_10_874 ();
 sg13g2_fill_1 FILLER_10_876 ();
 sg13g2_fill_1 FILLER_10_880 ();
 sg13g2_fill_2 FILLER_10_932 ();
 sg13g2_fill_2 FILLER_10_952 ();
 sg13g2_decap_8 FILLER_10_967 ();
 sg13g2_decap_4 FILLER_10_974 ();
 sg13g2_fill_1 FILLER_10_978 ();
 sg13g2_decap_8 FILLER_10_1023 ();
 sg13g2_decap_8 FILLER_10_1030 ();
 sg13g2_decap_8 FILLER_10_1037 ();
 sg13g2_fill_1 FILLER_10_1044 ();
 sg13g2_fill_2 FILLER_10_1064 ();
 sg13g2_fill_2 FILLER_10_1082 ();
 sg13g2_fill_1 FILLER_10_1084 ();
 sg13g2_fill_1 FILLER_10_1174 ();
 sg13g2_decap_4 FILLER_10_1211 ();
 sg13g2_decap_8 FILLER_10_1224 ();
 sg13g2_fill_2 FILLER_10_1235 ();
 sg13g2_fill_1 FILLER_10_1277 ();
 sg13g2_fill_2 FILLER_10_1295 ();
 sg13g2_fill_2 FILLER_10_1325 ();
 sg13g2_fill_1 FILLER_10_1327 ();
 sg13g2_fill_1 FILLER_10_1334 ();
 sg13g2_fill_1 FILLER_10_1340 ();
 sg13g2_fill_2 FILLER_10_1400 ();
 sg13g2_fill_1 FILLER_10_1402 ();
 sg13g2_fill_2 FILLER_10_1426 ();
 sg13g2_fill_2 FILLER_10_1450 ();
 sg13g2_decap_4 FILLER_10_1471 ();
 sg13g2_fill_2 FILLER_10_1546 ();
 sg13g2_fill_1 FILLER_10_1650 ();
 sg13g2_fill_1 FILLER_10_1692 ();
 sg13g2_fill_2 FILLER_10_1707 ();
 sg13g2_fill_2 FILLER_10_1715 ();
 sg13g2_fill_1 FILLER_10_1730 ();
 sg13g2_fill_1 FILLER_10_1758 ();
 sg13g2_fill_2 FILLER_10_1771 ();
 sg13g2_fill_1 FILLER_10_1773 ();
 sg13g2_decap_4 FILLER_10_1783 ();
 sg13g2_fill_2 FILLER_10_1836 ();
 sg13g2_fill_1 FILLER_10_1838 ();
 sg13g2_fill_2 FILLER_10_1896 ();
 sg13g2_fill_1 FILLER_10_1907 ();
 sg13g2_decap_4 FILLER_10_1945 ();
 sg13g2_fill_1 FILLER_10_2028 ();
 sg13g2_fill_2 FILLER_10_2068 ();
 sg13g2_fill_1 FILLER_10_2070 ();
 sg13g2_fill_1 FILLER_10_2102 ();
 sg13g2_fill_2 FILLER_10_2121 ();
 sg13g2_fill_2 FILLER_10_2129 ();
 sg13g2_fill_2 FILLER_10_2158 ();
 sg13g2_decap_8 FILLER_10_2178 ();
 sg13g2_decap_8 FILLER_10_2185 ();
 sg13g2_decap_8 FILLER_10_2192 ();
 sg13g2_decap_8 FILLER_10_2199 ();
 sg13g2_decap_8 FILLER_10_2206 ();
 sg13g2_decap_8 FILLER_10_2213 ();
 sg13g2_decap_8 FILLER_10_2220 ();
 sg13g2_decap_8 FILLER_10_2227 ();
 sg13g2_decap_8 FILLER_10_2234 ();
 sg13g2_decap_8 FILLER_10_2241 ();
 sg13g2_decap_8 FILLER_10_2248 ();
 sg13g2_decap_8 FILLER_10_2255 ();
 sg13g2_decap_8 FILLER_10_2262 ();
 sg13g2_decap_8 FILLER_10_2269 ();
 sg13g2_decap_8 FILLER_10_2276 ();
 sg13g2_decap_8 FILLER_10_2283 ();
 sg13g2_decap_8 FILLER_10_2290 ();
 sg13g2_decap_8 FILLER_10_2297 ();
 sg13g2_decap_8 FILLER_10_2304 ();
 sg13g2_decap_8 FILLER_10_2311 ();
 sg13g2_decap_8 FILLER_10_2318 ();
 sg13g2_decap_8 FILLER_10_2325 ();
 sg13g2_decap_8 FILLER_10_2332 ();
 sg13g2_decap_8 FILLER_10_2339 ();
 sg13g2_decap_8 FILLER_10_2346 ();
 sg13g2_decap_8 FILLER_10_2353 ();
 sg13g2_decap_8 FILLER_10_2360 ();
 sg13g2_decap_8 FILLER_10_2367 ();
 sg13g2_decap_8 FILLER_10_2374 ();
 sg13g2_decap_8 FILLER_10_2381 ();
 sg13g2_decap_8 FILLER_10_2388 ();
 sg13g2_decap_8 FILLER_10_2395 ();
 sg13g2_decap_8 FILLER_10_2402 ();
 sg13g2_decap_8 FILLER_10_2409 ();
 sg13g2_decap_8 FILLER_10_2416 ();
 sg13g2_decap_8 FILLER_10_2423 ();
 sg13g2_decap_8 FILLER_10_2430 ();
 sg13g2_decap_8 FILLER_10_2437 ();
 sg13g2_decap_8 FILLER_10_2444 ();
 sg13g2_decap_8 FILLER_10_2451 ();
 sg13g2_decap_8 FILLER_10_2458 ();
 sg13g2_decap_8 FILLER_10_2465 ();
 sg13g2_decap_8 FILLER_10_2472 ();
 sg13g2_decap_8 FILLER_10_2479 ();
 sg13g2_decap_8 FILLER_10_2486 ();
 sg13g2_decap_8 FILLER_10_2493 ();
 sg13g2_decap_8 FILLER_10_2500 ();
 sg13g2_decap_8 FILLER_10_2507 ();
 sg13g2_decap_8 FILLER_10_2514 ();
 sg13g2_decap_8 FILLER_10_2521 ();
 sg13g2_decap_8 FILLER_10_2528 ();
 sg13g2_decap_8 FILLER_10_2535 ();
 sg13g2_decap_8 FILLER_10_2542 ();
 sg13g2_decap_8 FILLER_10_2549 ();
 sg13g2_decap_8 FILLER_10_2556 ();
 sg13g2_decap_8 FILLER_10_2563 ();
 sg13g2_decap_8 FILLER_10_2570 ();
 sg13g2_decap_8 FILLER_10_2577 ();
 sg13g2_decap_8 FILLER_10_2584 ();
 sg13g2_decap_8 FILLER_10_2591 ();
 sg13g2_decap_8 FILLER_10_2598 ();
 sg13g2_decap_8 FILLER_10_2605 ();
 sg13g2_decap_8 FILLER_10_2612 ();
 sg13g2_decap_8 FILLER_10_2619 ();
 sg13g2_decap_8 FILLER_10_2626 ();
 sg13g2_decap_8 FILLER_10_2633 ();
 sg13g2_decap_8 FILLER_10_2640 ();
 sg13g2_decap_8 FILLER_10_2647 ();
 sg13g2_decap_8 FILLER_10_2654 ();
 sg13g2_decap_8 FILLER_10_2661 ();
 sg13g2_decap_4 FILLER_10_2668 ();
 sg13g2_fill_2 FILLER_10_2672 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_2 FILLER_11_85 ();
 sg13g2_fill_2 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_140 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_256 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_decap_4 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_2 FILLER_11_379 ();
 sg13g2_fill_2 FILLER_11_391 ();
 sg13g2_fill_2 FILLER_11_414 ();
 sg13g2_fill_2 FILLER_11_469 ();
 sg13g2_decap_4 FILLER_11_484 ();
 sg13g2_fill_1 FILLER_11_488 ();
 sg13g2_fill_2 FILLER_11_519 ();
 sg13g2_fill_2 FILLER_11_533 ();
 sg13g2_decap_8 FILLER_11_555 ();
 sg13g2_fill_1 FILLER_11_562 ();
 sg13g2_decap_4 FILLER_11_571 ();
 sg13g2_fill_2 FILLER_11_575 ();
 sg13g2_decap_4 FILLER_11_587 ();
 sg13g2_fill_2 FILLER_11_591 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_fill_1 FILLER_11_669 ();
 sg13g2_fill_2 FILLER_11_675 ();
 sg13g2_decap_8 FILLER_11_688 ();
 sg13g2_decap_8 FILLER_11_695 ();
 sg13g2_decap_8 FILLER_11_702 ();
 sg13g2_decap_8 FILLER_11_709 ();
 sg13g2_fill_2 FILLER_11_716 ();
 sg13g2_fill_1 FILLER_11_718 ();
 sg13g2_fill_2 FILLER_11_744 ();
 sg13g2_fill_1 FILLER_11_746 ();
 sg13g2_decap_4 FILLER_11_752 ();
 sg13g2_fill_1 FILLER_11_756 ();
 sg13g2_fill_1 FILLER_11_761 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_4 FILLER_11_849 ();
 sg13g2_fill_1 FILLER_11_853 ();
 sg13g2_fill_2 FILLER_11_885 ();
 sg13g2_fill_1 FILLER_11_887 ();
 sg13g2_fill_2 FILLER_11_938 ();
 sg13g2_fill_1 FILLER_11_943 ();
 sg13g2_fill_2 FILLER_11_957 ();
 sg13g2_decap_8 FILLER_11_972 ();
 sg13g2_decap_8 FILLER_11_979 ();
 sg13g2_fill_1 FILLER_11_986 ();
 sg13g2_decap_8 FILLER_11_1023 ();
 sg13g2_decap_8 FILLER_11_1030 ();
 sg13g2_decap_4 FILLER_11_1037 ();
 sg13g2_decap_8 FILLER_11_1072 ();
 sg13g2_decap_8 FILLER_11_1079 ();
 sg13g2_decap_8 FILLER_11_1086 ();
 sg13g2_fill_2 FILLER_11_1093 ();
 sg13g2_fill_1 FILLER_11_1095 ();
 sg13g2_decap_4 FILLER_11_1105 ();
 sg13g2_fill_2 FILLER_11_1109 ();
 sg13g2_fill_2 FILLER_11_1117 ();
 sg13g2_fill_1 FILLER_11_1119 ();
 sg13g2_fill_1 FILLER_11_1129 ();
 sg13g2_fill_2 FILLER_11_1172 ();
 sg13g2_decap_8 FILLER_11_1250 ();
 sg13g2_decap_4 FILLER_11_1257 ();
 sg13g2_fill_2 FILLER_11_1270 ();
 sg13g2_decap_8 FILLER_11_1347 ();
 sg13g2_fill_1 FILLER_11_1354 ();
 sg13g2_fill_1 FILLER_11_1388 ();
 sg13g2_fill_1 FILLER_11_1433 ();
 sg13g2_fill_1 FILLER_11_1493 ();
 sg13g2_fill_2 FILLER_11_1533 ();
 sg13g2_fill_1 FILLER_11_1535 ();
 sg13g2_fill_1 FILLER_11_1557 ();
 sg13g2_fill_1 FILLER_11_1580 ();
 sg13g2_fill_2 FILLER_11_1587 ();
 sg13g2_fill_2 FILLER_11_1611 ();
 sg13g2_fill_1 FILLER_11_1613 ();
 sg13g2_decap_8 FILLER_11_1635 ();
 sg13g2_decap_8 FILLER_11_1642 ();
 sg13g2_decap_8 FILLER_11_1649 ();
 sg13g2_fill_2 FILLER_11_1656 ();
 sg13g2_decap_8 FILLER_11_1668 ();
 sg13g2_decap_8 FILLER_11_1675 ();
 sg13g2_fill_2 FILLER_11_1682 ();
 sg13g2_decap_4 FILLER_11_1707 ();
 sg13g2_fill_1 FILLER_11_1711 ();
 sg13g2_fill_1 FILLER_11_1743 ();
 sg13g2_decap_4 FILLER_11_1782 ();
 sg13g2_decap_4 FILLER_11_1820 ();
 sg13g2_fill_1 FILLER_11_1824 ();
 sg13g2_fill_2 FILLER_11_1852 ();
 sg13g2_fill_1 FILLER_11_1854 ();
 sg13g2_fill_2 FILLER_11_1935 ();
 sg13g2_fill_1 FILLER_11_1937 ();
 sg13g2_fill_1 FILLER_11_1966 ();
 sg13g2_fill_2 FILLER_11_1980 ();
 sg13g2_fill_2 FILLER_11_2038 ();
 sg13g2_fill_2 FILLER_11_2074 ();
 sg13g2_fill_1 FILLER_11_2076 ();
 sg13g2_fill_1 FILLER_11_2094 ();
 sg13g2_fill_1 FILLER_11_2133 ();
 sg13g2_fill_2 FILLER_11_2157 ();
 sg13g2_decap_8 FILLER_11_2174 ();
 sg13g2_decap_8 FILLER_11_2181 ();
 sg13g2_decap_8 FILLER_11_2188 ();
 sg13g2_decap_8 FILLER_11_2195 ();
 sg13g2_decap_8 FILLER_11_2202 ();
 sg13g2_decap_8 FILLER_11_2209 ();
 sg13g2_decap_8 FILLER_11_2216 ();
 sg13g2_decap_8 FILLER_11_2223 ();
 sg13g2_decap_8 FILLER_11_2230 ();
 sg13g2_decap_8 FILLER_11_2237 ();
 sg13g2_decap_8 FILLER_11_2244 ();
 sg13g2_decap_8 FILLER_11_2251 ();
 sg13g2_decap_8 FILLER_11_2258 ();
 sg13g2_decap_8 FILLER_11_2265 ();
 sg13g2_decap_8 FILLER_11_2272 ();
 sg13g2_decap_8 FILLER_11_2279 ();
 sg13g2_decap_8 FILLER_11_2286 ();
 sg13g2_decap_8 FILLER_11_2293 ();
 sg13g2_decap_8 FILLER_11_2300 ();
 sg13g2_decap_8 FILLER_11_2307 ();
 sg13g2_decap_8 FILLER_11_2314 ();
 sg13g2_decap_8 FILLER_11_2321 ();
 sg13g2_decap_8 FILLER_11_2328 ();
 sg13g2_decap_8 FILLER_11_2335 ();
 sg13g2_decap_8 FILLER_11_2342 ();
 sg13g2_decap_8 FILLER_11_2349 ();
 sg13g2_decap_8 FILLER_11_2356 ();
 sg13g2_decap_8 FILLER_11_2363 ();
 sg13g2_decap_8 FILLER_11_2370 ();
 sg13g2_decap_8 FILLER_11_2377 ();
 sg13g2_decap_8 FILLER_11_2384 ();
 sg13g2_decap_8 FILLER_11_2391 ();
 sg13g2_decap_8 FILLER_11_2398 ();
 sg13g2_decap_8 FILLER_11_2405 ();
 sg13g2_decap_8 FILLER_11_2412 ();
 sg13g2_decap_8 FILLER_11_2419 ();
 sg13g2_decap_8 FILLER_11_2426 ();
 sg13g2_decap_8 FILLER_11_2433 ();
 sg13g2_decap_8 FILLER_11_2440 ();
 sg13g2_decap_8 FILLER_11_2447 ();
 sg13g2_decap_8 FILLER_11_2454 ();
 sg13g2_decap_8 FILLER_11_2461 ();
 sg13g2_decap_8 FILLER_11_2468 ();
 sg13g2_decap_8 FILLER_11_2475 ();
 sg13g2_decap_8 FILLER_11_2482 ();
 sg13g2_decap_8 FILLER_11_2489 ();
 sg13g2_decap_8 FILLER_11_2496 ();
 sg13g2_decap_8 FILLER_11_2503 ();
 sg13g2_decap_8 FILLER_11_2510 ();
 sg13g2_decap_8 FILLER_11_2517 ();
 sg13g2_decap_8 FILLER_11_2524 ();
 sg13g2_decap_8 FILLER_11_2531 ();
 sg13g2_decap_8 FILLER_11_2538 ();
 sg13g2_decap_8 FILLER_11_2545 ();
 sg13g2_decap_8 FILLER_11_2552 ();
 sg13g2_decap_8 FILLER_11_2559 ();
 sg13g2_decap_8 FILLER_11_2566 ();
 sg13g2_decap_8 FILLER_11_2573 ();
 sg13g2_decap_8 FILLER_11_2580 ();
 sg13g2_decap_8 FILLER_11_2587 ();
 sg13g2_decap_8 FILLER_11_2594 ();
 sg13g2_decap_8 FILLER_11_2601 ();
 sg13g2_decap_8 FILLER_11_2608 ();
 sg13g2_decap_8 FILLER_11_2615 ();
 sg13g2_decap_8 FILLER_11_2622 ();
 sg13g2_decap_8 FILLER_11_2629 ();
 sg13g2_decap_8 FILLER_11_2636 ();
 sg13g2_decap_8 FILLER_11_2643 ();
 sg13g2_decap_8 FILLER_11_2650 ();
 sg13g2_decap_8 FILLER_11_2657 ();
 sg13g2_decap_8 FILLER_11_2664 ();
 sg13g2_fill_2 FILLER_11_2671 ();
 sg13g2_fill_1 FILLER_11_2673 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_118 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_346 ();
 sg13g2_decap_4 FILLER_12_481 ();
 sg13g2_fill_2 FILLER_12_485 ();
 sg13g2_fill_2 FILLER_12_531 ();
 sg13g2_fill_2 FILLER_12_537 ();
 sg13g2_decap_8 FILLER_12_544 ();
 sg13g2_fill_2 FILLER_12_551 ();
 sg13g2_fill_1 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_558 ();
 sg13g2_decap_8 FILLER_12_565 ();
 sg13g2_decap_8 FILLER_12_572 ();
 sg13g2_decap_8 FILLER_12_579 ();
 sg13g2_decap_4 FILLER_12_586 ();
 sg13g2_fill_1 FILLER_12_600 ();
 sg13g2_fill_1 FILLER_12_605 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_643 ();
 sg13g2_decap_8 FILLER_12_650 ();
 sg13g2_fill_2 FILLER_12_657 ();
 sg13g2_fill_1 FILLER_12_664 ();
 sg13g2_fill_2 FILLER_12_677 ();
 sg13g2_decap_8 FILLER_12_685 ();
 sg13g2_decap_4 FILLER_12_692 ();
 sg13g2_fill_1 FILLER_12_696 ();
 sg13g2_decap_4 FILLER_12_707 ();
 sg13g2_fill_2 FILLER_12_711 ();
 sg13g2_fill_2 FILLER_12_748 ();
 sg13g2_fill_2 FILLER_12_789 ();
 sg13g2_fill_1 FILLER_12_791 ();
 sg13g2_fill_2 FILLER_12_820 ();
 sg13g2_fill_1 FILLER_12_835 ();
 sg13g2_fill_1 FILLER_12_848 ();
 sg13g2_fill_2 FILLER_12_867 ();
 sg13g2_fill_2 FILLER_12_884 ();
 sg13g2_fill_1 FILLER_12_944 ();
 sg13g2_decap_4 FILLER_12_972 ();
 sg13g2_fill_2 FILLER_12_976 ();
 sg13g2_decap_8 FILLER_12_987 ();
 sg13g2_fill_2 FILLER_12_994 ();
 sg13g2_decap_4 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1023 ();
 sg13g2_decap_8 FILLER_12_1029 ();
 sg13g2_fill_1 FILLER_12_1036 ();
 sg13g2_fill_1 FILLER_12_1076 ();
 sg13g2_fill_2 FILLER_12_1082 ();
 sg13g2_decap_8 FILLER_12_1100 ();
 sg13g2_decap_4 FILLER_12_1107 ();
 sg13g2_fill_2 FILLER_12_1111 ();
 sg13g2_fill_1 FILLER_12_1131 ();
 sg13g2_fill_1 FILLER_12_1167 ();
 sg13g2_fill_1 FILLER_12_1244 ();
 sg13g2_decap_4 FILLER_12_1263 ();
 sg13g2_decap_4 FILLER_12_1271 ();
 sg13g2_fill_1 FILLER_12_1275 ();
 sg13g2_fill_2 FILLER_12_1304 ();
 sg13g2_fill_1 FILLER_12_1306 ();
 sg13g2_decap_8 FILLER_12_1321 ();
 sg13g2_fill_1 FILLER_12_1328 ();
 sg13g2_decap_4 FILLER_12_1342 ();
 sg13g2_fill_1 FILLER_12_1389 ();
 sg13g2_fill_2 FILLER_12_1400 ();
 sg13g2_fill_1 FILLER_12_1402 ();
 sg13g2_fill_2 FILLER_12_1441 ();
 sg13g2_fill_1 FILLER_12_1443 ();
 sg13g2_fill_1 FILLER_12_1472 ();
 sg13g2_decap_4 FILLER_12_1489 ();
 sg13g2_fill_2 FILLER_12_1511 ();
 sg13g2_fill_1 FILLER_12_1522 ();
 sg13g2_decap_8 FILLER_12_1572 ();
 sg13g2_decap_8 FILLER_12_1579 ();
 sg13g2_fill_2 FILLER_12_1586 ();
 sg13g2_fill_2 FILLER_12_1596 ();
 sg13g2_fill_1 FILLER_12_1598 ();
 sg13g2_fill_2 FILLER_12_1618 ();
 sg13g2_decap_8 FILLER_12_1648 ();
 sg13g2_fill_2 FILLER_12_1655 ();
 sg13g2_fill_2 FILLER_12_1667 ();
 sg13g2_fill_1 FILLER_12_1669 ();
 sg13g2_fill_2 FILLER_12_1763 ();
 sg13g2_fill_1 FILLER_12_1765 ();
 sg13g2_fill_2 FILLER_12_1779 ();
 sg13g2_fill_1 FILLER_12_1781 ();
 sg13g2_fill_2 FILLER_12_1791 ();
 sg13g2_fill_2 FILLER_12_1829 ();
 sg13g2_fill_1 FILLER_12_1831 ();
 sg13g2_decap_4 FILLER_12_1899 ();
 sg13g2_fill_1 FILLER_12_1903 ();
 sg13g2_fill_1 FILLER_12_1924 ();
 sg13g2_decap_4 FILLER_12_1934 ();
 sg13g2_fill_1 FILLER_12_1975 ();
 sg13g2_fill_1 FILLER_12_2059 ();
 sg13g2_fill_2 FILLER_12_2083 ();
 sg13g2_fill_1 FILLER_12_2097 ();
 sg13g2_fill_2 FILLER_12_2138 ();
 sg13g2_fill_1 FILLER_12_2145 ();
 sg13g2_fill_2 FILLER_12_2151 ();
 sg13g2_fill_1 FILLER_12_2153 ();
 sg13g2_decap_8 FILLER_12_2195 ();
 sg13g2_decap_8 FILLER_12_2202 ();
 sg13g2_decap_8 FILLER_12_2209 ();
 sg13g2_decap_8 FILLER_12_2216 ();
 sg13g2_decap_8 FILLER_12_2223 ();
 sg13g2_decap_8 FILLER_12_2230 ();
 sg13g2_decap_8 FILLER_12_2237 ();
 sg13g2_decap_8 FILLER_12_2244 ();
 sg13g2_decap_8 FILLER_12_2251 ();
 sg13g2_decap_8 FILLER_12_2258 ();
 sg13g2_decap_8 FILLER_12_2265 ();
 sg13g2_decap_8 FILLER_12_2272 ();
 sg13g2_decap_8 FILLER_12_2279 ();
 sg13g2_decap_8 FILLER_12_2286 ();
 sg13g2_decap_8 FILLER_12_2293 ();
 sg13g2_decap_8 FILLER_12_2300 ();
 sg13g2_decap_8 FILLER_12_2307 ();
 sg13g2_decap_8 FILLER_12_2314 ();
 sg13g2_decap_8 FILLER_12_2321 ();
 sg13g2_decap_8 FILLER_12_2328 ();
 sg13g2_decap_8 FILLER_12_2335 ();
 sg13g2_decap_8 FILLER_12_2342 ();
 sg13g2_decap_8 FILLER_12_2349 ();
 sg13g2_decap_8 FILLER_12_2356 ();
 sg13g2_decap_8 FILLER_12_2363 ();
 sg13g2_decap_8 FILLER_12_2370 ();
 sg13g2_decap_8 FILLER_12_2377 ();
 sg13g2_decap_8 FILLER_12_2384 ();
 sg13g2_decap_8 FILLER_12_2391 ();
 sg13g2_decap_8 FILLER_12_2398 ();
 sg13g2_decap_8 FILLER_12_2405 ();
 sg13g2_decap_8 FILLER_12_2412 ();
 sg13g2_decap_8 FILLER_12_2419 ();
 sg13g2_decap_8 FILLER_12_2426 ();
 sg13g2_decap_8 FILLER_12_2433 ();
 sg13g2_decap_8 FILLER_12_2440 ();
 sg13g2_decap_8 FILLER_12_2447 ();
 sg13g2_decap_8 FILLER_12_2454 ();
 sg13g2_decap_8 FILLER_12_2461 ();
 sg13g2_decap_8 FILLER_12_2468 ();
 sg13g2_decap_8 FILLER_12_2475 ();
 sg13g2_decap_8 FILLER_12_2482 ();
 sg13g2_decap_8 FILLER_12_2489 ();
 sg13g2_decap_8 FILLER_12_2496 ();
 sg13g2_decap_8 FILLER_12_2503 ();
 sg13g2_decap_8 FILLER_12_2510 ();
 sg13g2_decap_8 FILLER_12_2517 ();
 sg13g2_decap_8 FILLER_12_2524 ();
 sg13g2_decap_8 FILLER_12_2531 ();
 sg13g2_decap_8 FILLER_12_2538 ();
 sg13g2_decap_8 FILLER_12_2545 ();
 sg13g2_decap_8 FILLER_12_2552 ();
 sg13g2_decap_8 FILLER_12_2559 ();
 sg13g2_decap_8 FILLER_12_2566 ();
 sg13g2_decap_8 FILLER_12_2573 ();
 sg13g2_decap_8 FILLER_12_2580 ();
 sg13g2_decap_8 FILLER_12_2587 ();
 sg13g2_decap_8 FILLER_12_2594 ();
 sg13g2_decap_8 FILLER_12_2601 ();
 sg13g2_decap_8 FILLER_12_2608 ();
 sg13g2_decap_8 FILLER_12_2615 ();
 sg13g2_decap_8 FILLER_12_2622 ();
 sg13g2_decap_8 FILLER_12_2629 ();
 sg13g2_decap_8 FILLER_12_2636 ();
 sg13g2_decap_8 FILLER_12_2643 ();
 sg13g2_decap_8 FILLER_12_2650 ();
 sg13g2_decap_8 FILLER_12_2657 ();
 sg13g2_decap_8 FILLER_12_2664 ();
 sg13g2_fill_2 FILLER_12_2671 ();
 sg13g2_fill_1 FILLER_12_2673 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_2 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_53 ();
 sg13g2_fill_2 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_159 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_decap_4 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_457 ();
 sg13g2_decap_8 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_484 ();
 sg13g2_decap_4 FILLER_13_491 ();
 sg13g2_decap_8 FILLER_13_526 ();
 sg13g2_decap_8 FILLER_13_533 ();
 sg13g2_fill_1 FILLER_13_587 ();
 sg13g2_fill_2 FILLER_13_601 ();
 sg13g2_fill_1 FILLER_13_603 ();
 sg13g2_decap_4 FILLER_13_619 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_fill_2 FILLER_13_649 ();
 sg13g2_fill_2 FILLER_13_661 ();
 sg13g2_fill_1 FILLER_13_663 ();
 sg13g2_decap_4 FILLER_13_672 ();
 sg13g2_fill_2 FILLER_13_681 ();
 sg13g2_fill_2 FILLER_13_704 ();
 sg13g2_decap_4 FILLER_13_740 ();
 sg13g2_fill_2 FILLER_13_755 ();
 sg13g2_fill_1 FILLER_13_764 ();
 sg13g2_fill_2 FILLER_13_779 ();
 sg13g2_fill_2 FILLER_13_789 ();
 sg13g2_fill_1 FILLER_13_791 ();
 sg13g2_fill_1 FILLER_13_801 ();
 sg13g2_decap_4 FILLER_13_811 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_fill_1 FILLER_13_863 ();
 sg13g2_fill_2 FILLER_13_898 ();
 sg13g2_fill_2 FILLER_13_941 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_4 FILLER_13_998 ();
 sg13g2_fill_1 FILLER_13_1002 ();
 sg13g2_decap_4 FILLER_13_1008 ();
 sg13g2_fill_1 FILLER_13_1012 ();
 sg13g2_decap_4 FILLER_13_1018 ();
 sg13g2_decap_8 FILLER_13_1035 ();
 sg13g2_fill_2 FILLER_13_1042 ();
 sg13g2_fill_1 FILLER_13_1051 ();
 sg13g2_fill_2 FILLER_13_1064 ();
 sg13g2_fill_1 FILLER_13_1066 ();
 sg13g2_decap_8 FILLER_13_1106 ();
 sg13g2_fill_2 FILLER_13_1113 ();
 sg13g2_fill_1 FILLER_13_1115 ();
 sg13g2_fill_2 FILLER_13_1167 ();
 sg13g2_fill_1 FILLER_13_1169 ();
 sg13g2_fill_1 FILLER_13_1184 ();
 sg13g2_fill_1 FILLER_13_1268 ();
 sg13g2_fill_1 FILLER_13_1307 ();
 sg13g2_decap_8 FILLER_13_1321 ();
 sg13g2_decap_4 FILLER_13_1328 ();
 sg13g2_fill_1 FILLER_13_1332 ();
 sg13g2_decap_8 FILLER_13_1342 ();
 sg13g2_fill_2 FILLER_13_1349 ();
 sg13g2_decap_4 FILLER_13_1356 ();
 sg13g2_fill_1 FILLER_13_1364 ();
 sg13g2_fill_2 FILLER_13_1379 ();
 sg13g2_fill_2 FILLER_13_1386 ();
 sg13g2_fill_1 FILLER_13_1388 ();
 sg13g2_decap_8 FILLER_13_1411 ();
 sg13g2_fill_2 FILLER_13_1418 ();
 sg13g2_fill_1 FILLER_13_1420 ();
 sg13g2_fill_2 FILLER_13_1478 ();
 sg13g2_fill_1 FILLER_13_1480 ();
 sg13g2_fill_1 FILLER_13_1527 ();
 sg13g2_fill_2 FILLER_13_1560 ();
 sg13g2_decap_8 FILLER_13_1590 ();
 sg13g2_decap_8 FILLER_13_1597 ();
 sg13g2_fill_2 FILLER_13_1604 ();
 sg13g2_decap_4 FILLER_13_1624 ();
 sg13g2_fill_2 FILLER_13_1628 ();
 sg13g2_decap_4 FILLER_13_1658 ();
 sg13g2_fill_2 FILLER_13_1662 ();
 sg13g2_fill_1 FILLER_13_1704 ();
 sg13g2_fill_1 FILLER_13_1751 ();
 sg13g2_fill_2 FILLER_13_1765 ();
 sg13g2_fill_1 FILLER_13_1767 ();
 sg13g2_fill_2 FILLER_13_1873 ();
 sg13g2_fill_1 FILLER_13_1875 ();
 sg13g2_fill_2 FILLER_13_1917 ();
 sg13g2_fill_1 FILLER_13_1919 ();
 sg13g2_decap_8 FILLER_13_1925 ();
 sg13g2_decap_8 FILLER_13_1932 ();
 sg13g2_fill_1 FILLER_13_1939 ();
 sg13g2_fill_1 FILLER_13_1963 ();
 sg13g2_fill_1 FILLER_13_2056 ();
 sg13g2_fill_1 FILLER_13_2091 ();
 sg13g2_fill_1 FILLER_13_2109 ();
 sg13g2_fill_1 FILLER_13_2125 ();
 sg13g2_fill_1 FILLER_13_2135 ();
 sg13g2_decap_8 FILLER_13_2204 ();
 sg13g2_decap_8 FILLER_13_2211 ();
 sg13g2_decap_8 FILLER_13_2218 ();
 sg13g2_decap_8 FILLER_13_2225 ();
 sg13g2_decap_8 FILLER_13_2232 ();
 sg13g2_decap_8 FILLER_13_2239 ();
 sg13g2_decap_8 FILLER_13_2246 ();
 sg13g2_decap_8 FILLER_13_2253 ();
 sg13g2_decap_8 FILLER_13_2260 ();
 sg13g2_decap_8 FILLER_13_2267 ();
 sg13g2_decap_8 FILLER_13_2274 ();
 sg13g2_decap_8 FILLER_13_2281 ();
 sg13g2_decap_8 FILLER_13_2288 ();
 sg13g2_decap_8 FILLER_13_2295 ();
 sg13g2_decap_8 FILLER_13_2302 ();
 sg13g2_decap_8 FILLER_13_2309 ();
 sg13g2_decap_8 FILLER_13_2316 ();
 sg13g2_decap_8 FILLER_13_2323 ();
 sg13g2_decap_8 FILLER_13_2330 ();
 sg13g2_decap_8 FILLER_13_2337 ();
 sg13g2_decap_8 FILLER_13_2344 ();
 sg13g2_decap_8 FILLER_13_2351 ();
 sg13g2_decap_8 FILLER_13_2358 ();
 sg13g2_decap_8 FILLER_13_2365 ();
 sg13g2_decap_8 FILLER_13_2372 ();
 sg13g2_decap_8 FILLER_13_2379 ();
 sg13g2_decap_8 FILLER_13_2386 ();
 sg13g2_decap_8 FILLER_13_2393 ();
 sg13g2_decap_8 FILLER_13_2400 ();
 sg13g2_decap_8 FILLER_13_2407 ();
 sg13g2_decap_8 FILLER_13_2414 ();
 sg13g2_decap_8 FILLER_13_2421 ();
 sg13g2_decap_8 FILLER_13_2428 ();
 sg13g2_decap_8 FILLER_13_2435 ();
 sg13g2_decap_8 FILLER_13_2442 ();
 sg13g2_decap_8 FILLER_13_2449 ();
 sg13g2_decap_8 FILLER_13_2456 ();
 sg13g2_decap_8 FILLER_13_2463 ();
 sg13g2_decap_8 FILLER_13_2470 ();
 sg13g2_decap_8 FILLER_13_2477 ();
 sg13g2_decap_8 FILLER_13_2484 ();
 sg13g2_decap_8 FILLER_13_2491 ();
 sg13g2_decap_8 FILLER_13_2498 ();
 sg13g2_decap_8 FILLER_13_2505 ();
 sg13g2_decap_8 FILLER_13_2512 ();
 sg13g2_decap_8 FILLER_13_2519 ();
 sg13g2_decap_8 FILLER_13_2526 ();
 sg13g2_decap_8 FILLER_13_2533 ();
 sg13g2_decap_8 FILLER_13_2540 ();
 sg13g2_decap_8 FILLER_13_2547 ();
 sg13g2_decap_8 FILLER_13_2554 ();
 sg13g2_decap_8 FILLER_13_2561 ();
 sg13g2_decap_8 FILLER_13_2568 ();
 sg13g2_decap_8 FILLER_13_2575 ();
 sg13g2_decap_8 FILLER_13_2582 ();
 sg13g2_decap_8 FILLER_13_2589 ();
 sg13g2_decap_8 FILLER_13_2596 ();
 sg13g2_decap_8 FILLER_13_2603 ();
 sg13g2_decap_8 FILLER_13_2610 ();
 sg13g2_decap_8 FILLER_13_2617 ();
 sg13g2_decap_8 FILLER_13_2624 ();
 sg13g2_decap_8 FILLER_13_2631 ();
 sg13g2_decap_8 FILLER_13_2638 ();
 sg13g2_decap_8 FILLER_13_2645 ();
 sg13g2_decap_8 FILLER_13_2652 ();
 sg13g2_decap_8 FILLER_13_2659 ();
 sg13g2_decap_8 FILLER_13_2666 ();
 sg13g2_fill_1 FILLER_13_2673 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_32 ();
 sg13g2_fill_1 FILLER_14_34 ();
 sg13g2_fill_2 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_169 ();
 sg13g2_decap_4 FILLER_14_215 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_306 ();
 sg13g2_decap_4 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_fill_2 FILLER_14_430 ();
 sg13g2_fill_1 FILLER_14_432 ();
 sg13g2_decap_8 FILLER_14_446 ();
 sg13g2_decap_8 FILLER_14_453 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_4 FILLER_14_483 ();
 sg13g2_fill_2 FILLER_14_487 ();
 sg13g2_decap_4 FILLER_14_496 ();
 sg13g2_fill_1 FILLER_14_500 ();
 sg13g2_fill_2 FILLER_14_519 ();
 sg13g2_fill_1 FILLER_14_521 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_586 ();
 sg13g2_decap_8 FILLER_14_597 ();
 sg13g2_fill_1 FILLER_14_604 ();
 sg13g2_fill_2 FILLER_14_633 ();
 sg13g2_fill_1 FILLER_14_635 ();
 sg13g2_decap_4 FILLER_14_644 ();
 sg13g2_fill_2 FILLER_14_653 ();
 sg13g2_fill_1 FILLER_14_680 ();
 sg13g2_decap_8 FILLER_14_687 ();
 sg13g2_decap_8 FILLER_14_694 ();
 sg13g2_decap_8 FILLER_14_701 ();
 sg13g2_decap_4 FILLER_14_708 ();
 sg13g2_fill_2 FILLER_14_712 ();
 sg13g2_decap_4 FILLER_14_740 ();
 sg13g2_fill_1 FILLER_14_773 ();
 sg13g2_fill_1 FILLER_14_779 ();
 sg13g2_fill_2 FILLER_14_785 ();
 sg13g2_fill_1 FILLER_14_787 ();
 sg13g2_fill_2 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_4 FILLER_14_852 ();
 sg13g2_fill_1 FILLER_14_892 ();
 sg13g2_fill_2 FILLER_14_933 ();
 sg13g2_fill_1 FILLER_14_962 ();
 sg13g2_fill_2 FILLER_14_976 ();
 sg13g2_decap_8 FILLER_14_987 ();
 sg13g2_decap_8 FILLER_14_994 ();
 sg13g2_decap_8 FILLER_14_1001 ();
 sg13g2_fill_1 FILLER_14_1008 ();
 sg13g2_fill_1 FILLER_14_1054 ();
 sg13g2_fill_1 FILLER_14_1065 ();
 sg13g2_decap_8 FILLER_14_1071 ();
 sg13g2_decap_4 FILLER_14_1078 ();
 sg13g2_fill_2 FILLER_14_1082 ();
 sg13g2_fill_2 FILLER_14_1091 ();
 sg13g2_fill_1 FILLER_14_1093 ();
 sg13g2_decap_4 FILLER_14_1119 ();
 sg13g2_fill_2 FILLER_14_1123 ();
 sg13g2_fill_2 FILLER_14_1171 ();
 sg13g2_decap_8 FILLER_14_1214 ();
 sg13g2_decap_4 FILLER_14_1221 ();
 sg13g2_fill_2 FILLER_14_1286 ();
 sg13g2_fill_1 FILLER_14_1315 ();
 sg13g2_fill_1 FILLER_14_1320 ();
 sg13g2_decap_4 FILLER_14_1331 ();
 sg13g2_fill_1 FILLER_14_1335 ();
 sg13g2_fill_1 FILLER_14_1381 ();
 sg13g2_decap_8 FILLER_14_1387 ();
 sg13g2_fill_2 FILLER_14_1394 ();
 sg13g2_decap_8 FILLER_14_1417 ();
 sg13g2_fill_1 FILLER_14_1424 ();
 sg13g2_decap_4 FILLER_14_1431 ();
 sg13g2_decap_4 FILLER_14_1472 ();
 sg13g2_fill_2 FILLER_14_1476 ();
 sg13g2_fill_2 FILLER_14_1505 ();
 sg13g2_fill_1 FILLER_14_1507 ();
 sg13g2_fill_2 FILLER_14_1549 ();
 sg13g2_decap_8 FILLER_14_1584 ();
 sg13g2_decap_4 FILLER_14_1591 ();
 sg13g2_fill_1 FILLER_14_1595 ();
 sg13g2_decap_4 FILLER_14_1600 ();
 sg13g2_decap_4 FILLER_14_1625 ();
 sg13g2_fill_2 FILLER_14_1629 ();
 sg13g2_decap_4 FILLER_14_1641 ();
 sg13g2_fill_2 FILLER_14_1645 ();
 sg13g2_decap_8 FILLER_14_1687 ();
 sg13g2_fill_1 FILLER_14_1694 ();
 sg13g2_fill_1 FILLER_14_1721 ();
 sg13g2_fill_2 FILLER_14_1742 ();
 sg13g2_fill_1 FILLER_14_1744 ();
 sg13g2_fill_2 FILLER_14_1787 ();
 sg13g2_fill_1 FILLER_14_1789 ();
 sg13g2_fill_2 FILLER_14_1823 ();
 sg13g2_fill_2 FILLER_14_1834 ();
 sg13g2_fill_2 FILLER_14_1873 ();
 sg13g2_fill_1 FILLER_14_1884 ();
 sg13g2_decap_4 FILLER_14_1913 ();
 sg13g2_decap_4 FILLER_14_1945 ();
 sg13g2_fill_1 FILLER_14_1959 ();
 sg13g2_fill_1 FILLER_14_2016 ();
 sg13g2_fill_2 FILLER_14_2038 ();
 sg13g2_fill_2 FILLER_14_2084 ();
 sg13g2_fill_1 FILLER_14_2086 ();
 sg13g2_fill_1 FILLER_14_2105 ();
 sg13g2_fill_2 FILLER_14_2169 ();
 sg13g2_fill_1 FILLER_14_2171 ();
 sg13g2_decap_8 FILLER_14_2221 ();
 sg13g2_decap_8 FILLER_14_2228 ();
 sg13g2_decap_8 FILLER_14_2235 ();
 sg13g2_decap_8 FILLER_14_2242 ();
 sg13g2_decap_8 FILLER_14_2249 ();
 sg13g2_decap_8 FILLER_14_2256 ();
 sg13g2_decap_8 FILLER_14_2263 ();
 sg13g2_decap_8 FILLER_14_2270 ();
 sg13g2_decap_8 FILLER_14_2277 ();
 sg13g2_decap_8 FILLER_14_2284 ();
 sg13g2_decap_8 FILLER_14_2291 ();
 sg13g2_decap_8 FILLER_14_2298 ();
 sg13g2_decap_8 FILLER_14_2305 ();
 sg13g2_decap_8 FILLER_14_2312 ();
 sg13g2_decap_8 FILLER_14_2319 ();
 sg13g2_decap_8 FILLER_14_2326 ();
 sg13g2_decap_8 FILLER_14_2333 ();
 sg13g2_decap_8 FILLER_14_2340 ();
 sg13g2_decap_8 FILLER_14_2347 ();
 sg13g2_decap_8 FILLER_14_2354 ();
 sg13g2_decap_8 FILLER_14_2361 ();
 sg13g2_decap_8 FILLER_14_2368 ();
 sg13g2_decap_8 FILLER_14_2375 ();
 sg13g2_decap_8 FILLER_14_2382 ();
 sg13g2_decap_8 FILLER_14_2389 ();
 sg13g2_decap_8 FILLER_14_2396 ();
 sg13g2_decap_8 FILLER_14_2403 ();
 sg13g2_decap_8 FILLER_14_2410 ();
 sg13g2_decap_8 FILLER_14_2417 ();
 sg13g2_decap_8 FILLER_14_2424 ();
 sg13g2_decap_8 FILLER_14_2431 ();
 sg13g2_decap_8 FILLER_14_2438 ();
 sg13g2_decap_8 FILLER_14_2445 ();
 sg13g2_decap_8 FILLER_14_2452 ();
 sg13g2_decap_8 FILLER_14_2459 ();
 sg13g2_decap_8 FILLER_14_2466 ();
 sg13g2_decap_8 FILLER_14_2473 ();
 sg13g2_decap_8 FILLER_14_2480 ();
 sg13g2_decap_8 FILLER_14_2487 ();
 sg13g2_decap_8 FILLER_14_2494 ();
 sg13g2_decap_8 FILLER_14_2501 ();
 sg13g2_decap_8 FILLER_14_2508 ();
 sg13g2_decap_8 FILLER_14_2515 ();
 sg13g2_decap_8 FILLER_14_2522 ();
 sg13g2_decap_8 FILLER_14_2529 ();
 sg13g2_decap_8 FILLER_14_2536 ();
 sg13g2_decap_8 FILLER_14_2543 ();
 sg13g2_decap_8 FILLER_14_2550 ();
 sg13g2_decap_8 FILLER_14_2557 ();
 sg13g2_decap_8 FILLER_14_2564 ();
 sg13g2_decap_8 FILLER_14_2571 ();
 sg13g2_decap_8 FILLER_14_2578 ();
 sg13g2_decap_8 FILLER_14_2585 ();
 sg13g2_decap_8 FILLER_14_2592 ();
 sg13g2_decap_8 FILLER_14_2599 ();
 sg13g2_decap_8 FILLER_14_2606 ();
 sg13g2_decap_8 FILLER_14_2613 ();
 sg13g2_decap_8 FILLER_14_2620 ();
 sg13g2_decap_8 FILLER_14_2627 ();
 sg13g2_decap_8 FILLER_14_2634 ();
 sg13g2_decap_8 FILLER_14_2641 ();
 sg13g2_decap_8 FILLER_14_2648 ();
 sg13g2_decap_8 FILLER_14_2655 ();
 sg13g2_decap_8 FILLER_14_2662 ();
 sg13g2_decap_4 FILLER_14_2669 ();
 sg13g2_fill_1 FILLER_14_2673 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_390 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_fill_1 FILLER_15_414 ();
 sg13g2_decap_4 FILLER_15_478 ();
 sg13g2_fill_1 FILLER_15_482 ();
 sg13g2_fill_2 FILLER_15_495 ();
 sg13g2_fill_1 FILLER_15_497 ();
 sg13g2_fill_2 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_fill_2 FILLER_15_550 ();
 sg13g2_decap_4 FILLER_15_565 ();
 sg13g2_fill_1 FILLER_15_569 ();
 sg13g2_decap_4 FILLER_15_580 ();
 sg13g2_fill_2 FILLER_15_584 ();
 sg13g2_decap_4 FILLER_15_603 ();
 sg13g2_decap_4 FILLER_15_615 ();
 sg13g2_fill_2 FILLER_15_624 ();
 sg13g2_decap_4 FILLER_15_631 ();
 sg13g2_fill_2 FILLER_15_640 ();
 sg13g2_fill_1 FILLER_15_642 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_fill_2 FILLER_15_661 ();
 sg13g2_fill_1 FILLER_15_663 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_4 FILLER_15_717 ();
 sg13g2_fill_1 FILLER_15_721 ();
 sg13g2_fill_1 FILLER_15_727 ();
 sg13g2_decap_8 FILLER_15_734 ();
 sg13g2_fill_2 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_783 ();
 sg13g2_decap_8 FILLER_15_790 ();
 sg13g2_fill_2 FILLER_15_797 ();
 sg13g2_fill_1 FILLER_15_799 ();
 sg13g2_fill_2 FILLER_15_900 ();
 sg13g2_fill_2 FILLER_15_937 ();
 sg13g2_fill_1 FILLER_15_971 ();
 sg13g2_fill_2 FILLER_15_1056 ();
 sg13g2_decap_8 FILLER_15_1064 ();
 sg13g2_decap_8 FILLER_15_1071 ();
 sg13g2_fill_2 FILLER_15_1078 ();
 sg13g2_fill_1 FILLER_15_1080 ();
 sg13g2_fill_2 FILLER_15_1138 ();
 sg13g2_fill_1 FILLER_15_1140 ();
 sg13g2_decap_4 FILLER_15_1214 ();
 sg13g2_fill_2 FILLER_15_1224 ();
 sg13g2_fill_2 FILLER_15_1412 ();
 sg13g2_fill_1 FILLER_15_1414 ();
 sg13g2_fill_2 FILLER_15_1420 ();
 sg13g2_fill_2 FILLER_15_1427 ();
 sg13g2_decap_4 FILLER_15_1466 ();
 sg13g2_fill_2 FILLER_15_1470 ();
 sg13g2_fill_1 FILLER_15_1519 ();
 sg13g2_fill_1 FILLER_15_1536 ();
 sg13g2_decap_8 FILLER_15_1550 ();
 sg13g2_fill_1 FILLER_15_1557 ();
 sg13g2_decap_8 FILLER_15_1568 ();
 sg13g2_fill_1 FILLER_15_1575 ();
 sg13g2_fill_2 FILLER_15_1598 ();
 sg13g2_decap_8 FILLER_15_1627 ();
 sg13g2_decap_8 FILLER_15_1634 ();
 sg13g2_decap_4 FILLER_15_1641 ();
 sg13g2_decap_8 FILLER_15_1683 ();
 sg13g2_fill_1 FILLER_15_1721 ();
 sg13g2_fill_2 FILLER_15_1736 ();
 sg13g2_fill_1 FILLER_15_1738 ();
 sg13g2_fill_2 FILLER_15_1744 ();
 sg13g2_fill_2 FILLER_15_1756 ();
 sg13g2_fill_2 FILLER_15_1764 ();
 sg13g2_fill_1 FILLER_15_1792 ();
 sg13g2_fill_2 FILLER_15_1802 ();
 sg13g2_fill_2 FILLER_15_1827 ();
 sg13g2_fill_1 FILLER_15_1829 ();
 sg13g2_fill_1 FILLER_15_1915 ();
 sg13g2_fill_1 FILLER_15_1983 ();
 sg13g2_fill_1 FILLER_15_1998 ();
 sg13g2_fill_1 FILLER_15_2047 ();
 sg13g2_fill_1 FILLER_15_2065 ();
 sg13g2_fill_2 FILLER_15_2071 ();
 sg13g2_fill_2 FILLER_15_2092 ();
 sg13g2_decap_4 FILLER_15_2155 ();
 sg13g2_fill_1 FILLER_15_2159 ();
 sg13g2_decap_8 FILLER_15_2204 ();
 sg13g2_fill_2 FILLER_15_2211 ();
 sg13g2_decap_4 FILLER_15_2218 ();
 sg13g2_decap_8 FILLER_15_2231 ();
 sg13g2_decap_8 FILLER_15_2238 ();
 sg13g2_decap_8 FILLER_15_2245 ();
 sg13g2_decap_8 FILLER_15_2252 ();
 sg13g2_decap_8 FILLER_15_2259 ();
 sg13g2_decap_8 FILLER_15_2266 ();
 sg13g2_decap_8 FILLER_15_2273 ();
 sg13g2_decap_8 FILLER_15_2280 ();
 sg13g2_decap_8 FILLER_15_2287 ();
 sg13g2_decap_8 FILLER_15_2294 ();
 sg13g2_decap_8 FILLER_15_2301 ();
 sg13g2_decap_8 FILLER_15_2308 ();
 sg13g2_decap_8 FILLER_15_2315 ();
 sg13g2_decap_8 FILLER_15_2322 ();
 sg13g2_decap_8 FILLER_15_2329 ();
 sg13g2_decap_8 FILLER_15_2336 ();
 sg13g2_decap_8 FILLER_15_2343 ();
 sg13g2_decap_8 FILLER_15_2350 ();
 sg13g2_decap_8 FILLER_15_2357 ();
 sg13g2_decap_8 FILLER_15_2364 ();
 sg13g2_decap_8 FILLER_15_2371 ();
 sg13g2_decap_8 FILLER_15_2378 ();
 sg13g2_decap_8 FILLER_15_2385 ();
 sg13g2_decap_8 FILLER_15_2392 ();
 sg13g2_decap_8 FILLER_15_2399 ();
 sg13g2_decap_8 FILLER_15_2406 ();
 sg13g2_decap_8 FILLER_15_2413 ();
 sg13g2_decap_8 FILLER_15_2420 ();
 sg13g2_decap_8 FILLER_15_2427 ();
 sg13g2_decap_8 FILLER_15_2434 ();
 sg13g2_decap_8 FILLER_15_2441 ();
 sg13g2_decap_8 FILLER_15_2448 ();
 sg13g2_decap_8 FILLER_15_2455 ();
 sg13g2_decap_8 FILLER_15_2462 ();
 sg13g2_decap_8 FILLER_15_2469 ();
 sg13g2_decap_8 FILLER_15_2476 ();
 sg13g2_decap_8 FILLER_15_2483 ();
 sg13g2_decap_8 FILLER_15_2490 ();
 sg13g2_decap_8 FILLER_15_2497 ();
 sg13g2_decap_8 FILLER_15_2504 ();
 sg13g2_decap_8 FILLER_15_2511 ();
 sg13g2_decap_8 FILLER_15_2518 ();
 sg13g2_decap_8 FILLER_15_2525 ();
 sg13g2_decap_8 FILLER_15_2532 ();
 sg13g2_decap_8 FILLER_15_2539 ();
 sg13g2_decap_8 FILLER_15_2546 ();
 sg13g2_decap_8 FILLER_15_2553 ();
 sg13g2_decap_8 FILLER_15_2560 ();
 sg13g2_decap_8 FILLER_15_2567 ();
 sg13g2_decap_8 FILLER_15_2574 ();
 sg13g2_decap_8 FILLER_15_2581 ();
 sg13g2_decap_8 FILLER_15_2588 ();
 sg13g2_decap_8 FILLER_15_2595 ();
 sg13g2_decap_8 FILLER_15_2602 ();
 sg13g2_decap_8 FILLER_15_2609 ();
 sg13g2_decap_8 FILLER_15_2616 ();
 sg13g2_decap_8 FILLER_15_2623 ();
 sg13g2_decap_8 FILLER_15_2630 ();
 sg13g2_decap_8 FILLER_15_2637 ();
 sg13g2_decap_8 FILLER_15_2644 ();
 sg13g2_decap_8 FILLER_15_2651 ();
 sg13g2_decap_8 FILLER_15_2658 ();
 sg13g2_decap_8 FILLER_15_2665 ();
 sg13g2_fill_2 FILLER_15_2672 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_decap_4 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_decap_4 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_401 ();
 sg13g2_fill_2 FILLER_16_439 ();
 sg13g2_fill_1 FILLER_16_441 ();
 sg13g2_decap_4 FILLER_16_473 ();
 sg13g2_fill_2 FILLER_16_477 ();
 sg13g2_fill_2 FILLER_16_505 ();
 sg13g2_decap_8 FILLER_16_538 ();
 sg13g2_fill_2 FILLER_16_563 ();
 sg13g2_fill_1 FILLER_16_565 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_fill_1 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_605 ();
 sg13g2_decap_4 FILLER_16_612 ();
 sg13g2_fill_1 FILLER_16_616 ();
 sg13g2_fill_1 FILLER_16_621 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_fill_1 FILLER_16_640 ();
 sg13g2_decap_8 FILLER_16_649 ();
 sg13g2_fill_1 FILLER_16_669 ();
 sg13g2_fill_2 FILLER_16_681 ();
 sg13g2_fill_1 FILLER_16_683 ();
 sg13g2_fill_1 FILLER_16_694 ();
 sg13g2_decap_4 FILLER_16_704 ();
 sg13g2_fill_1 FILLER_16_713 ();
 sg13g2_decap_8 FILLER_16_719 ();
 sg13g2_decap_8 FILLER_16_726 ();
 sg13g2_decap_4 FILLER_16_733 ();
 sg13g2_fill_1 FILLER_16_737 ();
 sg13g2_decap_4 FILLER_16_744 ();
 sg13g2_fill_1 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_4 FILLER_16_812 ();
 sg13g2_decap_4 FILLER_16_819 ();
 sg13g2_fill_2 FILLER_16_823 ();
 sg13g2_decap_4 FILLER_16_834 ();
 sg13g2_fill_2 FILLER_16_865 ();
 sg13g2_fill_2 FILLER_16_890 ();
 sg13g2_fill_1 FILLER_16_905 ();
 sg13g2_fill_2 FILLER_16_967 ();
 sg13g2_fill_1 FILLER_16_969 ();
 sg13g2_fill_2 FILLER_16_978 ();
 sg13g2_fill_2 FILLER_16_1032 ();
 sg13g2_decap_8 FILLER_16_1056 ();
 sg13g2_decap_8 FILLER_16_1063 ();
 sg13g2_decap_8 FILLER_16_1070 ();
 sg13g2_decap_8 FILLER_16_1077 ();
 sg13g2_fill_1 FILLER_16_1084 ();
 sg13g2_fill_1 FILLER_16_1133 ();
 sg13g2_fill_1 FILLER_16_1240 ();
 sg13g2_fill_1 FILLER_16_1264 ();
 sg13g2_fill_1 FILLER_16_1380 ();
 sg13g2_fill_1 FILLER_16_1386 ();
 sg13g2_fill_1 FILLER_16_1415 ();
 sg13g2_decap_4 FILLER_16_1437 ();
 sg13g2_fill_1 FILLER_16_1460 ();
 sg13g2_fill_2 FILLER_16_1490 ();
 sg13g2_fill_2 FILLER_16_1559 ();
 sg13g2_fill_1 FILLER_16_1561 ();
 sg13g2_decap_8 FILLER_16_1566 ();
 sg13g2_decap_4 FILLER_16_1578 ();
 sg13g2_fill_1 FILLER_16_1582 ();
 sg13g2_decap_8 FILLER_16_1587 ();
 sg13g2_fill_1 FILLER_16_1594 ();
 sg13g2_fill_1 FILLER_16_1633 ();
 sg13g2_fill_2 FILLER_16_1698 ();
 sg13g2_fill_2 FILLER_16_1740 ();
 sg13g2_fill_1 FILLER_16_1742 ();
 sg13g2_fill_2 FILLER_16_1775 ();
 sg13g2_fill_2 FILLER_16_1832 ();
 sg13g2_fill_2 FILLER_16_1862 ();
 sg13g2_fill_1 FILLER_16_1869 ();
 sg13g2_fill_2 FILLER_16_1945 ();
 sg13g2_fill_2 FILLER_16_2023 ();
 sg13g2_fill_2 FILLER_16_2045 ();
 sg13g2_fill_1 FILLER_16_2047 ();
 sg13g2_fill_2 FILLER_16_2060 ();
 sg13g2_fill_1 FILLER_16_2062 ();
 sg13g2_fill_1 FILLER_16_2149 ();
 sg13g2_fill_2 FILLER_16_2200 ();
 sg13g2_decap_8 FILLER_16_2238 ();
 sg13g2_decap_8 FILLER_16_2245 ();
 sg13g2_decap_8 FILLER_16_2252 ();
 sg13g2_decap_8 FILLER_16_2259 ();
 sg13g2_decap_8 FILLER_16_2266 ();
 sg13g2_decap_8 FILLER_16_2273 ();
 sg13g2_decap_8 FILLER_16_2280 ();
 sg13g2_decap_8 FILLER_16_2287 ();
 sg13g2_decap_8 FILLER_16_2294 ();
 sg13g2_decap_8 FILLER_16_2301 ();
 sg13g2_decap_8 FILLER_16_2308 ();
 sg13g2_decap_8 FILLER_16_2315 ();
 sg13g2_decap_8 FILLER_16_2322 ();
 sg13g2_decap_8 FILLER_16_2329 ();
 sg13g2_decap_8 FILLER_16_2336 ();
 sg13g2_decap_8 FILLER_16_2343 ();
 sg13g2_decap_8 FILLER_16_2350 ();
 sg13g2_decap_8 FILLER_16_2357 ();
 sg13g2_decap_8 FILLER_16_2364 ();
 sg13g2_decap_8 FILLER_16_2371 ();
 sg13g2_decap_8 FILLER_16_2378 ();
 sg13g2_decap_8 FILLER_16_2385 ();
 sg13g2_decap_8 FILLER_16_2392 ();
 sg13g2_decap_8 FILLER_16_2399 ();
 sg13g2_decap_8 FILLER_16_2406 ();
 sg13g2_decap_8 FILLER_16_2413 ();
 sg13g2_decap_8 FILLER_16_2420 ();
 sg13g2_decap_8 FILLER_16_2427 ();
 sg13g2_decap_8 FILLER_16_2434 ();
 sg13g2_decap_8 FILLER_16_2441 ();
 sg13g2_decap_8 FILLER_16_2448 ();
 sg13g2_decap_8 FILLER_16_2455 ();
 sg13g2_decap_8 FILLER_16_2462 ();
 sg13g2_decap_8 FILLER_16_2469 ();
 sg13g2_decap_8 FILLER_16_2476 ();
 sg13g2_decap_8 FILLER_16_2483 ();
 sg13g2_decap_8 FILLER_16_2490 ();
 sg13g2_decap_8 FILLER_16_2497 ();
 sg13g2_decap_8 FILLER_16_2504 ();
 sg13g2_decap_8 FILLER_16_2511 ();
 sg13g2_decap_8 FILLER_16_2518 ();
 sg13g2_decap_8 FILLER_16_2525 ();
 sg13g2_decap_8 FILLER_16_2532 ();
 sg13g2_decap_8 FILLER_16_2539 ();
 sg13g2_decap_8 FILLER_16_2546 ();
 sg13g2_decap_8 FILLER_16_2553 ();
 sg13g2_decap_8 FILLER_16_2560 ();
 sg13g2_decap_8 FILLER_16_2567 ();
 sg13g2_decap_8 FILLER_16_2574 ();
 sg13g2_decap_8 FILLER_16_2581 ();
 sg13g2_decap_8 FILLER_16_2588 ();
 sg13g2_decap_8 FILLER_16_2595 ();
 sg13g2_decap_8 FILLER_16_2602 ();
 sg13g2_decap_8 FILLER_16_2609 ();
 sg13g2_decap_8 FILLER_16_2616 ();
 sg13g2_decap_8 FILLER_16_2623 ();
 sg13g2_decap_8 FILLER_16_2630 ();
 sg13g2_decap_8 FILLER_16_2637 ();
 sg13g2_decap_8 FILLER_16_2644 ();
 sg13g2_decap_8 FILLER_16_2651 ();
 sg13g2_decap_8 FILLER_16_2658 ();
 sg13g2_decap_8 FILLER_16_2665 ();
 sg13g2_fill_2 FILLER_16_2672 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_31 ();
 sg13g2_decap_8 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_155 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_decap_4 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_decap_4 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_decap_4 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_361 ();
 sg13g2_fill_1 FILLER_17_404 ();
 sg13g2_fill_2 FILLER_17_461 ();
 sg13g2_fill_1 FILLER_17_463 ();
 sg13g2_fill_1 FILLER_17_473 ();
 sg13g2_decap_4 FILLER_17_527 ();
 sg13g2_fill_1 FILLER_17_531 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_fill_2 FILLER_17_560 ();
 sg13g2_fill_1 FILLER_17_562 ();
 sg13g2_fill_1 FILLER_17_568 ();
 sg13g2_decap_8 FILLER_17_573 ();
 sg13g2_decap_4 FILLER_17_580 ();
 sg13g2_decap_4 FILLER_17_588 ();
 sg13g2_fill_2 FILLER_17_592 ();
 sg13g2_decap_4 FILLER_17_599 ();
 sg13g2_fill_2 FILLER_17_603 ();
 sg13g2_decap_8 FILLER_17_610 ();
 sg13g2_decap_8 FILLER_17_617 ();
 sg13g2_fill_2 FILLER_17_624 ();
 sg13g2_fill_1 FILLER_17_626 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_fill_1 FILLER_17_648 ();
 sg13g2_fill_2 FILLER_17_675 ();
 sg13g2_fill_1 FILLER_17_688 ();
 sg13g2_decap_8 FILLER_17_699 ();
 sg13g2_fill_2 FILLER_17_706 ();
 sg13g2_fill_1 FILLER_17_708 ();
 sg13g2_decap_8 FILLER_17_724 ();
 sg13g2_decap_4 FILLER_17_731 ();
 sg13g2_fill_2 FILLER_17_735 ();
 sg13g2_decap_4 FILLER_17_748 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_4 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_fill_1 FILLER_17_830 ();
 sg13g2_fill_1 FILLER_17_891 ();
 sg13g2_fill_2 FILLER_17_926 ();
 sg13g2_fill_1 FILLER_17_959 ();
 sg13g2_fill_2 FILLER_17_993 ();
 sg13g2_fill_1 FILLER_17_1010 ();
 sg13g2_fill_1 FILLER_17_1020 ();
 sg13g2_decap_4 FILLER_17_1045 ();
 sg13g2_fill_1 FILLER_17_1049 ();
 sg13g2_decap_4 FILLER_17_1086 ();
 sg13g2_fill_1 FILLER_17_1090 ();
 sg13g2_decap_4 FILLER_17_1094 ();
 sg13g2_fill_2 FILLER_17_1167 ();
 sg13g2_fill_1 FILLER_17_1217 ();
 sg13g2_fill_2 FILLER_17_1242 ();
 sg13g2_fill_2 FILLER_17_1253 ();
 sg13g2_fill_1 FILLER_17_1255 ();
 sg13g2_fill_2 FILLER_17_1310 ();
 sg13g2_fill_1 FILLER_17_1354 ();
 sg13g2_fill_1 FILLER_17_1364 ();
 sg13g2_fill_1 FILLER_17_1425 ();
 sg13g2_fill_2 FILLER_17_1473 ();
 sg13g2_fill_1 FILLER_17_1491 ();
 sg13g2_fill_1 FILLER_17_1510 ();
 sg13g2_fill_1 FILLER_17_1556 ();
 sg13g2_fill_2 FILLER_17_1562 ();
 sg13g2_fill_1 FILLER_17_1564 ();
 sg13g2_fill_2 FILLER_17_1571 ();
 sg13g2_fill_1 FILLER_17_1573 ();
 sg13g2_decap_4 FILLER_17_1587 ();
 sg13g2_fill_2 FILLER_17_1591 ();
 sg13g2_fill_2 FILLER_17_1623 ();
 sg13g2_fill_1 FILLER_17_1625 ();
 sg13g2_fill_1 FILLER_17_1632 ();
 sg13g2_fill_2 FILLER_17_1659 ();
 sg13g2_fill_1 FILLER_17_1661 ();
 sg13g2_fill_2 FILLER_17_1729 ();
 sg13g2_fill_1 FILLER_17_1741 ();
 sg13g2_fill_1 FILLER_17_1755 ();
 sg13g2_fill_2 FILLER_17_1787 ();
 sg13g2_fill_1 FILLER_17_1865 ();
 sg13g2_fill_2 FILLER_17_1875 ();
 sg13g2_fill_2 FILLER_17_1913 ();
 sg13g2_fill_1 FILLER_17_1915 ();
 sg13g2_decap_8 FILLER_17_1960 ();
 sg13g2_decap_4 FILLER_17_1967 ();
 sg13g2_fill_2 FILLER_17_1971 ();
 sg13g2_fill_2 FILLER_17_2050 ();
 sg13g2_fill_1 FILLER_17_2094 ();
 sg13g2_fill_2 FILLER_17_2125 ();
 sg13g2_fill_1 FILLER_17_2143 ();
 sg13g2_fill_2 FILLER_17_2155 ();
 sg13g2_fill_1 FILLER_17_2202 ();
 sg13g2_decap_8 FILLER_17_2236 ();
 sg13g2_decap_8 FILLER_17_2243 ();
 sg13g2_decap_8 FILLER_17_2250 ();
 sg13g2_decap_8 FILLER_17_2257 ();
 sg13g2_decap_8 FILLER_17_2264 ();
 sg13g2_decap_8 FILLER_17_2271 ();
 sg13g2_decap_8 FILLER_17_2278 ();
 sg13g2_decap_8 FILLER_17_2285 ();
 sg13g2_decap_8 FILLER_17_2292 ();
 sg13g2_decap_8 FILLER_17_2299 ();
 sg13g2_decap_8 FILLER_17_2306 ();
 sg13g2_decap_8 FILLER_17_2313 ();
 sg13g2_decap_8 FILLER_17_2320 ();
 sg13g2_decap_8 FILLER_17_2327 ();
 sg13g2_decap_8 FILLER_17_2334 ();
 sg13g2_decap_8 FILLER_17_2341 ();
 sg13g2_decap_8 FILLER_17_2348 ();
 sg13g2_decap_8 FILLER_17_2355 ();
 sg13g2_decap_8 FILLER_17_2362 ();
 sg13g2_decap_8 FILLER_17_2369 ();
 sg13g2_decap_8 FILLER_17_2376 ();
 sg13g2_decap_8 FILLER_17_2383 ();
 sg13g2_decap_8 FILLER_17_2390 ();
 sg13g2_decap_8 FILLER_17_2397 ();
 sg13g2_decap_8 FILLER_17_2404 ();
 sg13g2_decap_8 FILLER_17_2411 ();
 sg13g2_decap_8 FILLER_17_2418 ();
 sg13g2_decap_8 FILLER_17_2425 ();
 sg13g2_decap_8 FILLER_17_2432 ();
 sg13g2_decap_8 FILLER_17_2439 ();
 sg13g2_decap_8 FILLER_17_2446 ();
 sg13g2_decap_8 FILLER_17_2453 ();
 sg13g2_decap_8 FILLER_17_2460 ();
 sg13g2_decap_8 FILLER_17_2467 ();
 sg13g2_decap_8 FILLER_17_2474 ();
 sg13g2_decap_8 FILLER_17_2481 ();
 sg13g2_decap_8 FILLER_17_2488 ();
 sg13g2_decap_8 FILLER_17_2495 ();
 sg13g2_decap_8 FILLER_17_2502 ();
 sg13g2_decap_8 FILLER_17_2509 ();
 sg13g2_decap_8 FILLER_17_2516 ();
 sg13g2_decap_8 FILLER_17_2523 ();
 sg13g2_decap_8 FILLER_17_2530 ();
 sg13g2_decap_8 FILLER_17_2537 ();
 sg13g2_decap_8 FILLER_17_2544 ();
 sg13g2_decap_8 FILLER_17_2551 ();
 sg13g2_decap_8 FILLER_17_2558 ();
 sg13g2_decap_8 FILLER_17_2565 ();
 sg13g2_decap_8 FILLER_17_2572 ();
 sg13g2_decap_8 FILLER_17_2579 ();
 sg13g2_decap_8 FILLER_17_2586 ();
 sg13g2_decap_8 FILLER_17_2593 ();
 sg13g2_decap_8 FILLER_17_2600 ();
 sg13g2_decap_8 FILLER_17_2607 ();
 sg13g2_decap_8 FILLER_17_2614 ();
 sg13g2_decap_8 FILLER_17_2621 ();
 sg13g2_decap_8 FILLER_17_2628 ();
 sg13g2_decap_8 FILLER_17_2635 ();
 sg13g2_decap_8 FILLER_17_2642 ();
 sg13g2_decap_8 FILLER_17_2649 ();
 sg13g2_decap_8 FILLER_17_2656 ();
 sg13g2_decap_8 FILLER_17_2663 ();
 sg13g2_decap_4 FILLER_17_2670 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_decap_4 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_2 FILLER_18_305 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_4 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_2 FILLER_18_398 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_decap_4 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_460 ();
 sg13g2_decap_8 FILLER_18_467 ();
 sg13g2_decap_4 FILLER_18_474 ();
 sg13g2_decap_8 FILLER_18_500 ();
 sg13g2_decap_8 FILLER_18_517 ();
 sg13g2_decap_4 FILLER_18_524 ();
 sg13g2_fill_2 FILLER_18_528 ();
 sg13g2_decap_8 FILLER_18_551 ();
 sg13g2_decap_8 FILLER_18_558 ();
 sg13g2_decap_8 FILLER_18_565 ();
 sg13g2_decap_4 FILLER_18_572 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_fill_1 FILLER_18_602 ();
 sg13g2_fill_1 FILLER_18_608 ();
 sg13g2_fill_1 FILLER_18_627 ();
 sg13g2_decap_4 FILLER_18_633 ();
 sg13g2_fill_1 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_642 ();
 sg13g2_decap_8 FILLER_18_649 ();
 sg13g2_fill_2 FILLER_18_656 ();
 sg13g2_fill_1 FILLER_18_658 ();
 sg13g2_fill_2 FILLER_18_669 ();
 sg13g2_fill_1 FILLER_18_671 ();
 sg13g2_fill_1 FILLER_18_687 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_fill_2 FILLER_18_700 ();
 sg13g2_fill_1 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_733 ();
 sg13g2_fill_2 FILLER_18_740 ();
 sg13g2_fill_1 FILLER_18_742 ();
 sg13g2_fill_1 FILLER_18_748 ();
 sg13g2_fill_1 FILLER_18_756 ();
 sg13g2_fill_1 FILLER_18_771 ();
 sg13g2_fill_2 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_fill_1 FILLER_18_840 ();
 sg13g2_fill_2 FILLER_18_844 ();
 sg13g2_fill_1 FILLER_18_846 ();
 sg13g2_decap_4 FILLER_18_853 ();
 sg13g2_fill_2 FILLER_18_961 ();
 sg13g2_fill_1 FILLER_18_976 ();
 sg13g2_fill_2 FILLER_18_983 ();
 sg13g2_decap_8 FILLER_18_1047 ();
 sg13g2_fill_2 FILLER_18_1054 ();
 sg13g2_fill_1 FILLER_18_1056 ();
 sg13g2_decap_4 FILLER_18_1096 ();
 sg13g2_fill_2 FILLER_18_1153 ();
 sg13g2_fill_1 FILLER_18_1155 ();
 sg13g2_fill_2 FILLER_18_1174 ();
 sg13g2_fill_1 FILLER_18_1176 ();
 sg13g2_fill_2 FILLER_18_1297 ();
 sg13g2_fill_2 FILLER_18_1335 ();
 sg13g2_fill_2 FILLER_18_1382 ();
 sg13g2_fill_1 FILLER_18_1458 ();
 sg13g2_fill_2 FILLER_18_1486 ();
 sg13g2_fill_1 FILLER_18_1488 ();
 sg13g2_decap_8 FILLER_18_1595 ();
 sg13g2_decap_4 FILLER_18_1602 ();
 sg13g2_fill_1 FILLER_18_1606 ();
 sg13g2_fill_1 FILLER_18_1642 ();
 sg13g2_fill_1 FILLER_18_1660 ();
 sg13g2_fill_2 FILLER_18_1752 ();
 sg13g2_fill_1 FILLER_18_1754 ();
 sg13g2_fill_2 FILLER_18_1825 ();
 sg13g2_fill_2 FILLER_18_1831 ();
 sg13g2_fill_1 FILLER_18_1833 ();
 sg13g2_fill_2 FILLER_18_1861 ();
 sg13g2_fill_1 FILLER_18_1863 ();
 sg13g2_fill_2 FILLER_18_1929 ();
 sg13g2_decap_8 FILLER_18_1959 ();
 sg13g2_decap_4 FILLER_18_1966 ();
 sg13g2_fill_2 FILLER_18_2024 ();
 sg13g2_fill_1 FILLER_18_2026 ();
 sg13g2_fill_1 FILLER_18_2055 ();
 sg13g2_fill_2 FILLER_18_2069 ();
 sg13g2_fill_2 FILLER_18_2110 ();
 sg13g2_fill_1 FILLER_18_2153 ();
 sg13g2_fill_1 FILLER_18_2158 ();
 sg13g2_fill_1 FILLER_18_2210 ();
 sg13g2_decap_8 FILLER_18_2239 ();
 sg13g2_decap_8 FILLER_18_2246 ();
 sg13g2_decap_8 FILLER_18_2253 ();
 sg13g2_decap_8 FILLER_18_2260 ();
 sg13g2_decap_8 FILLER_18_2267 ();
 sg13g2_decap_8 FILLER_18_2274 ();
 sg13g2_decap_8 FILLER_18_2281 ();
 sg13g2_decap_8 FILLER_18_2288 ();
 sg13g2_decap_8 FILLER_18_2295 ();
 sg13g2_decap_8 FILLER_18_2302 ();
 sg13g2_decap_8 FILLER_18_2309 ();
 sg13g2_decap_8 FILLER_18_2316 ();
 sg13g2_decap_8 FILLER_18_2323 ();
 sg13g2_decap_8 FILLER_18_2330 ();
 sg13g2_decap_8 FILLER_18_2337 ();
 sg13g2_decap_8 FILLER_18_2344 ();
 sg13g2_decap_8 FILLER_18_2351 ();
 sg13g2_decap_8 FILLER_18_2358 ();
 sg13g2_decap_8 FILLER_18_2365 ();
 sg13g2_decap_8 FILLER_18_2372 ();
 sg13g2_decap_8 FILLER_18_2379 ();
 sg13g2_decap_8 FILLER_18_2386 ();
 sg13g2_decap_8 FILLER_18_2393 ();
 sg13g2_decap_8 FILLER_18_2400 ();
 sg13g2_decap_8 FILLER_18_2407 ();
 sg13g2_decap_8 FILLER_18_2414 ();
 sg13g2_decap_8 FILLER_18_2421 ();
 sg13g2_decap_8 FILLER_18_2428 ();
 sg13g2_decap_8 FILLER_18_2435 ();
 sg13g2_decap_8 FILLER_18_2442 ();
 sg13g2_decap_8 FILLER_18_2449 ();
 sg13g2_decap_8 FILLER_18_2456 ();
 sg13g2_decap_8 FILLER_18_2463 ();
 sg13g2_decap_8 FILLER_18_2470 ();
 sg13g2_decap_8 FILLER_18_2477 ();
 sg13g2_decap_8 FILLER_18_2484 ();
 sg13g2_decap_8 FILLER_18_2491 ();
 sg13g2_decap_8 FILLER_18_2498 ();
 sg13g2_decap_8 FILLER_18_2505 ();
 sg13g2_decap_8 FILLER_18_2512 ();
 sg13g2_decap_8 FILLER_18_2519 ();
 sg13g2_decap_8 FILLER_18_2526 ();
 sg13g2_decap_8 FILLER_18_2533 ();
 sg13g2_decap_8 FILLER_18_2540 ();
 sg13g2_decap_8 FILLER_18_2547 ();
 sg13g2_decap_8 FILLER_18_2554 ();
 sg13g2_decap_8 FILLER_18_2561 ();
 sg13g2_decap_8 FILLER_18_2568 ();
 sg13g2_decap_8 FILLER_18_2575 ();
 sg13g2_decap_8 FILLER_18_2582 ();
 sg13g2_decap_8 FILLER_18_2589 ();
 sg13g2_decap_8 FILLER_18_2596 ();
 sg13g2_decap_8 FILLER_18_2603 ();
 sg13g2_decap_8 FILLER_18_2610 ();
 sg13g2_decap_8 FILLER_18_2617 ();
 sg13g2_decap_8 FILLER_18_2624 ();
 sg13g2_decap_8 FILLER_18_2631 ();
 sg13g2_decap_8 FILLER_18_2638 ();
 sg13g2_decap_8 FILLER_18_2645 ();
 sg13g2_decap_8 FILLER_18_2652 ();
 sg13g2_decap_8 FILLER_18_2659 ();
 sg13g2_decap_8 FILLER_18_2666 ();
 sg13g2_fill_1 FILLER_18_2673 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_decap_4 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_decap_4 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_399 ();
 sg13g2_fill_1 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_19_433 ();
 sg13g2_fill_1 FILLER_19_440 ();
 sg13g2_decap_4 FILLER_19_454 ();
 sg13g2_fill_2 FILLER_19_458 ();
 sg13g2_decap_8 FILLER_19_473 ();
 sg13g2_decap_4 FILLER_19_480 ();
 sg13g2_fill_1 FILLER_19_484 ();
 sg13g2_fill_2 FILLER_19_490 ();
 sg13g2_fill_1 FILLER_19_492 ();
 sg13g2_decap_4 FILLER_19_498 ();
 sg13g2_fill_1 FILLER_19_502 ();
 sg13g2_decap_4 FILLER_19_518 ();
 sg13g2_fill_2 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_555 ();
 sg13g2_fill_2 FILLER_19_583 ();
 sg13g2_decap_8 FILLER_19_589 ();
 sg13g2_fill_1 FILLER_19_596 ();
 sg13g2_fill_2 FILLER_19_616 ();
 sg13g2_fill_1 FILLER_19_618 ();
 sg13g2_fill_1 FILLER_19_632 ();
 sg13g2_fill_2 FILLER_19_638 ();
 sg13g2_decap_4 FILLER_19_660 ();
 sg13g2_fill_2 FILLER_19_664 ();
 sg13g2_fill_2 FILLER_19_692 ();
 sg13g2_fill_1 FILLER_19_694 ();
 sg13g2_fill_2 FILLER_19_742 ();
 sg13g2_fill_1 FILLER_19_744 ();
 sg13g2_fill_1 FILLER_19_786 ();
 sg13g2_fill_1 FILLER_19_819 ();
 sg13g2_decap_4 FILLER_19_848 ();
 sg13g2_fill_2 FILLER_19_885 ();
 sg13g2_fill_2 FILLER_19_899 ();
 sg13g2_fill_2 FILLER_19_956 ();
 sg13g2_fill_1 FILLER_19_958 ();
 sg13g2_fill_1 FILLER_19_1012 ();
 sg13g2_decap_4 FILLER_19_1088 ();
 sg13g2_fill_2 FILLER_19_1218 ();
 sg13g2_fill_1 FILLER_19_1220 ();
 sg13g2_fill_2 FILLER_19_1246 ();
 sg13g2_fill_2 FILLER_19_1276 ();
 sg13g2_fill_1 FILLER_19_1278 ();
 sg13g2_fill_2 FILLER_19_1298 ();
 sg13g2_fill_1 FILLER_19_1300 ();
 sg13g2_fill_1 FILLER_19_1317 ();
 sg13g2_fill_1 FILLER_19_1364 ();
 sg13g2_fill_2 FILLER_19_1384 ();
 sg13g2_decap_4 FILLER_19_1408 ();
 sg13g2_fill_2 FILLER_19_1412 ();
 sg13g2_fill_2 FILLER_19_1469 ();
 sg13g2_fill_1 FILLER_19_1496 ();
 sg13g2_decap_8 FILLER_19_1575 ();
 sg13g2_decap_4 FILLER_19_1582 ();
 sg13g2_decap_8 FILLER_19_1594 ();
 sg13g2_fill_1 FILLER_19_1601 ();
 sg13g2_decap_8 FILLER_19_1608 ();
 sg13g2_fill_2 FILLER_19_1620 ();
 sg13g2_decap_4 FILLER_19_1650 ();
 sg13g2_fill_1 FILLER_19_1654 ();
 sg13g2_fill_2 FILLER_19_1687 ();
 sg13g2_fill_1 FILLER_19_1689 ();
 sg13g2_fill_2 FILLER_19_1829 ();
 sg13g2_fill_1 FILLER_19_1911 ();
 sg13g2_fill_2 FILLER_19_1953 ();
 sg13g2_fill_1 FILLER_19_1955 ();
 sg13g2_decap_8 FILLER_19_1965 ();
 sg13g2_fill_2 FILLER_19_1972 ();
 sg13g2_fill_1 FILLER_19_2021 ();
 sg13g2_fill_2 FILLER_19_2040 ();
 sg13g2_fill_1 FILLER_19_2042 ();
 sg13g2_decap_8 FILLER_19_2071 ();
 sg13g2_fill_2 FILLER_19_2206 ();
 sg13g2_fill_1 FILLER_19_2222 ();
 sg13g2_decap_8 FILLER_19_2241 ();
 sg13g2_decap_8 FILLER_19_2248 ();
 sg13g2_decap_8 FILLER_19_2255 ();
 sg13g2_decap_8 FILLER_19_2262 ();
 sg13g2_decap_8 FILLER_19_2269 ();
 sg13g2_decap_8 FILLER_19_2276 ();
 sg13g2_decap_8 FILLER_19_2283 ();
 sg13g2_decap_8 FILLER_19_2290 ();
 sg13g2_decap_8 FILLER_19_2297 ();
 sg13g2_decap_8 FILLER_19_2304 ();
 sg13g2_decap_8 FILLER_19_2311 ();
 sg13g2_decap_8 FILLER_19_2318 ();
 sg13g2_decap_8 FILLER_19_2325 ();
 sg13g2_decap_8 FILLER_19_2332 ();
 sg13g2_decap_8 FILLER_19_2339 ();
 sg13g2_decap_8 FILLER_19_2346 ();
 sg13g2_decap_8 FILLER_19_2353 ();
 sg13g2_decap_8 FILLER_19_2360 ();
 sg13g2_decap_8 FILLER_19_2367 ();
 sg13g2_decap_8 FILLER_19_2374 ();
 sg13g2_decap_8 FILLER_19_2381 ();
 sg13g2_decap_8 FILLER_19_2388 ();
 sg13g2_decap_8 FILLER_19_2395 ();
 sg13g2_decap_8 FILLER_19_2402 ();
 sg13g2_decap_8 FILLER_19_2409 ();
 sg13g2_decap_8 FILLER_19_2416 ();
 sg13g2_decap_8 FILLER_19_2423 ();
 sg13g2_decap_8 FILLER_19_2430 ();
 sg13g2_decap_8 FILLER_19_2437 ();
 sg13g2_decap_8 FILLER_19_2444 ();
 sg13g2_decap_8 FILLER_19_2451 ();
 sg13g2_decap_8 FILLER_19_2458 ();
 sg13g2_decap_8 FILLER_19_2465 ();
 sg13g2_decap_8 FILLER_19_2472 ();
 sg13g2_decap_8 FILLER_19_2479 ();
 sg13g2_decap_8 FILLER_19_2486 ();
 sg13g2_decap_8 FILLER_19_2493 ();
 sg13g2_decap_8 FILLER_19_2500 ();
 sg13g2_decap_8 FILLER_19_2507 ();
 sg13g2_decap_8 FILLER_19_2514 ();
 sg13g2_decap_8 FILLER_19_2521 ();
 sg13g2_decap_8 FILLER_19_2528 ();
 sg13g2_decap_8 FILLER_19_2535 ();
 sg13g2_decap_8 FILLER_19_2542 ();
 sg13g2_decap_8 FILLER_19_2549 ();
 sg13g2_decap_8 FILLER_19_2556 ();
 sg13g2_decap_8 FILLER_19_2563 ();
 sg13g2_decap_8 FILLER_19_2570 ();
 sg13g2_decap_8 FILLER_19_2577 ();
 sg13g2_decap_8 FILLER_19_2584 ();
 sg13g2_decap_8 FILLER_19_2591 ();
 sg13g2_decap_8 FILLER_19_2598 ();
 sg13g2_decap_8 FILLER_19_2605 ();
 sg13g2_decap_8 FILLER_19_2612 ();
 sg13g2_decap_8 FILLER_19_2619 ();
 sg13g2_decap_8 FILLER_19_2626 ();
 sg13g2_decap_8 FILLER_19_2633 ();
 sg13g2_decap_8 FILLER_19_2640 ();
 sg13g2_decap_8 FILLER_19_2647 ();
 sg13g2_decap_8 FILLER_19_2654 ();
 sg13g2_decap_8 FILLER_19_2661 ();
 sg13g2_decap_4 FILLER_19_2668 ();
 sg13g2_fill_2 FILLER_19_2672 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_26 ();
 sg13g2_fill_2 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_105 ();
 sg13g2_decap_4 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_232 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_412 ();
 sg13g2_fill_2 FILLER_20_440 ();
 sg13g2_fill_1 FILLER_20_442 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_4 FILLER_20_455 ();
 sg13g2_fill_2 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_489 ();
 sg13g2_decap_8 FILLER_20_496 ();
 sg13g2_fill_2 FILLER_20_503 ();
 sg13g2_fill_1 FILLER_20_514 ();
 sg13g2_fill_2 FILLER_20_519 ();
 sg13g2_fill_1 FILLER_20_535 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_fill_1 FILLER_20_582 ();
 sg13g2_decap_4 FILLER_20_593 ();
 sg13g2_fill_1 FILLER_20_597 ();
 sg13g2_decap_8 FILLER_20_611 ();
 sg13g2_decap_8 FILLER_20_618 ();
 sg13g2_decap_8 FILLER_20_625 ();
 sg13g2_decap_8 FILLER_20_632 ();
 sg13g2_decap_8 FILLER_20_639 ();
 sg13g2_decap_4 FILLER_20_646 ();
 sg13g2_fill_1 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_4 FILLER_20_670 ();
 sg13g2_fill_2 FILLER_20_674 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_4 FILLER_20_700 ();
 sg13g2_fill_2 FILLER_20_704 ();
 sg13g2_decap_4 FILLER_20_737 ();
 sg13g2_fill_1 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_fill_1 FILLER_20_784 ();
 sg13g2_decap_4 FILLER_20_856 ();
 sg13g2_fill_1 FILLER_20_860 ();
 sg13g2_fill_1 FILLER_20_865 ();
 sg13g2_fill_2 FILLER_20_901 ();
 sg13g2_fill_2 FILLER_20_944 ();
 sg13g2_fill_2 FILLER_20_992 ();
 sg13g2_fill_2 FILLER_20_1002 ();
 sg13g2_fill_2 FILLER_20_1015 ();
 sg13g2_decap_8 FILLER_20_1036 ();
 sg13g2_fill_2 FILLER_20_1043 ();
 sg13g2_fill_1 FILLER_20_1079 ();
 sg13g2_fill_2 FILLER_20_1106 ();
 sg13g2_fill_2 FILLER_20_1206 ();
 sg13g2_fill_2 FILLER_20_1270 ();
 sg13g2_fill_1 FILLER_20_1272 ();
 sg13g2_fill_1 FILLER_20_1278 ();
 sg13g2_fill_2 FILLER_20_1321 ();
 sg13g2_fill_1 FILLER_20_1323 ();
 sg13g2_fill_1 FILLER_20_1376 ();
 sg13g2_fill_1 FILLER_20_1392 ();
 sg13g2_decap_8 FILLER_20_1406 ();
 sg13g2_fill_2 FILLER_20_1413 ();
 sg13g2_fill_1 FILLER_20_1425 ();
 sg13g2_decap_8 FILLER_20_1547 ();
 sg13g2_fill_2 FILLER_20_1554 ();
 sg13g2_decap_8 FILLER_20_1575 ();
 sg13g2_decap_8 FILLER_20_1582 ();
 sg13g2_decap_8 FILLER_20_1589 ();
 sg13g2_fill_1 FILLER_20_1596 ();
 sg13g2_fill_2 FILLER_20_1604 ();
 sg13g2_fill_2 FILLER_20_1628 ();
 sg13g2_fill_1 FILLER_20_1697 ();
 sg13g2_fill_1 FILLER_20_1705 ();
 sg13g2_fill_2 FILLER_20_1714 ();
 sg13g2_fill_1 FILLER_20_1716 ();
 sg13g2_fill_2 FILLER_20_1728 ();
 sg13g2_fill_1 FILLER_20_1768 ();
 sg13g2_fill_1 FILLER_20_1815 ();
 sg13g2_fill_1 FILLER_20_1905 ();
 sg13g2_fill_2 FILLER_20_1915 ();
 sg13g2_fill_1 FILLER_20_1917 ();
 sg13g2_decap_4 FILLER_20_1964 ();
 sg13g2_fill_2 FILLER_20_1968 ();
 sg13g2_fill_2 FILLER_20_1997 ();
 sg13g2_fill_2 FILLER_20_2017 ();
 sg13g2_fill_1 FILLER_20_2019 ();
 sg13g2_fill_2 FILLER_20_2096 ();
 sg13g2_fill_2 FILLER_20_2143 ();
 sg13g2_fill_2 FILLER_20_2155 ();
 sg13g2_fill_1 FILLER_20_2166 ();
 sg13g2_fill_2 FILLER_20_2208 ();
 sg13g2_fill_1 FILLER_20_2210 ();
 sg13g2_decap_8 FILLER_20_2224 ();
 sg13g2_decap_4 FILLER_20_2231 ();
 sg13g2_decap_8 FILLER_20_2244 ();
 sg13g2_decap_8 FILLER_20_2251 ();
 sg13g2_decap_8 FILLER_20_2258 ();
 sg13g2_decap_8 FILLER_20_2265 ();
 sg13g2_decap_8 FILLER_20_2272 ();
 sg13g2_decap_8 FILLER_20_2279 ();
 sg13g2_decap_8 FILLER_20_2286 ();
 sg13g2_decap_8 FILLER_20_2293 ();
 sg13g2_decap_8 FILLER_20_2300 ();
 sg13g2_decap_8 FILLER_20_2307 ();
 sg13g2_decap_8 FILLER_20_2314 ();
 sg13g2_decap_8 FILLER_20_2321 ();
 sg13g2_decap_8 FILLER_20_2328 ();
 sg13g2_decap_8 FILLER_20_2335 ();
 sg13g2_decap_8 FILLER_20_2342 ();
 sg13g2_decap_8 FILLER_20_2349 ();
 sg13g2_decap_8 FILLER_20_2356 ();
 sg13g2_decap_8 FILLER_20_2363 ();
 sg13g2_decap_8 FILLER_20_2370 ();
 sg13g2_decap_8 FILLER_20_2377 ();
 sg13g2_decap_8 FILLER_20_2384 ();
 sg13g2_decap_8 FILLER_20_2391 ();
 sg13g2_decap_8 FILLER_20_2398 ();
 sg13g2_decap_8 FILLER_20_2405 ();
 sg13g2_decap_8 FILLER_20_2412 ();
 sg13g2_decap_8 FILLER_20_2419 ();
 sg13g2_decap_8 FILLER_20_2426 ();
 sg13g2_decap_8 FILLER_20_2433 ();
 sg13g2_decap_8 FILLER_20_2440 ();
 sg13g2_decap_8 FILLER_20_2447 ();
 sg13g2_decap_8 FILLER_20_2454 ();
 sg13g2_decap_8 FILLER_20_2461 ();
 sg13g2_decap_8 FILLER_20_2468 ();
 sg13g2_decap_8 FILLER_20_2475 ();
 sg13g2_decap_8 FILLER_20_2482 ();
 sg13g2_decap_8 FILLER_20_2489 ();
 sg13g2_decap_8 FILLER_20_2496 ();
 sg13g2_decap_8 FILLER_20_2503 ();
 sg13g2_decap_8 FILLER_20_2510 ();
 sg13g2_decap_8 FILLER_20_2517 ();
 sg13g2_decap_8 FILLER_20_2524 ();
 sg13g2_decap_8 FILLER_20_2531 ();
 sg13g2_decap_8 FILLER_20_2538 ();
 sg13g2_decap_8 FILLER_20_2545 ();
 sg13g2_decap_8 FILLER_20_2552 ();
 sg13g2_decap_8 FILLER_20_2559 ();
 sg13g2_decap_8 FILLER_20_2566 ();
 sg13g2_decap_8 FILLER_20_2573 ();
 sg13g2_decap_8 FILLER_20_2580 ();
 sg13g2_decap_8 FILLER_20_2587 ();
 sg13g2_decap_8 FILLER_20_2594 ();
 sg13g2_decap_8 FILLER_20_2601 ();
 sg13g2_decap_8 FILLER_20_2608 ();
 sg13g2_decap_8 FILLER_20_2615 ();
 sg13g2_decap_8 FILLER_20_2622 ();
 sg13g2_decap_8 FILLER_20_2629 ();
 sg13g2_decap_8 FILLER_20_2636 ();
 sg13g2_decap_8 FILLER_20_2643 ();
 sg13g2_decap_8 FILLER_20_2650 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_8 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2671 ();
 sg13g2_fill_1 FILLER_20_2673 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_9 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_96 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_decap_4 FILLER_21_132 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_399 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_21_430 ();
 sg13g2_fill_1 FILLER_21_459 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_fill_2 FILLER_21_508 ();
 sg13g2_fill_1 FILLER_21_516 ();
 sg13g2_fill_2 FILLER_21_540 ();
 sg13g2_fill_2 FILLER_21_560 ();
 sg13g2_fill_1 FILLER_21_562 ();
 sg13g2_decap_4 FILLER_21_581 ();
 sg13g2_fill_1 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_608 ();
 sg13g2_decap_8 FILLER_21_615 ();
 sg13g2_decap_8 FILLER_21_622 ();
 sg13g2_decap_8 FILLER_21_629 ();
 sg13g2_decap_4 FILLER_21_636 ();
 sg13g2_fill_1 FILLER_21_640 ();
 sg13g2_decap_8 FILLER_21_661 ();
 sg13g2_decap_4 FILLER_21_668 ();
 sg13g2_fill_1 FILLER_21_672 ();
 sg13g2_decap_4 FILLER_21_683 ();
 sg13g2_fill_1 FILLER_21_687 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_fill_2 FILLER_21_719 ();
 sg13g2_fill_1 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_739 ();
 sg13g2_decap_4 FILLER_21_746 ();
 sg13g2_decap_4 FILLER_21_768 ();
 sg13g2_fill_2 FILLER_21_772 ();
 sg13g2_decap_4 FILLER_21_780 ();
 sg13g2_fill_2 FILLER_21_903 ();
 sg13g2_decap_4 FILLER_21_912 ();
 sg13g2_fill_2 FILLER_21_916 ();
 sg13g2_decap_8 FILLER_21_936 ();
 sg13g2_fill_2 FILLER_21_943 ();
 sg13g2_fill_2 FILLER_21_960 ();
 sg13g2_fill_2 FILLER_21_975 ();
 sg13g2_fill_1 FILLER_21_977 ();
 sg13g2_fill_1 FILLER_21_981 ();
 sg13g2_fill_1 FILLER_21_1035 ();
 sg13g2_fill_1 FILLER_21_1094 ();
 sg13g2_fill_2 FILLER_21_1101 ();
 sg13g2_fill_2 FILLER_21_1120 ();
 sg13g2_fill_1 FILLER_21_1122 ();
 sg13g2_fill_2 FILLER_21_1148 ();
 sg13g2_fill_1 FILLER_21_1159 ();
 sg13g2_fill_2 FILLER_21_1211 ();
 sg13g2_fill_1 FILLER_21_1268 ();
 sg13g2_fill_1 FILLER_21_1283 ();
 sg13g2_fill_2 FILLER_21_1297 ();
 sg13g2_fill_1 FILLER_21_1377 ();
 sg13g2_decap_8 FILLER_21_1398 ();
 sg13g2_decap_4 FILLER_21_1405 ();
 sg13g2_fill_2 FILLER_21_1460 ();
 sg13g2_fill_1 FILLER_21_1462 ();
 sg13g2_fill_2 FILLER_21_1468 ();
 sg13g2_fill_1 FILLER_21_1495 ();
 sg13g2_fill_2 FILLER_21_1511 ();
 sg13g2_fill_1 FILLER_21_1513 ();
 sg13g2_decap_4 FILLER_21_1537 ();
 sg13g2_decap_8 FILLER_21_1554 ();
 sg13g2_fill_2 FILLER_21_1595 ();
 sg13g2_fill_2 FILLER_21_1601 ();
 sg13g2_fill_1 FILLER_21_1603 ();
 sg13g2_fill_2 FILLER_21_1631 ();
 sg13g2_fill_1 FILLER_21_1633 ();
 sg13g2_fill_1 FILLER_21_1652 ();
 sg13g2_fill_1 FILLER_21_1716 ();
 sg13g2_fill_2 FILLER_21_1767 ();
 sg13g2_fill_1 FILLER_21_1769 ();
 sg13g2_fill_1 FILLER_21_1779 ();
 sg13g2_fill_2 FILLER_21_1809 ();
 sg13g2_fill_1 FILLER_21_1848 ();
 sg13g2_fill_2 FILLER_21_1858 ();
 sg13g2_fill_2 FILLER_21_1914 ();
 sg13g2_fill_2 FILLER_21_1970 ();
 sg13g2_fill_1 FILLER_21_1972 ();
 sg13g2_fill_1 FILLER_21_2017 ();
 sg13g2_fill_2 FILLER_21_2048 ();
 sg13g2_decap_4 FILLER_21_2103 ();
 sg13g2_fill_2 FILLER_21_2164 ();
 sg13g2_fill_2 FILLER_21_2199 ();
 sg13g2_decap_8 FILLER_21_2248 ();
 sg13g2_decap_8 FILLER_21_2255 ();
 sg13g2_decap_8 FILLER_21_2262 ();
 sg13g2_decap_8 FILLER_21_2269 ();
 sg13g2_decap_8 FILLER_21_2276 ();
 sg13g2_decap_8 FILLER_21_2283 ();
 sg13g2_decap_8 FILLER_21_2290 ();
 sg13g2_decap_8 FILLER_21_2297 ();
 sg13g2_decap_8 FILLER_21_2304 ();
 sg13g2_decap_8 FILLER_21_2311 ();
 sg13g2_decap_8 FILLER_21_2318 ();
 sg13g2_decap_8 FILLER_21_2325 ();
 sg13g2_decap_8 FILLER_21_2332 ();
 sg13g2_decap_8 FILLER_21_2339 ();
 sg13g2_decap_8 FILLER_21_2346 ();
 sg13g2_decap_8 FILLER_21_2353 ();
 sg13g2_decap_8 FILLER_21_2360 ();
 sg13g2_decap_8 FILLER_21_2367 ();
 sg13g2_decap_8 FILLER_21_2374 ();
 sg13g2_decap_8 FILLER_21_2381 ();
 sg13g2_decap_8 FILLER_21_2388 ();
 sg13g2_decap_8 FILLER_21_2395 ();
 sg13g2_decap_8 FILLER_21_2402 ();
 sg13g2_decap_8 FILLER_21_2409 ();
 sg13g2_decap_8 FILLER_21_2416 ();
 sg13g2_decap_8 FILLER_21_2423 ();
 sg13g2_decap_8 FILLER_21_2430 ();
 sg13g2_decap_8 FILLER_21_2437 ();
 sg13g2_decap_8 FILLER_21_2444 ();
 sg13g2_decap_8 FILLER_21_2451 ();
 sg13g2_decap_8 FILLER_21_2458 ();
 sg13g2_decap_8 FILLER_21_2465 ();
 sg13g2_decap_8 FILLER_21_2472 ();
 sg13g2_decap_8 FILLER_21_2479 ();
 sg13g2_decap_8 FILLER_21_2486 ();
 sg13g2_decap_8 FILLER_21_2493 ();
 sg13g2_decap_8 FILLER_21_2500 ();
 sg13g2_decap_8 FILLER_21_2507 ();
 sg13g2_decap_8 FILLER_21_2514 ();
 sg13g2_decap_8 FILLER_21_2521 ();
 sg13g2_decap_8 FILLER_21_2528 ();
 sg13g2_decap_8 FILLER_21_2535 ();
 sg13g2_decap_8 FILLER_21_2542 ();
 sg13g2_decap_8 FILLER_21_2549 ();
 sg13g2_decap_8 FILLER_21_2556 ();
 sg13g2_decap_8 FILLER_21_2563 ();
 sg13g2_decap_8 FILLER_21_2570 ();
 sg13g2_decap_8 FILLER_21_2577 ();
 sg13g2_decap_8 FILLER_21_2584 ();
 sg13g2_decap_8 FILLER_21_2591 ();
 sg13g2_decap_8 FILLER_21_2598 ();
 sg13g2_decap_8 FILLER_21_2605 ();
 sg13g2_decap_8 FILLER_21_2612 ();
 sg13g2_decap_8 FILLER_21_2619 ();
 sg13g2_decap_8 FILLER_21_2626 ();
 sg13g2_decap_8 FILLER_21_2633 ();
 sg13g2_decap_8 FILLER_21_2640 ();
 sg13g2_decap_8 FILLER_21_2647 ();
 sg13g2_decap_8 FILLER_21_2654 ();
 sg13g2_decap_8 FILLER_21_2661 ();
 sg13g2_decap_4 FILLER_21_2668 ();
 sg13g2_fill_2 FILLER_21_2672 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_47 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_173 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_2 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_432 ();
 sg13g2_decap_4 FILLER_22_446 ();
 sg13g2_fill_2 FILLER_22_450 ();
 sg13g2_decap_4 FILLER_22_476 ();
 sg13g2_fill_1 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_496 ();
 sg13g2_decap_8 FILLER_22_503 ();
 sg13g2_decap_8 FILLER_22_510 ();
 sg13g2_decap_8 FILLER_22_517 ();
 sg13g2_fill_2 FILLER_22_524 ();
 sg13g2_decap_8 FILLER_22_545 ();
 sg13g2_fill_2 FILLER_22_552 ();
 sg13g2_fill_1 FILLER_22_554 ();
 sg13g2_fill_2 FILLER_22_560 ();
 sg13g2_fill_2 FILLER_22_566 ();
 sg13g2_decap_4 FILLER_22_573 ();
 sg13g2_fill_2 FILLER_22_591 ();
 sg13g2_fill_1 FILLER_22_593 ();
 sg13g2_fill_2 FILLER_22_607 ();
 sg13g2_decap_4 FILLER_22_626 ();
 sg13g2_fill_1 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_636 ();
 sg13g2_decap_4 FILLER_22_643 ();
 sg13g2_fill_2 FILLER_22_660 ();
 sg13g2_decap_8 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_705 ();
 sg13g2_fill_2 FILLER_22_712 ();
 sg13g2_fill_1 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_fill_1 FILLER_22_753 ();
 sg13g2_fill_2 FILLER_22_816 ();
 sg13g2_fill_1 FILLER_22_818 ();
 sg13g2_decap_4 FILLER_22_900 ();
 sg13g2_fill_1 FILLER_22_904 ();
 sg13g2_fill_1 FILLER_22_946 ();
 sg13g2_decap_8 FILLER_22_978 ();
 sg13g2_fill_1 FILLER_22_985 ();
 sg13g2_fill_1 FILLER_22_1034 ();
 sg13g2_fill_2 FILLER_22_1076 ();
 sg13g2_fill_2 FILLER_22_1105 ();
 sg13g2_fill_1 FILLER_22_1107 ();
 sg13g2_fill_1 FILLER_22_1168 ();
 sg13g2_fill_2 FILLER_22_1182 ();
 sg13g2_fill_1 FILLER_22_1249 ();
 sg13g2_fill_2 FILLER_22_1296 ();
 sg13g2_fill_1 FILLER_22_1298 ();
 sg13g2_fill_1 FILLER_22_1307 ();
 sg13g2_decap_4 FILLER_22_1314 ();
 sg13g2_fill_2 FILLER_22_1318 ();
 sg13g2_fill_1 FILLER_22_1337 ();
 sg13g2_fill_1 FILLER_22_1352 ();
 sg13g2_decap_4 FILLER_22_1389 ();
 sg13g2_fill_1 FILLER_22_1406 ();
 sg13g2_fill_2 FILLER_22_1419 ();
 sg13g2_fill_1 FILLER_22_1421 ();
 sg13g2_decap_8 FILLER_22_1440 ();
 sg13g2_decap_8 FILLER_22_1447 ();
 sg13g2_decap_8 FILLER_22_1454 ();
 sg13g2_decap_4 FILLER_22_1461 ();
 sg13g2_fill_2 FILLER_22_1465 ();
 sg13g2_fill_2 FILLER_22_1499 ();
 sg13g2_fill_2 FILLER_22_1525 ();
 sg13g2_fill_1 FILLER_22_1527 ();
 sg13g2_decap_4 FILLER_22_1541 ();
 sg13g2_fill_1 FILLER_22_1545 ();
 sg13g2_fill_2 FILLER_22_1564 ();
 sg13g2_fill_2 FILLER_22_1572 ();
 sg13g2_fill_2 FILLER_22_1591 ();
 sg13g2_fill_2 FILLER_22_1625 ();
 sg13g2_decap_4 FILLER_22_1677 ();
 sg13g2_fill_1 FILLER_22_1708 ();
 sg13g2_fill_2 FILLER_22_1748 ();
 sg13g2_fill_1 FILLER_22_1800 ();
 sg13g2_fill_2 FILLER_22_1833 ();
 sg13g2_fill_2 FILLER_22_1853 ();
 sg13g2_fill_1 FILLER_22_1864 ();
 sg13g2_fill_2 FILLER_22_1878 ();
 sg13g2_fill_1 FILLER_22_1889 ();
 sg13g2_fill_2 FILLER_22_2042 ();
 sg13g2_fill_1 FILLER_22_2044 ();
 sg13g2_fill_1 FILLER_22_2086 ();
 sg13g2_decap_8 FILLER_22_2100 ();
 sg13g2_fill_2 FILLER_22_2107 ();
 sg13g2_fill_1 FILLER_22_2109 ();
 sg13g2_fill_1 FILLER_22_2168 ();
 sg13g2_fill_2 FILLER_22_2184 ();
 sg13g2_fill_2 FILLER_22_2214 ();
 sg13g2_fill_1 FILLER_22_2216 ();
 sg13g2_decap_8 FILLER_22_2245 ();
 sg13g2_decap_8 FILLER_22_2252 ();
 sg13g2_decap_8 FILLER_22_2259 ();
 sg13g2_decap_8 FILLER_22_2266 ();
 sg13g2_decap_8 FILLER_22_2273 ();
 sg13g2_decap_8 FILLER_22_2280 ();
 sg13g2_decap_8 FILLER_22_2287 ();
 sg13g2_decap_8 FILLER_22_2294 ();
 sg13g2_decap_8 FILLER_22_2301 ();
 sg13g2_decap_8 FILLER_22_2308 ();
 sg13g2_decap_8 FILLER_22_2315 ();
 sg13g2_decap_8 FILLER_22_2322 ();
 sg13g2_decap_8 FILLER_22_2329 ();
 sg13g2_decap_8 FILLER_22_2336 ();
 sg13g2_decap_8 FILLER_22_2343 ();
 sg13g2_decap_8 FILLER_22_2350 ();
 sg13g2_decap_8 FILLER_22_2357 ();
 sg13g2_decap_8 FILLER_22_2364 ();
 sg13g2_decap_8 FILLER_22_2371 ();
 sg13g2_decap_8 FILLER_22_2378 ();
 sg13g2_decap_8 FILLER_22_2385 ();
 sg13g2_decap_8 FILLER_22_2392 ();
 sg13g2_decap_8 FILLER_22_2399 ();
 sg13g2_decap_8 FILLER_22_2406 ();
 sg13g2_decap_8 FILLER_22_2413 ();
 sg13g2_decap_8 FILLER_22_2420 ();
 sg13g2_decap_8 FILLER_22_2427 ();
 sg13g2_decap_8 FILLER_22_2434 ();
 sg13g2_decap_8 FILLER_22_2441 ();
 sg13g2_decap_8 FILLER_22_2448 ();
 sg13g2_decap_8 FILLER_22_2455 ();
 sg13g2_decap_8 FILLER_22_2462 ();
 sg13g2_decap_8 FILLER_22_2469 ();
 sg13g2_decap_8 FILLER_22_2476 ();
 sg13g2_decap_8 FILLER_22_2483 ();
 sg13g2_decap_8 FILLER_22_2490 ();
 sg13g2_decap_8 FILLER_22_2497 ();
 sg13g2_decap_8 FILLER_22_2504 ();
 sg13g2_decap_8 FILLER_22_2511 ();
 sg13g2_decap_8 FILLER_22_2518 ();
 sg13g2_decap_8 FILLER_22_2525 ();
 sg13g2_decap_8 FILLER_22_2532 ();
 sg13g2_decap_8 FILLER_22_2539 ();
 sg13g2_decap_8 FILLER_22_2546 ();
 sg13g2_decap_8 FILLER_22_2553 ();
 sg13g2_decap_8 FILLER_22_2560 ();
 sg13g2_decap_8 FILLER_22_2567 ();
 sg13g2_decap_8 FILLER_22_2574 ();
 sg13g2_decap_8 FILLER_22_2581 ();
 sg13g2_decap_8 FILLER_22_2588 ();
 sg13g2_decap_8 FILLER_22_2595 ();
 sg13g2_decap_8 FILLER_22_2602 ();
 sg13g2_decap_8 FILLER_22_2609 ();
 sg13g2_decap_8 FILLER_22_2616 ();
 sg13g2_decap_8 FILLER_22_2623 ();
 sg13g2_decap_8 FILLER_22_2630 ();
 sg13g2_decap_8 FILLER_22_2637 ();
 sg13g2_decap_8 FILLER_22_2644 ();
 sg13g2_decap_8 FILLER_22_2651 ();
 sg13g2_decap_8 FILLER_22_2658 ();
 sg13g2_decap_8 FILLER_22_2665 ();
 sg13g2_fill_2 FILLER_22_2672 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_90 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_2 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_4 FILLER_23_452 ();
 sg13g2_fill_1 FILLER_23_456 ();
 sg13g2_decap_8 FILLER_23_512 ();
 sg13g2_fill_2 FILLER_23_519 ();
 sg13g2_decap_8 FILLER_23_524 ();
 sg13g2_fill_2 FILLER_23_531 ();
 sg13g2_decap_4 FILLER_23_579 ();
 sg13g2_fill_2 FILLER_23_583 ();
 sg13g2_fill_2 FILLER_23_630 ();
 sg13g2_fill_1 FILLER_23_632 ();
 sg13g2_fill_2 FILLER_23_638 ();
 sg13g2_fill_2 FILLER_23_666 ();
 sg13g2_fill_1 FILLER_23_668 ();
 sg13g2_fill_1 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_695 ();
 sg13g2_fill_1 FILLER_23_702 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_743 ();
 sg13g2_fill_2 FILLER_23_804 ();
 sg13g2_fill_2 FILLER_23_819 ();
 sg13g2_fill_1 FILLER_23_878 ();
 sg13g2_decap_8 FILLER_23_897 ();
 sg13g2_decap_8 FILLER_23_904 ();
 sg13g2_decap_4 FILLER_23_911 ();
 sg13g2_fill_1 FILLER_23_915 ();
 sg13g2_decap_8 FILLER_23_980 ();
 sg13g2_decap_4 FILLER_23_987 ();
 sg13g2_fill_1 FILLER_23_1043 ();
 sg13g2_fill_1 FILLER_23_1058 ();
 sg13g2_decap_4 FILLER_23_1083 ();
 sg13g2_fill_1 FILLER_23_1096 ();
 sg13g2_decap_4 FILLER_23_1106 ();
 sg13g2_fill_2 FILLER_23_1110 ();
 sg13g2_fill_2 FILLER_23_1152 ();
 sg13g2_fill_1 FILLER_23_1154 ();
 sg13g2_fill_2 FILLER_23_1196 ();
 sg13g2_fill_1 FILLER_23_1198 ();
 sg13g2_fill_1 FILLER_23_1213 ();
 sg13g2_fill_1 FILLER_23_1229 ();
 sg13g2_fill_1 FILLER_23_1242 ();
 sg13g2_fill_2 FILLER_23_1283 ();
 sg13g2_fill_1 FILLER_23_1285 ();
 sg13g2_decap_8 FILLER_23_1305 ();
 sg13g2_decap_8 FILLER_23_1312 ();
 sg13g2_fill_2 FILLER_23_1319 ();
 sg13g2_fill_1 FILLER_23_1321 ();
 sg13g2_fill_1 FILLER_23_1340 ();
 sg13g2_fill_1 FILLER_23_1357 ();
 sg13g2_decap_4 FILLER_23_1367 ();
 sg13g2_fill_1 FILLER_23_1371 ();
 sg13g2_fill_1 FILLER_23_1377 ();
 sg13g2_fill_2 FILLER_23_1409 ();
 sg13g2_fill_1 FILLER_23_1411 ();
 sg13g2_fill_1 FILLER_23_1516 ();
 sg13g2_fill_2 FILLER_23_1543 ();
 sg13g2_fill_1 FILLER_23_1545 ();
 sg13g2_fill_2 FILLER_23_1611 ();
 sg13g2_fill_1 FILLER_23_1670 ();
 sg13g2_decap_8 FILLER_23_1681 ();
 sg13g2_fill_1 FILLER_23_1729 ();
 sg13g2_fill_1 FILLER_23_1761 ();
 sg13g2_fill_2 FILLER_23_1801 ();
 sg13g2_fill_1 FILLER_23_1803 ();
 sg13g2_fill_2 FILLER_23_1813 ();
 sg13g2_fill_2 FILLER_23_1829 ();
 sg13g2_fill_2 FILLER_23_1840 ();
 sg13g2_decap_4 FILLER_23_1861 ();
 sg13g2_fill_1 FILLER_23_1877 ();
 sg13g2_fill_1 FILLER_23_1883 ();
 sg13g2_fill_2 FILLER_23_1893 ();
 sg13g2_fill_1 FILLER_23_1936 ();
 sg13g2_decap_4 FILLER_23_1959 ();
 sg13g2_fill_1 FILLER_23_1963 ();
 sg13g2_decap_8 FILLER_23_1973 ();
 sg13g2_decap_4 FILLER_23_1980 ();
 sg13g2_fill_1 FILLER_23_1984 ();
 sg13g2_fill_2 FILLER_23_1998 ();
 sg13g2_fill_2 FILLER_23_2009 ();
 sg13g2_fill_1 FILLER_23_2050 ();
 sg13g2_fill_2 FILLER_23_2060 ();
 sg13g2_fill_2 FILLER_23_2121 ();
 sg13g2_fill_1 FILLER_23_2123 ();
 sg13g2_fill_1 FILLER_23_2134 ();
 sg13g2_fill_2 FILLER_23_2169 ();
 sg13g2_fill_1 FILLER_23_2203 ();
 sg13g2_fill_2 FILLER_23_2213 ();
 sg13g2_fill_1 FILLER_23_2215 ();
 sg13g2_fill_2 FILLER_23_2225 ();
 sg13g2_fill_1 FILLER_23_2227 ();
 sg13g2_decap_8 FILLER_23_2241 ();
 sg13g2_decap_8 FILLER_23_2248 ();
 sg13g2_decap_8 FILLER_23_2255 ();
 sg13g2_decap_8 FILLER_23_2262 ();
 sg13g2_decap_8 FILLER_23_2269 ();
 sg13g2_decap_8 FILLER_23_2276 ();
 sg13g2_decap_8 FILLER_23_2283 ();
 sg13g2_decap_8 FILLER_23_2290 ();
 sg13g2_decap_8 FILLER_23_2297 ();
 sg13g2_decap_8 FILLER_23_2304 ();
 sg13g2_decap_8 FILLER_23_2311 ();
 sg13g2_decap_8 FILLER_23_2318 ();
 sg13g2_decap_8 FILLER_23_2325 ();
 sg13g2_decap_8 FILLER_23_2332 ();
 sg13g2_decap_8 FILLER_23_2339 ();
 sg13g2_decap_8 FILLER_23_2346 ();
 sg13g2_decap_8 FILLER_23_2353 ();
 sg13g2_decap_8 FILLER_23_2360 ();
 sg13g2_decap_8 FILLER_23_2367 ();
 sg13g2_decap_8 FILLER_23_2374 ();
 sg13g2_decap_8 FILLER_23_2381 ();
 sg13g2_decap_8 FILLER_23_2388 ();
 sg13g2_decap_8 FILLER_23_2395 ();
 sg13g2_decap_8 FILLER_23_2402 ();
 sg13g2_decap_8 FILLER_23_2409 ();
 sg13g2_decap_8 FILLER_23_2416 ();
 sg13g2_decap_8 FILLER_23_2423 ();
 sg13g2_decap_8 FILLER_23_2430 ();
 sg13g2_decap_8 FILLER_23_2437 ();
 sg13g2_decap_8 FILLER_23_2444 ();
 sg13g2_decap_8 FILLER_23_2451 ();
 sg13g2_decap_8 FILLER_23_2458 ();
 sg13g2_decap_8 FILLER_23_2465 ();
 sg13g2_decap_8 FILLER_23_2472 ();
 sg13g2_decap_8 FILLER_23_2479 ();
 sg13g2_decap_8 FILLER_23_2486 ();
 sg13g2_decap_8 FILLER_23_2493 ();
 sg13g2_decap_8 FILLER_23_2500 ();
 sg13g2_decap_8 FILLER_23_2507 ();
 sg13g2_decap_8 FILLER_23_2514 ();
 sg13g2_decap_8 FILLER_23_2521 ();
 sg13g2_decap_8 FILLER_23_2528 ();
 sg13g2_decap_8 FILLER_23_2535 ();
 sg13g2_decap_8 FILLER_23_2542 ();
 sg13g2_decap_8 FILLER_23_2549 ();
 sg13g2_decap_8 FILLER_23_2556 ();
 sg13g2_decap_8 FILLER_23_2563 ();
 sg13g2_decap_8 FILLER_23_2570 ();
 sg13g2_decap_8 FILLER_23_2577 ();
 sg13g2_decap_8 FILLER_23_2584 ();
 sg13g2_decap_8 FILLER_23_2591 ();
 sg13g2_decap_8 FILLER_23_2598 ();
 sg13g2_decap_8 FILLER_23_2605 ();
 sg13g2_decap_8 FILLER_23_2612 ();
 sg13g2_decap_8 FILLER_23_2619 ();
 sg13g2_decap_8 FILLER_23_2626 ();
 sg13g2_decap_8 FILLER_23_2633 ();
 sg13g2_decap_8 FILLER_23_2640 ();
 sg13g2_decap_8 FILLER_23_2647 ();
 sg13g2_decap_8 FILLER_23_2654 ();
 sg13g2_decap_8 FILLER_23_2661 ();
 sg13g2_decap_4 FILLER_23_2668 ();
 sg13g2_fill_2 FILLER_23_2672 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_fill_2 FILLER_24_75 ();
 sg13g2_fill_1 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_251 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_416 ();
 sg13g2_fill_1 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_449 ();
 sg13g2_fill_1 FILLER_24_456 ();
 sg13g2_fill_1 FILLER_24_497 ();
 sg13g2_fill_2 FILLER_24_505 ();
 sg13g2_fill_1 FILLER_24_507 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_fill_1 FILLER_24_515 ();
 sg13g2_decap_4 FILLER_24_520 ();
 sg13g2_fill_2 FILLER_24_524 ();
 sg13g2_fill_2 FILLER_24_532 ();
 sg13g2_fill_1 FILLER_24_534 ();
 sg13g2_fill_2 FILLER_24_544 ();
 sg13g2_fill_2 FILLER_24_551 ();
 sg13g2_fill_1 FILLER_24_553 ();
 sg13g2_fill_1 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_563 ();
 sg13g2_fill_2 FILLER_24_570 ();
 sg13g2_fill_1 FILLER_24_572 ();
 sg13g2_decap_4 FILLER_24_583 ();
 sg13g2_fill_1 FILLER_24_597 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_fill_2 FILLER_24_609 ();
 sg13g2_fill_1 FILLER_24_611 ();
 sg13g2_fill_1 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_640 ();
 sg13g2_decap_8 FILLER_24_647 ();
 sg13g2_decap_8 FILLER_24_654 ();
 sg13g2_decap_8 FILLER_24_661 ();
 sg13g2_fill_1 FILLER_24_693 ();
 sg13g2_fill_2 FILLER_24_699 ();
 sg13g2_fill_1 FILLER_24_701 ();
 sg13g2_fill_1 FILLER_24_708 ();
 sg13g2_decap_4 FILLER_24_776 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_fill_1 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_889 ();
 sg13g2_fill_2 FILLER_24_896 ();
 sg13g2_fill_1 FILLER_24_903 ();
 sg13g2_fill_2 FILLER_24_951 ();
 sg13g2_fill_2 FILLER_24_966 ();
 sg13g2_decap_8 FILLER_24_1014 ();
 sg13g2_decap_8 FILLER_24_1021 ();
 sg13g2_fill_2 FILLER_24_1028 ();
 sg13g2_fill_1 FILLER_24_1058 ();
 sg13g2_fill_2 FILLER_24_1147 ();
 sg13g2_decap_8 FILLER_24_1195 ();
 sg13g2_decap_4 FILLER_24_1202 ();
 sg13g2_fill_2 FILLER_24_1206 ();
 sg13g2_fill_2 FILLER_24_1257 ();
 sg13g2_fill_2 FILLER_24_1321 ();
 sg13g2_fill_1 FILLER_24_1323 ();
 sg13g2_fill_1 FILLER_24_1356 ();
 sg13g2_fill_2 FILLER_24_1361 ();
 sg13g2_fill_1 FILLER_24_1363 ();
 sg13g2_fill_1 FILLER_24_1430 ();
 sg13g2_fill_2 FILLER_24_1463 ();
 sg13g2_decap_4 FILLER_24_1509 ();
 sg13g2_fill_1 FILLER_24_1532 ();
 sg13g2_fill_2 FILLER_24_1546 ();
 sg13g2_fill_1 FILLER_24_1548 ();
 sg13g2_decap_4 FILLER_24_1567 ();
 sg13g2_fill_2 FILLER_24_1571 ();
 sg13g2_fill_2 FILLER_24_1577 ();
 sg13g2_fill_1 FILLER_24_1579 ();
 sg13g2_fill_2 FILLER_24_1598 ();
 sg13g2_fill_2 FILLER_24_1623 ();
 sg13g2_fill_2 FILLER_24_1701 ();
 sg13g2_fill_1 FILLER_24_1779 ();
 sg13g2_fill_2 FILLER_24_1794 ();
 sg13g2_fill_1 FILLER_24_1796 ();
 sg13g2_decap_8 FILLER_24_1828 ();
 sg13g2_fill_2 FILLER_24_1835 ();
 sg13g2_fill_2 FILLER_24_1869 ();
 sg13g2_fill_1 FILLER_24_1871 ();
 sg13g2_fill_2 FILLER_24_1884 ();
 sg13g2_fill_1 FILLER_24_1886 ();
 sg13g2_fill_1 FILLER_24_1908 ();
 sg13g2_decap_4 FILLER_24_1922 ();
 sg13g2_decap_8 FILLER_24_1949 ();
 sg13g2_decap_4 FILLER_24_1956 ();
 sg13g2_decap_8 FILLER_24_1973 ();
 sg13g2_decap_8 FILLER_24_1980 ();
 sg13g2_decap_4 FILLER_24_1987 ();
 sg13g2_fill_2 FILLER_24_2038 ();
 sg13g2_fill_1 FILLER_24_2040 ();
 sg13g2_decap_4 FILLER_24_2074 ();
 sg13g2_fill_2 FILLER_24_2106 ();
 sg13g2_fill_1 FILLER_24_2108 ();
 sg13g2_fill_2 FILLER_24_2118 ();
 sg13g2_fill_1 FILLER_24_2148 ();
 sg13g2_fill_2 FILLER_24_2154 ();
 sg13g2_fill_1 FILLER_24_2161 ();
 sg13g2_fill_1 FILLER_24_2213 ();
 sg13g2_fill_2 FILLER_24_2232 ();
 sg13g2_fill_1 FILLER_24_2234 ();
 sg13g2_decap_8 FILLER_24_2244 ();
 sg13g2_decap_8 FILLER_24_2251 ();
 sg13g2_decap_8 FILLER_24_2258 ();
 sg13g2_decap_8 FILLER_24_2265 ();
 sg13g2_decap_8 FILLER_24_2272 ();
 sg13g2_decap_8 FILLER_24_2279 ();
 sg13g2_decap_8 FILLER_24_2286 ();
 sg13g2_decap_8 FILLER_24_2293 ();
 sg13g2_decap_8 FILLER_24_2300 ();
 sg13g2_decap_8 FILLER_24_2307 ();
 sg13g2_decap_8 FILLER_24_2314 ();
 sg13g2_decap_8 FILLER_24_2321 ();
 sg13g2_decap_8 FILLER_24_2328 ();
 sg13g2_decap_8 FILLER_24_2335 ();
 sg13g2_decap_8 FILLER_24_2342 ();
 sg13g2_decap_8 FILLER_24_2349 ();
 sg13g2_decap_8 FILLER_24_2356 ();
 sg13g2_decap_8 FILLER_24_2363 ();
 sg13g2_decap_8 FILLER_24_2370 ();
 sg13g2_decap_8 FILLER_24_2377 ();
 sg13g2_decap_8 FILLER_24_2384 ();
 sg13g2_decap_8 FILLER_24_2391 ();
 sg13g2_decap_8 FILLER_24_2398 ();
 sg13g2_decap_8 FILLER_24_2405 ();
 sg13g2_decap_8 FILLER_24_2412 ();
 sg13g2_decap_8 FILLER_24_2419 ();
 sg13g2_decap_8 FILLER_24_2426 ();
 sg13g2_decap_8 FILLER_24_2433 ();
 sg13g2_decap_8 FILLER_24_2440 ();
 sg13g2_decap_8 FILLER_24_2447 ();
 sg13g2_decap_8 FILLER_24_2454 ();
 sg13g2_decap_8 FILLER_24_2461 ();
 sg13g2_decap_8 FILLER_24_2468 ();
 sg13g2_decap_8 FILLER_24_2475 ();
 sg13g2_decap_8 FILLER_24_2482 ();
 sg13g2_decap_8 FILLER_24_2489 ();
 sg13g2_decap_8 FILLER_24_2496 ();
 sg13g2_decap_8 FILLER_24_2503 ();
 sg13g2_decap_8 FILLER_24_2510 ();
 sg13g2_decap_8 FILLER_24_2517 ();
 sg13g2_decap_8 FILLER_24_2524 ();
 sg13g2_decap_8 FILLER_24_2531 ();
 sg13g2_decap_8 FILLER_24_2538 ();
 sg13g2_decap_8 FILLER_24_2545 ();
 sg13g2_decap_8 FILLER_24_2552 ();
 sg13g2_decap_8 FILLER_24_2559 ();
 sg13g2_decap_8 FILLER_24_2566 ();
 sg13g2_decap_8 FILLER_24_2573 ();
 sg13g2_decap_8 FILLER_24_2580 ();
 sg13g2_decap_8 FILLER_24_2587 ();
 sg13g2_decap_8 FILLER_24_2594 ();
 sg13g2_decap_8 FILLER_24_2601 ();
 sg13g2_decap_8 FILLER_24_2608 ();
 sg13g2_decap_8 FILLER_24_2615 ();
 sg13g2_decap_8 FILLER_24_2622 ();
 sg13g2_decap_8 FILLER_24_2629 ();
 sg13g2_decap_8 FILLER_24_2636 ();
 sg13g2_decap_8 FILLER_24_2643 ();
 sg13g2_decap_8 FILLER_24_2650 ();
 sg13g2_decap_8 FILLER_24_2657 ();
 sg13g2_decap_8 FILLER_24_2664 ();
 sg13g2_fill_2 FILLER_24_2671 ();
 sg13g2_fill_1 FILLER_24_2673 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_fill_2 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_398 ();
 sg13g2_fill_2 FILLER_25_409 ();
 sg13g2_fill_1 FILLER_25_411 ();
 sg13g2_decap_4 FILLER_25_417 ();
 sg13g2_fill_1 FILLER_25_421 ();
 sg13g2_decap_4 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_435 ();
 sg13g2_decap_4 FILLER_25_442 ();
 sg13g2_decap_8 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_480 ();
 sg13g2_decap_4 FILLER_25_487 ();
 sg13g2_fill_2 FILLER_25_491 ();
 sg13g2_fill_1 FILLER_25_497 ();
 sg13g2_fill_2 FILLER_25_530 ();
 sg13g2_decap_8 FILLER_25_545 ();
 sg13g2_decap_4 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_564 ();
 sg13g2_fill_1 FILLER_25_571 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_decap_8 FILLER_25_589 ();
 sg13g2_decap_8 FILLER_25_596 ();
 sg13g2_decap_8 FILLER_25_603 ();
 sg13g2_fill_2 FILLER_25_610 ();
 sg13g2_decap_4 FILLER_25_617 ();
 sg13g2_decap_8 FILLER_25_655 ();
 sg13g2_decap_8 FILLER_25_662 ();
 sg13g2_fill_1 FILLER_25_669 ();
 sg13g2_fill_1 FILLER_25_675 ();
 sg13g2_decap_4 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_740 ();
 sg13g2_decap_4 FILLER_25_747 ();
 sg13g2_fill_1 FILLER_25_751 ();
 sg13g2_decap_4 FILLER_25_793 ();
 sg13g2_fill_2 FILLER_25_797 ();
 sg13g2_fill_2 FILLER_25_805 ();
 sg13g2_decap_4 FILLER_25_811 ();
 sg13g2_fill_1 FILLER_25_833 ();
 sg13g2_fill_1 FILLER_25_852 ();
 sg13g2_decap_4 FILLER_25_888 ();
 sg13g2_fill_2 FILLER_25_892 ();
 sg13g2_fill_2 FILLER_25_899 ();
 sg13g2_fill_1 FILLER_25_901 ();
 sg13g2_fill_2 FILLER_25_970 ();
 sg13g2_fill_1 FILLER_25_972 ();
 sg13g2_fill_2 FILLER_25_976 ();
 sg13g2_decap_4 FILLER_25_984 ();
 sg13g2_fill_1 FILLER_25_988 ();
 sg13g2_decap_8 FILLER_25_1024 ();
 sg13g2_decap_8 FILLER_25_1031 ();
 sg13g2_fill_2 FILLER_25_1038 ();
 sg13g2_fill_1 FILLER_25_1040 ();
 sg13g2_fill_2 FILLER_25_1062 ();
 sg13g2_fill_1 FILLER_25_1064 ();
 sg13g2_decap_8 FILLER_25_1079 ();
 sg13g2_decap_8 FILLER_25_1086 ();
 sg13g2_decap_8 FILLER_25_1093 ();
 sg13g2_fill_2 FILLER_25_1100 ();
 sg13g2_fill_1 FILLER_25_1161 ();
 sg13g2_fill_2 FILLER_25_1175 ();
 sg13g2_fill_2 FILLER_25_1190 ();
 sg13g2_decap_4 FILLER_25_1201 ();
 sg13g2_fill_1 FILLER_25_1205 ();
 sg13g2_fill_1 FILLER_25_1239 ();
 sg13g2_fill_2 FILLER_25_1291 ();
 sg13g2_fill_1 FILLER_25_1293 ();
 sg13g2_decap_4 FILLER_25_1337 ();
 sg13g2_fill_2 FILLER_25_1381 ();
 sg13g2_fill_1 FILLER_25_1383 ();
 sg13g2_fill_2 FILLER_25_1417 ();
 sg13g2_fill_1 FILLER_25_1419 ();
 sg13g2_fill_1 FILLER_25_1457 ();
 sg13g2_fill_2 FILLER_25_1510 ();
 sg13g2_fill_2 FILLER_25_1532 ();
 sg13g2_fill_2 FILLER_25_1567 ();
 sg13g2_fill_2 FILLER_25_1616 ();
 sg13g2_fill_2 FILLER_25_1686 ();
 sg13g2_decap_8 FILLER_25_1793 ();
 sg13g2_decap_8 FILLER_25_1800 ();
 sg13g2_fill_1 FILLER_25_1807 ();
 sg13g2_fill_2 FILLER_25_1877 ();
 sg13g2_fill_1 FILLER_25_1879 ();
 sg13g2_fill_1 FILLER_25_1892 ();
 sg13g2_fill_1 FILLER_25_1903 ();
 sg13g2_fill_1 FILLER_25_1923 ();
 sg13g2_fill_1 FILLER_25_1956 ();
 sg13g2_fill_2 FILLER_25_1984 ();
 sg13g2_fill_2 FILLER_25_2039 ();
 sg13g2_decap_4 FILLER_25_2078 ();
 sg13g2_fill_1 FILLER_25_2082 ();
 sg13g2_fill_1 FILLER_25_2154 ();
 sg13g2_fill_2 FILLER_25_2178 ();
 sg13g2_fill_1 FILLER_25_2195 ();
 sg13g2_fill_2 FILLER_25_2219 ();
 sg13g2_decap_8 FILLER_25_2249 ();
 sg13g2_decap_8 FILLER_25_2256 ();
 sg13g2_decap_8 FILLER_25_2263 ();
 sg13g2_decap_8 FILLER_25_2270 ();
 sg13g2_decap_8 FILLER_25_2277 ();
 sg13g2_decap_8 FILLER_25_2284 ();
 sg13g2_decap_8 FILLER_25_2291 ();
 sg13g2_decap_8 FILLER_25_2298 ();
 sg13g2_decap_8 FILLER_25_2305 ();
 sg13g2_decap_8 FILLER_25_2312 ();
 sg13g2_decap_8 FILLER_25_2319 ();
 sg13g2_decap_8 FILLER_25_2326 ();
 sg13g2_decap_8 FILLER_25_2333 ();
 sg13g2_decap_8 FILLER_25_2340 ();
 sg13g2_decap_8 FILLER_25_2347 ();
 sg13g2_decap_8 FILLER_25_2354 ();
 sg13g2_decap_8 FILLER_25_2361 ();
 sg13g2_decap_8 FILLER_25_2368 ();
 sg13g2_decap_8 FILLER_25_2375 ();
 sg13g2_decap_8 FILLER_25_2382 ();
 sg13g2_decap_8 FILLER_25_2389 ();
 sg13g2_decap_8 FILLER_25_2396 ();
 sg13g2_decap_8 FILLER_25_2403 ();
 sg13g2_decap_8 FILLER_25_2410 ();
 sg13g2_decap_8 FILLER_25_2417 ();
 sg13g2_decap_8 FILLER_25_2424 ();
 sg13g2_decap_8 FILLER_25_2431 ();
 sg13g2_decap_8 FILLER_25_2438 ();
 sg13g2_decap_8 FILLER_25_2445 ();
 sg13g2_decap_8 FILLER_25_2452 ();
 sg13g2_decap_8 FILLER_25_2459 ();
 sg13g2_decap_8 FILLER_25_2466 ();
 sg13g2_decap_8 FILLER_25_2473 ();
 sg13g2_decap_8 FILLER_25_2480 ();
 sg13g2_decap_8 FILLER_25_2487 ();
 sg13g2_decap_8 FILLER_25_2494 ();
 sg13g2_decap_8 FILLER_25_2501 ();
 sg13g2_decap_8 FILLER_25_2508 ();
 sg13g2_decap_8 FILLER_25_2515 ();
 sg13g2_decap_8 FILLER_25_2522 ();
 sg13g2_decap_8 FILLER_25_2529 ();
 sg13g2_decap_8 FILLER_25_2536 ();
 sg13g2_decap_8 FILLER_25_2543 ();
 sg13g2_decap_8 FILLER_25_2550 ();
 sg13g2_decap_8 FILLER_25_2557 ();
 sg13g2_decap_8 FILLER_25_2564 ();
 sg13g2_decap_8 FILLER_25_2571 ();
 sg13g2_decap_8 FILLER_25_2578 ();
 sg13g2_decap_8 FILLER_25_2585 ();
 sg13g2_decap_8 FILLER_25_2592 ();
 sg13g2_decap_8 FILLER_25_2599 ();
 sg13g2_decap_8 FILLER_25_2606 ();
 sg13g2_decap_8 FILLER_25_2613 ();
 sg13g2_decap_8 FILLER_25_2620 ();
 sg13g2_decap_8 FILLER_25_2627 ();
 sg13g2_decap_8 FILLER_25_2634 ();
 sg13g2_decap_8 FILLER_25_2641 ();
 sg13g2_decap_8 FILLER_25_2648 ();
 sg13g2_decap_8 FILLER_25_2655 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_decap_4 FILLER_25_2669 ();
 sg13g2_fill_1 FILLER_25_2673 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_38 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_2 FILLER_26_421 ();
 sg13g2_fill_1 FILLER_26_423 ();
 sg13g2_decap_8 FILLER_26_445 ();
 sg13g2_fill_2 FILLER_26_452 ();
 sg13g2_decap_8 FILLER_26_458 ();
 sg13g2_decap_8 FILLER_26_465 ();
 sg13g2_fill_1 FILLER_26_472 ();
 sg13g2_decap_4 FILLER_26_479 ();
 sg13g2_fill_1 FILLER_26_521 ();
 sg13g2_fill_2 FILLER_26_558 ();
 sg13g2_decap_8 FILLER_26_565 ();
 sg13g2_decap_8 FILLER_26_572 ();
 sg13g2_fill_1 FILLER_26_579 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_633 ();
 sg13g2_decap_4 FILLER_26_640 ();
 sg13g2_fill_2 FILLER_26_644 ();
 sg13g2_fill_2 FILLER_26_664 ();
 sg13g2_fill_1 FILLER_26_666 ();
 sg13g2_decap_4 FILLER_26_671 ();
 sg13g2_fill_2 FILLER_26_675 ();
 sg13g2_fill_2 FILLER_26_699 ();
 sg13g2_decap_8 FILLER_26_744 ();
 sg13g2_fill_1 FILLER_26_756 ();
 sg13g2_decap_4 FILLER_26_763 ();
 sg13g2_fill_1 FILLER_26_767 ();
 sg13g2_fill_2 FILLER_26_774 ();
 sg13g2_decap_8 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_fill_1 FILLER_26_822 ();
 sg13g2_fill_1 FILLER_26_836 ();
 sg13g2_fill_1 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_881 ();
 sg13g2_fill_1 FILLER_26_888 ();
 sg13g2_fill_2 FILLER_26_924 ();
 sg13g2_fill_1 FILLER_26_961 ();
 sg13g2_fill_2 FILLER_26_975 ();
 sg13g2_fill_1 FILLER_26_977 ();
 sg13g2_fill_2 FILLER_26_987 ();
 sg13g2_fill_2 FILLER_26_1006 ();
 sg13g2_decap_8 FILLER_26_1032 ();
 sg13g2_fill_2 FILLER_26_1039 ();
 sg13g2_fill_1 FILLER_26_1072 ();
 sg13g2_decap_8 FILLER_26_1079 ();
 sg13g2_decap_8 FILLER_26_1086 ();
 sg13g2_decap_4 FILLER_26_1093 ();
 sg13g2_fill_2 FILLER_26_1097 ();
 sg13g2_fill_1 FILLER_26_1105 ();
 sg13g2_fill_2 FILLER_26_1152 ();
 sg13g2_fill_1 FILLER_26_1154 ();
 sg13g2_fill_1 FILLER_26_1209 ();
 sg13g2_fill_1 FILLER_26_1249 ();
 sg13g2_fill_2 FILLER_26_1269 ();
 sg13g2_fill_1 FILLER_26_1302 ();
 sg13g2_decap_8 FILLER_26_1335 ();
 sg13g2_decap_8 FILLER_26_1342 ();
 sg13g2_fill_2 FILLER_26_1349 ();
 sg13g2_decap_8 FILLER_26_1364 ();
 sg13g2_decap_4 FILLER_26_1463 ();
 sg13g2_fill_1 FILLER_26_1504 ();
 sg13g2_fill_1 FILLER_26_1523 ();
 sg13g2_decap_8 FILLER_26_1529 ();
 sg13g2_decap_4 FILLER_26_1536 ();
 sg13g2_fill_1 FILLER_26_1546 ();
 sg13g2_fill_2 FILLER_26_1594 ();
 sg13g2_fill_2 FILLER_26_1606 ();
 sg13g2_fill_1 FILLER_26_1608 ();
 sg13g2_fill_2 FILLER_26_1614 ();
 sg13g2_fill_2 FILLER_26_1630 ();
 sg13g2_fill_2 FILLER_26_1654 ();
 sg13g2_fill_1 FILLER_26_1656 ();
 sg13g2_decap_4 FILLER_26_1705 ();
 sg13g2_fill_2 FILLER_26_1714 ();
 sg13g2_fill_2 FILLER_26_1766 ();
 sg13g2_fill_1 FILLER_26_1768 ();
 sg13g2_fill_2 FILLER_26_1778 ();
 sg13g2_decap_8 FILLER_26_1794 ();
 sg13g2_decap_8 FILLER_26_1869 ();
 sg13g2_decap_4 FILLER_26_1876 ();
 sg13g2_fill_2 FILLER_26_1880 ();
 sg13g2_decap_8 FILLER_26_1918 ();
 sg13g2_fill_2 FILLER_26_1925 ();
 sg13g2_fill_1 FILLER_26_1927 ();
 sg13g2_fill_1 FILLER_26_1959 ();
 sg13g2_fill_1 FILLER_26_1969 ();
 sg13g2_fill_1 FILLER_26_1987 ();
 sg13g2_decap_8 FILLER_26_2078 ();
 sg13g2_decap_8 FILLER_26_2085 ();
 sg13g2_fill_1 FILLER_26_2105 ();
 sg13g2_fill_1 FILLER_26_2111 ();
 sg13g2_fill_2 FILLER_26_2121 ();
 sg13g2_decap_4 FILLER_26_2158 ();
 sg13g2_fill_1 FILLER_26_2162 ();
 sg13g2_fill_1 FILLER_26_2169 ();
 sg13g2_decap_8 FILLER_26_2237 ();
 sg13g2_decap_8 FILLER_26_2244 ();
 sg13g2_decap_8 FILLER_26_2251 ();
 sg13g2_decap_8 FILLER_26_2258 ();
 sg13g2_decap_8 FILLER_26_2265 ();
 sg13g2_decap_8 FILLER_26_2272 ();
 sg13g2_decap_8 FILLER_26_2279 ();
 sg13g2_decap_8 FILLER_26_2286 ();
 sg13g2_decap_8 FILLER_26_2293 ();
 sg13g2_decap_8 FILLER_26_2300 ();
 sg13g2_decap_8 FILLER_26_2307 ();
 sg13g2_decap_8 FILLER_26_2314 ();
 sg13g2_decap_8 FILLER_26_2321 ();
 sg13g2_decap_8 FILLER_26_2328 ();
 sg13g2_decap_8 FILLER_26_2335 ();
 sg13g2_decap_8 FILLER_26_2342 ();
 sg13g2_decap_8 FILLER_26_2349 ();
 sg13g2_decap_8 FILLER_26_2356 ();
 sg13g2_decap_8 FILLER_26_2363 ();
 sg13g2_decap_8 FILLER_26_2370 ();
 sg13g2_decap_8 FILLER_26_2377 ();
 sg13g2_decap_8 FILLER_26_2384 ();
 sg13g2_decap_8 FILLER_26_2391 ();
 sg13g2_decap_8 FILLER_26_2398 ();
 sg13g2_decap_8 FILLER_26_2405 ();
 sg13g2_decap_8 FILLER_26_2412 ();
 sg13g2_decap_8 FILLER_26_2419 ();
 sg13g2_decap_8 FILLER_26_2426 ();
 sg13g2_decap_8 FILLER_26_2433 ();
 sg13g2_decap_8 FILLER_26_2440 ();
 sg13g2_decap_8 FILLER_26_2447 ();
 sg13g2_decap_8 FILLER_26_2454 ();
 sg13g2_decap_8 FILLER_26_2461 ();
 sg13g2_decap_8 FILLER_26_2468 ();
 sg13g2_decap_8 FILLER_26_2475 ();
 sg13g2_decap_8 FILLER_26_2482 ();
 sg13g2_decap_8 FILLER_26_2489 ();
 sg13g2_decap_8 FILLER_26_2496 ();
 sg13g2_decap_8 FILLER_26_2503 ();
 sg13g2_decap_8 FILLER_26_2510 ();
 sg13g2_decap_8 FILLER_26_2517 ();
 sg13g2_decap_8 FILLER_26_2524 ();
 sg13g2_decap_8 FILLER_26_2531 ();
 sg13g2_decap_8 FILLER_26_2538 ();
 sg13g2_decap_8 FILLER_26_2545 ();
 sg13g2_decap_8 FILLER_26_2552 ();
 sg13g2_decap_8 FILLER_26_2559 ();
 sg13g2_decap_8 FILLER_26_2566 ();
 sg13g2_decap_8 FILLER_26_2573 ();
 sg13g2_decap_8 FILLER_26_2580 ();
 sg13g2_decap_8 FILLER_26_2587 ();
 sg13g2_decap_8 FILLER_26_2594 ();
 sg13g2_decap_8 FILLER_26_2601 ();
 sg13g2_decap_8 FILLER_26_2608 ();
 sg13g2_decap_8 FILLER_26_2615 ();
 sg13g2_decap_8 FILLER_26_2622 ();
 sg13g2_decap_8 FILLER_26_2629 ();
 sg13g2_decap_8 FILLER_26_2636 ();
 sg13g2_decap_8 FILLER_26_2643 ();
 sg13g2_decap_8 FILLER_26_2650 ();
 sg13g2_decap_8 FILLER_26_2657 ();
 sg13g2_decap_8 FILLER_26_2664 ();
 sg13g2_fill_2 FILLER_26_2671 ();
 sg13g2_fill_1 FILLER_26_2673 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_40 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_fill_1 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_468 ();
 sg13g2_fill_2 FILLER_27_545 ();
 sg13g2_fill_1 FILLER_27_547 ();
 sg13g2_decap_8 FILLER_27_562 ();
 sg13g2_decap_8 FILLER_27_569 ();
 sg13g2_decap_4 FILLER_27_595 ();
 sg13g2_fill_1 FILLER_27_599 ();
 sg13g2_decap_4 FILLER_27_636 ();
 sg13g2_fill_1 FILLER_27_640 ();
 sg13g2_decap_4 FILLER_27_645 ();
 sg13g2_fill_1 FILLER_27_649 ();
 sg13g2_decap_4 FILLER_27_661 ();
 sg13g2_fill_2 FILLER_27_696 ();
 sg13g2_fill_1 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_fill_2 FILLER_27_772 ();
 sg13g2_decap_4 FILLER_27_790 ();
 sg13g2_fill_1 FILLER_27_829 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_4 FILLER_27_977 ();
 sg13g2_fill_2 FILLER_27_981 ();
 sg13g2_fill_2 FILLER_27_996 ();
 sg13g2_fill_1 FILLER_27_998 ();
 sg13g2_fill_2 FILLER_27_1018 ();
 sg13g2_decap_4 FILLER_27_1025 ();
 sg13g2_fill_2 FILLER_27_1056 ();
 sg13g2_fill_1 FILLER_27_1058 ();
 sg13g2_fill_1 FILLER_27_1064 ();
 sg13g2_decap_8 FILLER_27_1078 ();
 sg13g2_fill_2 FILLER_27_1085 ();
 sg13g2_fill_1 FILLER_27_1087 ();
 sg13g2_fill_2 FILLER_27_1094 ();
 sg13g2_fill_2 FILLER_27_1141 ();
 sg13g2_fill_1 FILLER_27_1143 ();
 sg13g2_fill_2 FILLER_27_1161 ();
 sg13g2_fill_2 FILLER_27_1183 ();
 sg13g2_fill_2 FILLER_27_1253 ();
 sg13g2_fill_2 FILLER_27_1333 ();
 sg13g2_decap_4 FILLER_27_1344 ();
 sg13g2_fill_1 FILLER_27_1348 ();
 sg13g2_fill_1 FILLER_27_1368 ();
 sg13g2_fill_1 FILLER_27_1382 ();
 sg13g2_fill_2 FILLER_27_1396 ();
 sg13g2_fill_2 FILLER_27_1410 ();
 sg13g2_fill_1 FILLER_27_1412 ();
 sg13g2_fill_2 FILLER_27_1417 ();
 sg13g2_fill_1 FILLER_27_1419 ();
 sg13g2_fill_1 FILLER_27_1452 ();
 sg13g2_decap_8 FILLER_27_1458 ();
 sg13g2_fill_2 FILLER_27_1465 ();
 sg13g2_decap_8 FILLER_27_1472 ();
 sg13g2_decap_8 FILLER_27_1479 ();
 sg13g2_fill_2 FILLER_27_1486 ();
 sg13g2_fill_1 FILLER_27_1501 ();
 sg13g2_fill_1 FILLER_27_1579 ();
 sg13g2_fill_2 FILLER_27_1586 ();
 sg13g2_fill_1 FILLER_27_1601 ();
 sg13g2_fill_1 FILLER_27_1641 ();
 sg13g2_fill_1 FILLER_27_1708 ();
 sg13g2_fill_2 FILLER_27_1727 ();
 sg13g2_fill_1 FILLER_27_1729 ();
 sg13g2_fill_2 FILLER_27_1743 ();
 sg13g2_fill_1 FILLER_27_1763 ();
 sg13g2_fill_1 FILLER_27_1780 ();
 sg13g2_fill_1 FILLER_27_1792 ();
 sg13g2_fill_1 FILLER_27_1805 ();
 sg13g2_fill_1 FILLER_27_1816 ();
 sg13g2_decap_4 FILLER_27_1837 ();
 sg13g2_decap_8 FILLER_27_1859 ();
 sg13g2_decap_4 FILLER_27_1866 ();
 sg13g2_fill_1 FILLER_27_1879 ();
 sg13g2_decap_8 FILLER_27_1908 ();
 sg13g2_decap_8 FILLER_27_1915 ();
 sg13g2_decap_4 FILLER_27_1930 ();
 sg13g2_fill_2 FILLER_27_1971 ();
 sg13g2_fill_1 FILLER_27_1973 ();
 sg13g2_decap_8 FILLER_27_1979 ();
 sg13g2_decap_8 FILLER_27_1986 ();
 sg13g2_fill_2 FILLER_27_1993 ();
 sg13g2_fill_1 FILLER_27_1995 ();
 sg13g2_decap_8 FILLER_27_2018 ();
 sg13g2_fill_2 FILLER_27_2025 ();
 sg13g2_fill_1 FILLER_27_2037 ();
 sg13g2_fill_1 FILLER_27_2043 ();
 sg13g2_fill_2 FILLER_27_2100 ();
 sg13g2_fill_1 FILLER_27_2102 ();
 sg13g2_decap_8 FILLER_27_2164 ();
 sg13g2_decap_8 FILLER_27_2237 ();
 sg13g2_decap_8 FILLER_27_2244 ();
 sg13g2_decap_8 FILLER_27_2251 ();
 sg13g2_decap_8 FILLER_27_2258 ();
 sg13g2_decap_8 FILLER_27_2265 ();
 sg13g2_decap_8 FILLER_27_2272 ();
 sg13g2_decap_8 FILLER_27_2279 ();
 sg13g2_decap_8 FILLER_27_2286 ();
 sg13g2_decap_8 FILLER_27_2293 ();
 sg13g2_decap_8 FILLER_27_2300 ();
 sg13g2_decap_8 FILLER_27_2307 ();
 sg13g2_decap_8 FILLER_27_2314 ();
 sg13g2_decap_8 FILLER_27_2321 ();
 sg13g2_decap_8 FILLER_27_2328 ();
 sg13g2_decap_8 FILLER_27_2335 ();
 sg13g2_decap_8 FILLER_27_2342 ();
 sg13g2_decap_8 FILLER_27_2349 ();
 sg13g2_decap_8 FILLER_27_2356 ();
 sg13g2_decap_8 FILLER_27_2363 ();
 sg13g2_decap_8 FILLER_27_2370 ();
 sg13g2_decap_8 FILLER_27_2377 ();
 sg13g2_decap_8 FILLER_27_2384 ();
 sg13g2_decap_8 FILLER_27_2391 ();
 sg13g2_decap_8 FILLER_27_2398 ();
 sg13g2_decap_8 FILLER_27_2405 ();
 sg13g2_decap_8 FILLER_27_2412 ();
 sg13g2_decap_8 FILLER_27_2419 ();
 sg13g2_decap_8 FILLER_27_2426 ();
 sg13g2_decap_8 FILLER_27_2433 ();
 sg13g2_decap_8 FILLER_27_2440 ();
 sg13g2_decap_8 FILLER_27_2447 ();
 sg13g2_decap_8 FILLER_27_2454 ();
 sg13g2_decap_8 FILLER_27_2461 ();
 sg13g2_decap_8 FILLER_27_2468 ();
 sg13g2_decap_8 FILLER_27_2475 ();
 sg13g2_decap_8 FILLER_27_2482 ();
 sg13g2_decap_8 FILLER_27_2489 ();
 sg13g2_decap_8 FILLER_27_2496 ();
 sg13g2_decap_8 FILLER_27_2503 ();
 sg13g2_decap_8 FILLER_27_2510 ();
 sg13g2_decap_8 FILLER_27_2517 ();
 sg13g2_decap_8 FILLER_27_2524 ();
 sg13g2_decap_8 FILLER_27_2531 ();
 sg13g2_decap_8 FILLER_27_2538 ();
 sg13g2_decap_8 FILLER_27_2545 ();
 sg13g2_decap_8 FILLER_27_2552 ();
 sg13g2_decap_8 FILLER_27_2559 ();
 sg13g2_decap_8 FILLER_27_2566 ();
 sg13g2_decap_8 FILLER_27_2573 ();
 sg13g2_decap_8 FILLER_27_2580 ();
 sg13g2_decap_8 FILLER_27_2587 ();
 sg13g2_decap_8 FILLER_27_2594 ();
 sg13g2_decap_8 FILLER_27_2601 ();
 sg13g2_decap_8 FILLER_27_2608 ();
 sg13g2_decap_8 FILLER_27_2615 ();
 sg13g2_decap_8 FILLER_27_2622 ();
 sg13g2_decap_8 FILLER_27_2629 ();
 sg13g2_decap_8 FILLER_27_2636 ();
 sg13g2_decap_8 FILLER_27_2643 ();
 sg13g2_decap_8 FILLER_27_2650 ();
 sg13g2_decap_8 FILLER_27_2657 ();
 sg13g2_decap_8 FILLER_27_2664 ();
 sg13g2_fill_2 FILLER_27_2671 ();
 sg13g2_fill_1 FILLER_27_2673 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_fill_2 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_457 ();
 sg13g2_fill_2 FILLER_28_508 ();
 sg13g2_fill_2 FILLER_28_544 ();
 sg13g2_decap_8 FILLER_28_563 ();
 sg13g2_decap_8 FILLER_28_570 ();
 sg13g2_decap_8 FILLER_28_577 ();
 sg13g2_fill_2 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_decap_4 FILLER_28_608 ();
 sg13g2_fill_2 FILLER_28_612 ();
 sg13g2_fill_2 FILLER_28_628 ();
 sg13g2_decap_8 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_645 ();
 sg13g2_fill_1 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_744 ();
 sg13g2_fill_1 FILLER_28_751 ();
 sg13g2_decap_8 FILLER_28_800 ();
 sg13g2_fill_1 FILLER_28_864 ();
 sg13g2_decap_8 FILLER_28_880 ();
 sg13g2_decap_8 FILLER_28_887 ();
 sg13g2_fill_1 FILLER_28_894 ();
 sg13g2_fill_2 FILLER_28_945 ();
 sg13g2_fill_2 FILLER_28_1037 ();
 sg13g2_fill_2 FILLER_28_1053 ();
 sg13g2_decap_8 FILLER_28_1077 ();
 sg13g2_decap_8 FILLER_28_1084 ();
 sg13g2_fill_1 FILLER_28_1091 ();
 sg13g2_fill_2 FILLER_28_1215 ();
 sg13g2_fill_1 FILLER_28_1217 ();
 sg13g2_fill_1 FILLER_28_1249 ();
 sg13g2_fill_2 FILLER_28_1263 ();
 sg13g2_fill_2 FILLER_28_1316 ();
 sg13g2_fill_2 FILLER_28_1323 ();
 sg13g2_decap_8 FILLER_28_1348 ();
 sg13g2_decap_8 FILLER_28_1355 ();
 sg13g2_decap_4 FILLER_28_1362 ();
 sg13g2_fill_2 FILLER_28_1415 ();
 sg13g2_fill_1 FILLER_28_1417 ();
 sg13g2_fill_2 FILLER_28_1436 ();
 sg13g2_decap_4 FILLER_28_1474 ();
 sg13g2_fill_1 FILLER_28_1478 ();
 sg13g2_decap_8 FILLER_28_1497 ();
 sg13g2_fill_1 FILLER_28_1504 ();
 sg13g2_fill_2 FILLER_28_1531 ();
 sg13g2_fill_2 FILLER_28_1606 ();
 sg13g2_fill_2 FILLER_28_1650 ();
 sg13g2_fill_1 FILLER_28_1667 ();
 sg13g2_fill_1 FILLER_28_1709 ();
 sg13g2_fill_2 FILLER_28_1731 ();
 sg13g2_fill_2 FILLER_28_1767 ();
 sg13g2_fill_2 FILLER_28_1796 ();
 sg13g2_fill_1 FILLER_28_1798 ();
 sg13g2_fill_2 FILLER_28_1815 ();
 sg13g2_fill_1 FILLER_28_1817 ();
 sg13g2_decap_8 FILLER_28_1845 ();
 sg13g2_fill_2 FILLER_28_1852 ();
 sg13g2_fill_1 FILLER_28_1854 ();
 sg13g2_fill_2 FILLER_28_1868 ();
 sg13g2_fill_1 FILLER_28_1870 ();
 sg13g2_fill_2 FILLER_28_1884 ();
 sg13g2_fill_1 FILLER_28_1886 ();
 sg13g2_fill_2 FILLER_28_1902 ();
 sg13g2_decap_8 FILLER_28_1913 ();
 sg13g2_fill_1 FILLER_28_1920 ();
 sg13g2_fill_2 FILLER_28_1942 ();
 sg13g2_fill_2 FILLER_28_1962 ();
 sg13g2_fill_1 FILLER_28_1964 ();
 sg13g2_fill_1 FILLER_28_1975 ();
 sg13g2_decap_8 FILLER_28_2003 ();
 sg13g2_decap_4 FILLER_28_2010 ();
 sg13g2_fill_2 FILLER_28_2014 ();
 sg13g2_fill_1 FILLER_28_2042 ();
 sg13g2_fill_2 FILLER_28_2071 ();
 sg13g2_fill_1 FILLER_28_2073 ();
 sg13g2_fill_2 FILLER_28_2111 ();
 sg13g2_fill_1 FILLER_28_2113 ();
 sg13g2_decap_8 FILLER_28_2155 ();
 sg13g2_decap_8 FILLER_28_2162 ();
 sg13g2_fill_1 FILLER_28_2169 ();
 sg13g2_fill_2 FILLER_28_2184 ();
 sg13g2_fill_1 FILLER_28_2219 ();
 sg13g2_decap_8 FILLER_28_2253 ();
 sg13g2_decap_8 FILLER_28_2260 ();
 sg13g2_decap_8 FILLER_28_2267 ();
 sg13g2_decap_8 FILLER_28_2274 ();
 sg13g2_decap_8 FILLER_28_2281 ();
 sg13g2_decap_8 FILLER_28_2288 ();
 sg13g2_decap_8 FILLER_28_2295 ();
 sg13g2_decap_8 FILLER_28_2302 ();
 sg13g2_decap_8 FILLER_28_2309 ();
 sg13g2_decap_8 FILLER_28_2316 ();
 sg13g2_decap_8 FILLER_28_2323 ();
 sg13g2_decap_8 FILLER_28_2330 ();
 sg13g2_decap_8 FILLER_28_2337 ();
 sg13g2_decap_8 FILLER_28_2344 ();
 sg13g2_decap_8 FILLER_28_2351 ();
 sg13g2_decap_8 FILLER_28_2358 ();
 sg13g2_decap_8 FILLER_28_2365 ();
 sg13g2_decap_8 FILLER_28_2372 ();
 sg13g2_decap_8 FILLER_28_2379 ();
 sg13g2_decap_8 FILLER_28_2386 ();
 sg13g2_decap_8 FILLER_28_2393 ();
 sg13g2_decap_8 FILLER_28_2400 ();
 sg13g2_decap_8 FILLER_28_2407 ();
 sg13g2_decap_8 FILLER_28_2414 ();
 sg13g2_decap_8 FILLER_28_2421 ();
 sg13g2_decap_8 FILLER_28_2428 ();
 sg13g2_decap_8 FILLER_28_2435 ();
 sg13g2_decap_8 FILLER_28_2442 ();
 sg13g2_decap_8 FILLER_28_2449 ();
 sg13g2_decap_8 FILLER_28_2456 ();
 sg13g2_decap_8 FILLER_28_2463 ();
 sg13g2_decap_8 FILLER_28_2470 ();
 sg13g2_decap_8 FILLER_28_2477 ();
 sg13g2_decap_8 FILLER_28_2484 ();
 sg13g2_decap_8 FILLER_28_2491 ();
 sg13g2_decap_8 FILLER_28_2498 ();
 sg13g2_decap_8 FILLER_28_2505 ();
 sg13g2_decap_8 FILLER_28_2512 ();
 sg13g2_decap_8 FILLER_28_2519 ();
 sg13g2_decap_8 FILLER_28_2526 ();
 sg13g2_decap_8 FILLER_28_2533 ();
 sg13g2_decap_8 FILLER_28_2540 ();
 sg13g2_decap_8 FILLER_28_2547 ();
 sg13g2_decap_8 FILLER_28_2554 ();
 sg13g2_decap_8 FILLER_28_2561 ();
 sg13g2_decap_8 FILLER_28_2568 ();
 sg13g2_decap_8 FILLER_28_2575 ();
 sg13g2_decap_8 FILLER_28_2582 ();
 sg13g2_decap_8 FILLER_28_2589 ();
 sg13g2_decap_8 FILLER_28_2596 ();
 sg13g2_decap_8 FILLER_28_2603 ();
 sg13g2_decap_8 FILLER_28_2610 ();
 sg13g2_decap_8 FILLER_28_2617 ();
 sg13g2_decap_8 FILLER_28_2624 ();
 sg13g2_decap_8 FILLER_28_2631 ();
 sg13g2_decap_8 FILLER_28_2638 ();
 sg13g2_decap_8 FILLER_28_2645 ();
 sg13g2_decap_8 FILLER_28_2652 ();
 sg13g2_decap_8 FILLER_28_2659 ();
 sg13g2_decap_8 FILLER_28_2666 ();
 sg13g2_fill_1 FILLER_28_2673 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_fill_1 FILLER_29_41 ();
 sg13g2_decap_4 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_fill_1 FILLER_29_404 ();
 sg13g2_fill_2 FILLER_29_441 ();
 sg13g2_fill_1 FILLER_29_494 ();
 sg13g2_fill_2 FILLER_29_521 ();
 sg13g2_fill_2 FILLER_29_556 ();
 sg13g2_fill_1 FILLER_29_558 ();
 sg13g2_decap_8 FILLER_29_563 ();
 sg13g2_decap_8 FILLER_29_570 ();
 sg13g2_decap_4 FILLER_29_591 ();
 sg13g2_fill_2 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_4 FILLER_29_623 ();
 sg13g2_fill_2 FILLER_29_627 ();
 sg13g2_fill_2 FILLER_29_634 ();
 sg13g2_fill_2 FILLER_29_647 ();
 sg13g2_fill_1 FILLER_29_649 ();
 sg13g2_fill_1 FILLER_29_660 ();
 sg13g2_fill_1 FILLER_29_674 ();
 sg13g2_fill_2 FILLER_29_680 ();
 sg13g2_fill_1 FILLER_29_682 ();
 sg13g2_fill_1 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_698 ();
 sg13g2_decap_8 FILLER_29_705 ();
 sg13g2_fill_1 FILLER_29_712 ();
 sg13g2_decap_4 FILLER_29_736 ();
 sg13g2_fill_1 FILLER_29_740 ();
 sg13g2_fill_1 FILLER_29_863 ();
 sg13g2_decap_4 FILLER_29_871 ();
 sg13g2_fill_2 FILLER_29_889 ();
 sg13g2_fill_2 FILLER_29_917 ();
 sg13g2_fill_2 FILLER_29_961 ();
 sg13g2_fill_1 FILLER_29_963 ();
 sg13g2_fill_1 FILLER_29_996 ();
 sg13g2_fill_1 FILLER_29_1006 ();
 sg13g2_decap_4 FILLER_29_1033 ();
 sg13g2_fill_1 FILLER_29_1041 ();
 sg13g2_fill_1 FILLER_29_1050 ();
 sg13g2_decap_4 FILLER_29_1082 ();
 sg13g2_fill_2 FILLER_29_1086 ();
 sg13g2_fill_2 FILLER_29_1113 ();
 sg13g2_fill_1 FILLER_29_1115 ();
 sg13g2_decap_4 FILLER_29_1188 ();
 sg13g2_decap_4 FILLER_29_1201 ();
 sg13g2_fill_1 FILLER_29_1205 ();
 sg13g2_fill_1 FILLER_29_1246 ();
 sg13g2_fill_2 FILLER_29_1308 ();
 sg13g2_fill_1 FILLER_29_1328 ();
 sg13g2_decap_8 FILLER_29_1355 ();
 sg13g2_fill_2 FILLER_29_1362 ();
 sg13g2_fill_1 FILLER_29_1364 ();
 sg13g2_fill_2 FILLER_29_1417 ();
 sg13g2_fill_2 FILLER_29_1432 ();
 sg13g2_fill_1 FILLER_29_1434 ();
 sg13g2_fill_2 FILLER_29_1508 ();
 sg13g2_fill_2 FILLER_29_1533 ();
 sg13g2_fill_1 FILLER_29_1555 ();
 sg13g2_fill_1 FILLER_29_1607 ();
 sg13g2_fill_1 FILLER_29_1626 ();
 sg13g2_fill_2 FILLER_29_1713 ();
 sg13g2_fill_1 FILLER_29_1743 ();
 sg13g2_fill_1 FILLER_29_1785 ();
 sg13g2_fill_2 FILLER_29_1829 ();
 sg13g2_fill_1 FILLER_29_1831 ();
 sg13g2_fill_2 FILLER_29_1860 ();
 sg13g2_fill_2 FILLER_29_1899 ();
 sg13g2_decap_4 FILLER_29_1905 ();
 sg13g2_fill_2 FILLER_29_1909 ();
 sg13g2_fill_2 FILLER_29_1951 ();
 sg13g2_decap_8 FILLER_29_2007 ();
 sg13g2_decap_4 FILLER_29_2014 ();
 sg13g2_fill_2 FILLER_29_2065 ();
 sg13g2_decap_8 FILLER_29_2108 ();
 sg13g2_decap_8 FILLER_29_2115 ();
 sg13g2_fill_1 FILLER_29_2122 ();
 sg13g2_decap_4 FILLER_29_2154 ();
 sg13g2_fill_2 FILLER_29_2158 ();
 sg13g2_fill_1 FILLER_29_2173 ();
 sg13g2_fill_1 FILLER_29_2187 ();
 sg13g2_decap_8 FILLER_29_2247 ();
 sg13g2_decap_8 FILLER_29_2254 ();
 sg13g2_decap_8 FILLER_29_2261 ();
 sg13g2_decap_8 FILLER_29_2268 ();
 sg13g2_decap_8 FILLER_29_2275 ();
 sg13g2_decap_8 FILLER_29_2282 ();
 sg13g2_decap_8 FILLER_29_2289 ();
 sg13g2_decap_8 FILLER_29_2296 ();
 sg13g2_decap_8 FILLER_29_2303 ();
 sg13g2_decap_8 FILLER_29_2310 ();
 sg13g2_decap_8 FILLER_29_2317 ();
 sg13g2_decap_8 FILLER_29_2324 ();
 sg13g2_decap_8 FILLER_29_2331 ();
 sg13g2_decap_8 FILLER_29_2338 ();
 sg13g2_decap_8 FILLER_29_2345 ();
 sg13g2_decap_8 FILLER_29_2352 ();
 sg13g2_decap_8 FILLER_29_2359 ();
 sg13g2_decap_8 FILLER_29_2366 ();
 sg13g2_decap_8 FILLER_29_2373 ();
 sg13g2_decap_8 FILLER_29_2380 ();
 sg13g2_decap_8 FILLER_29_2387 ();
 sg13g2_decap_8 FILLER_29_2394 ();
 sg13g2_decap_8 FILLER_29_2401 ();
 sg13g2_decap_8 FILLER_29_2408 ();
 sg13g2_decap_8 FILLER_29_2415 ();
 sg13g2_decap_8 FILLER_29_2422 ();
 sg13g2_decap_8 FILLER_29_2429 ();
 sg13g2_decap_8 FILLER_29_2436 ();
 sg13g2_decap_8 FILLER_29_2443 ();
 sg13g2_decap_8 FILLER_29_2450 ();
 sg13g2_decap_8 FILLER_29_2457 ();
 sg13g2_decap_8 FILLER_29_2464 ();
 sg13g2_decap_8 FILLER_29_2471 ();
 sg13g2_decap_8 FILLER_29_2478 ();
 sg13g2_decap_8 FILLER_29_2485 ();
 sg13g2_decap_8 FILLER_29_2492 ();
 sg13g2_decap_8 FILLER_29_2499 ();
 sg13g2_decap_8 FILLER_29_2506 ();
 sg13g2_decap_8 FILLER_29_2513 ();
 sg13g2_decap_8 FILLER_29_2520 ();
 sg13g2_decap_8 FILLER_29_2527 ();
 sg13g2_decap_8 FILLER_29_2534 ();
 sg13g2_decap_8 FILLER_29_2541 ();
 sg13g2_decap_8 FILLER_29_2548 ();
 sg13g2_decap_8 FILLER_29_2555 ();
 sg13g2_decap_8 FILLER_29_2562 ();
 sg13g2_decap_8 FILLER_29_2569 ();
 sg13g2_decap_8 FILLER_29_2576 ();
 sg13g2_decap_8 FILLER_29_2583 ();
 sg13g2_decap_8 FILLER_29_2590 ();
 sg13g2_decap_8 FILLER_29_2597 ();
 sg13g2_decap_8 FILLER_29_2604 ();
 sg13g2_decap_8 FILLER_29_2611 ();
 sg13g2_decap_8 FILLER_29_2618 ();
 sg13g2_decap_8 FILLER_29_2625 ();
 sg13g2_decap_8 FILLER_29_2632 ();
 sg13g2_decap_8 FILLER_29_2639 ();
 sg13g2_decap_8 FILLER_29_2646 ();
 sg13g2_decap_8 FILLER_29_2653 ();
 sg13g2_decap_8 FILLER_29_2660 ();
 sg13g2_decap_8 FILLER_29_2667 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_11 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_85 ();
 sg13g2_decap_4 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_394 ();
 sg13g2_fill_2 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_451 ();
 sg13g2_fill_2 FILLER_30_502 ();
 sg13g2_fill_2 FILLER_30_533 ();
 sg13g2_fill_1 FILLER_30_535 ();
 sg13g2_fill_2 FILLER_30_541 ();
 sg13g2_fill_1 FILLER_30_543 ();
 sg13g2_decap_8 FILLER_30_565 ();
 sg13g2_fill_1 FILLER_30_572 ();
 sg13g2_decap_4 FILLER_30_606 ();
 sg13g2_fill_1 FILLER_30_610 ();
 sg13g2_fill_2 FILLER_30_616 ();
 sg13g2_fill_2 FILLER_30_632 ();
 sg13g2_fill_2 FILLER_30_662 ();
 sg13g2_fill_1 FILLER_30_664 ();
 sg13g2_decap_4 FILLER_30_672 ();
 sg13g2_fill_1 FILLER_30_676 ();
 sg13g2_decap_4 FILLER_30_696 ();
 sg13g2_fill_1 FILLER_30_700 ();
 sg13g2_fill_2 FILLER_30_740 ();
 sg13g2_fill_1 FILLER_30_742 ();
 sg13g2_fill_1 FILLER_30_776 ();
 sg13g2_fill_1 FILLER_30_796 ();
 sg13g2_fill_1 FILLER_30_851 ();
 sg13g2_fill_2 FILLER_30_880 ();
 sg13g2_fill_1 FILLER_30_927 ();
 sg13g2_fill_2 FILLER_30_983 ();
 sg13g2_decap_8 FILLER_30_1010 ();
 sg13g2_decap_8 FILLER_30_1017 ();
 sg13g2_decap_8 FILLER_30_1024 ();
 sg13g2_fill_2 FILLER_30_1031 ();
 sg13g2_decap_8 FILLER_30_1036 ();
 sg13g2_decap_8 FILLER_30_1043 ();
 sg13g2_decap_8 FILLER_30_1085 ();
 sg13g2_decap_4 FILLER_30_1092 ();
 sg13g2_fill_2 FILLER_30_1105 ();
 sg13g2_fill_1 FILLER_30_1107 ();
 sg13g2_fill_1 FILLER_30_1113 ();
 sg13g2_fill_1 FILLER_30_1159 ();
 sg13g2_decap_8 FILLER_30_1181 ();
 sg13g2_fill_1 FILLER_30_1188 ();
 sg13g2_fill_2 FILLER_30_1321 ();
 sg13g2_fill_1 FILLER_30_1323 ();
 sg13g2_fill_2 FILLER_30_1337 ();
 sg13g2_fill_1 FILLER_30_1367 ();
 sg13g2_decap_4 FILLER_30_1378 ();
 sg13g2_decap_4 FILLER_30_1393 ();
 sg13g2_fill_2 FILLER_30_1424 ();
 sg13g2_fill_1 FILLER_30_1426 ();
 sg13g2_decap_4 FILLER_30_1468 ();
 sg13g2_decap_8 FILLER_30_1494 ();
 sg13g2_fill_2 FILLER_30_1501 ();
 sg13g2_fill_1 FILLER_30_1558 ();
 sg13g2_fill_1 FILLER_30_1575 ();
 sg13g2_decap_4 FILLER_30_1665 ();
 sg13g2_fill_1 FILLER_30_1714 ();
 sg13g2_fill_2 FILLER_30_1749 ();
 sg13g2_decap_4 FILLER_30_1827 ();
 sg13g2_decap_8 FILLER_30_1858 ();
 sg13g2_decap_8 FILLER_30_1865 ();
 sg13g2_fill_1 FILLER_30_1872 ();
 sg13g2_decap_4 FILLER_30_1882 ();
 sg13g2_fill_1 FILLER_30_1886 ();
 sg13g2_decap_4 FILLER_30_1891 ();
 sg13g2_decap_4 FILLER_30_1993 ();
 sg13g2_fill_1 FILLER_30_2013 ();
 sg13g2_fill_1 FILLER_30_2055 ();
 sg13g2_decap_8 FILLER_30_2106 ();
 sg13g2_fill_2 FILLER_30_2113 ();
 sg13g2_fill_1 FILLER_30_2164 ();
 sg13g2_fill_2 FILLER_30_2169 ();
 sg13g2_fill_2 FILLER_30_2225 ();
 sg13g2_fill_2 FILLER_30_2240 ();
 sg13g2_fill_1 FILLER_30_2242 ();
 sg13g2_decap_8 FILLER_30_2252 ();
 sg13g2_decap_8 FILLER_30_2259 ();
 sg13g2_decap_8 FILLER_30_2266 ();
 sg13g2_decap_8 FILLER_30_2273 ();
 sg13g2_decap_8 FILLER_30_2280 ();
 sg13g2_decap_8 FILLER_30_2287 ();
 sg13g2_decap_8 FILLER_30_2294 ();
 sg13g2_decap_8 FILLER_30_2301 ();
 sg13g2_decap_8 FILLER_30_2308 ();
 sg13g2_decap_8 FILLER_30_2315 ();
 sg13g2_decap_8 FILLER_30_2322 ();
 sg13g2_decap_8 FILLER_30_2329 ();
 sg13g2_decap_8 FILLER_30_2336 ();
 sg13g2_decap_8 FILLER_30_2343 ();
 sg13g2_decap_8 FILLER_30_2350 ();
 sg13g2_decap_8 FILLER_30_2357 ();
 sg13g2_decap_8 FILLER_30_2364 ();
 sg13g2_decap_8 FILLER_30_2371 ();
 sg13g2_decap_8 FILLER_30_2378 ();
 sg13g2_decap_8 FILLER_30_2385 ();
 sg13g2_decap_8 FILLER_30_2392 ();
 sg13g2_decap_8 FILLER_30_2399 ();
 sg13g2_decap_8 FILLER_30_2406 ();
 sg13g2_decap_8 FILLER_30_2413 ();
 sg13g2_decap_8 FILLER_30_2420 ();
 sg13g2_decap_8 FILLER_30_2427 ();
 sg13g2_decap_8 FILLER_30_2434 ();
 sg13g2_decap_8 FILLER_30_2441 ();
 sg13g2_decap_8 FILLER_30_2448 ();
 sg13g2_decap_8 FILLER_30_2455 ();
 sg13g2_decap_8 FILLER_30_2462 ();
 sg13g2_decap_8 FILLER_30_2469 ();
 sg13g2_decap_8 FILLER_30_2476 ();
 sg13g2_decap_8 FILLER_30_2483 ();
 sg13g2_decap_8 FILLER_30_2490 ();
 sg13g2_decap_8 FILLER_30_2497 ();
 sg13g2_decap_8 FILLER_30_2504 ();
 sg13g2_decap_8 FILLER_30_2511 ();
 sg13g2_decap_8 FILLER_30_2518 ();
 sg13g2_decap_8 FILLER_30_2525 ();
 sg13g2_decap_8 FILLER_30_2532 ();
 sg13g2_decap_8 FILLER_30_2539 ();
 sg13g2_decap_8 FILLER_30_2546 ();
 sg13g2_decap_8 FILLER_30_2553 ();
 sg13g2_decap_8 FILLER_30_2560 ();
 sg13g2_decap_8 FILLER_30_2567 ();
 sg13g2_decap_8 FILLER_30_2574 ();
 sg13g2_decap_8 FILLER_30_2581 ();
 sg13g2_decap_8 FILLER_30_2588 ();
 sg13g2_decap_8 FILLER_30_2595 ();
 sg13g2_decap_8 FILLER_30_2602 ();
 sg13g2_decap_8 FILLER_30_2609 ();
 sg13g2_decap_8 FILLER_30_2616 ();
 sg13g2_decap_8 FILLER_30_2623 ();
 sg13g2_decap_8 FILLER_30_2630 ();
 sg13g2_decap_8 FILLER_30_2637 ();
 sg13g2_decap_8 FILLER_30_2644 ();
 sg13g2_decap_8 FILLER_30_2651 ();
 sg13g2_decap_8 FILLER_30_2658 ();
 sg13g2_decap_8 FILLER_30_2665 ();
 sg13g2_fill_2 FILLER_30_2672 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_160 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_457 ();
 sg13g2_fill_1 FILLER_31_459 ();
 sg13g2_decap_8 FILLER_31_482 ();
 sg13g2_decap_8 FILLER_31_489 ();
 sg13g2_fill_2 FILLER_31_514 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_2 FILLER_31_535 ();
 sg13g2_fill_1 FILLER_31_537 ();
 sg13g2_decap_8 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_fill_2 FILLER_31_563 ();
 sg13g2_fill_1 FILLER_31_565 ();
 sg13g2_fill_2 FILLER_31_597 ();
 sg13g2_decap_8 FILLER_31_631 ();
 sg13g2_decap_8 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_645 ();
 sg13g2_decap_4 FILLER_31_652 ();
 sg13g2_fill_1 FILLER_31_676 ();
 sg13g2_decap_8 FILLER_31_704 ();
 sg13g2_fill_2 FILLER_31_728 ();
 sg13g2_fill_1 FILLER_31_730 ();
 sg13g2_fill_1 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_763 ();
 sg13g2_fill_2 FILLER_31_777 ();
 sg13g2_fill_2 FILLER_31_801 ();
 sg13g2_fill_1 FILLER_31_803 ();
 sg13g2_fill_2 FILLER_31_850 ();
 sg13g2_fill_1 FILLER_31_852 ();
 sg13g2_decap_4 FILLER_31_1003 ();
 sg13g2_decap_4 FILLER_31_1043 ();
 sg13g2_fill_2 FILLER_31_1047 ();
 sg13g2_decap_4 FILLER_31_1053 ();
 sg13g2_fill_1 FILLER_31_1057 ();
 sg13g2_decap_8 FILLER_31_1083 ();
 sg13g2_fill_1 FILLER_31_1090 ();
 sg13g2_decap_8 FILLER_31_1095 ();
 sg13g2_fill_1 FILLER_31_1102 ();
 sg13g2_fill_2 FILLER_31_1108 ();
 sg13g2_fill_1 FILLER_31_1110 ();
 sg13g2_decap_8 FILLER_31_1131 ();
 sg13g2_fill_2 FILLER_31_1138 ();
 sg13g2_fill_1 FILLER_31_1178 ();
 sg13g2_fill_2 FILLER_31_1223 ();
 sg13g2_fill_1 FILLER_31_1225 ();
 sg13g2_fill_2 FILLER_31_1269 ();
 sg13g2_fill_2 FILLER_31_1279 ();
 sg13g2_fill_2 FILLER_31_1290 ();
 sg13g2_fill_1 FILLER_31_1302 ();
 sg13g2_fill_2 FILLER_31_1315 ();
 sg13g2_fill_1 FILLER_31_1317 ();
 sg13g2_fill_1 FILLER_31_1328 ();
 sg13g2_decap_8 FILLER_31_1342 ();
 sg13g2_decap_8 FILLER_31_1349 ();
 sg13g2_fill_1 FILLER_31_1383 ();
 sg13g2_decap_4 FILLER_31_1389 ();
 sg13g2_fill_1 FILLER_31_1393 ();
 sg13g2_decap_4 FILLER_31_1439 ();
 sg13g2_fill_2 FILLER_31_1443 ();
 sg13g2_decap_8 FILLER_31_1458 ();
 sg13g2_decap_4 FILLER_31_1465 ();
 sg13g2_fill_2 FILLER_31_1469 ();
 sg13g2_fill_2 FILLER_31_1505 ();
 sg13g2_fill_1 FILLER_31_1544 ();
 sg13g2_decap_4 FILLER_31_1555 ();
 sg13g2_fill_2 FILLER_31_1576 ();
 sg13g2_decap_4 FILLER_31_1609 ();
 sg13g2_fill_1 FILLER_31_1631 ();
 sg13g2_fill_2 FILLER_31_1711 ();
 sg13g2_fill_1 FILLER_31_1713 ();
 sg13g2_decap_8 FILLER_31_1740 ();
 sg13g2_decap_4 FILLER_31_1747 ();
 sg13g2_fill_2 FILLER_31_1751 ();
 sg13g2_fill_1 FILLER_31_1786 ();
 sg13g2_fill_2 FILLER_31_1814 ();
 sg13g2_decap_8 FILLER_31_1869 ();
 sg13g2_decap_4 FILLER_31_1876 ();
 sg13g2_fill_2 FILLER_31_1880 ();
 sg13g2_decap_4 FILLER_31_1887 ();
 sg13g2_fill_2 FILLER_31_1891 ();
 sg13g2_fill_1 FILLER_31_1941 ();
 sg13g2_fill_2 FILLER_31_2003 ();
 sg13g2_fill_2 FILLER_31_2031 ();
 sg13g2_fill_1 FILLER_31_2033 ();
 sg13g2_decap_4 FILLER_31_2061 ();
 sg13g2_fill_1 FILLER_31_2065 ();
 sg13g2_fill_1 FILLER_31_2098 ();
 sg13g2_fill_1 FILLER_31_2112 ();
 sg13g2_fill_2 FILLER_31_2137 ();
 sg13g2_fill_2 FILLER_31_2149 ();
 sg13g2_fill_1 FILLER_31_2168 ();
 sg13g2_decap_4 FILLER_31_2218 ();
 sg13g2_fill_1 FILLER_31_2222 ();
 sg13g2_decap_8 FILLER_31_2256 ();
 sg13g2_decap_8 FILLER_31_2263 ();
 sg13g2_decap_8 FILLER_31_2270 ();
 sg13g2_decap_8 FILLER_31_2277 ();
 sg13g2_decap_8 FILLER_31_2284 ();
 sg13g2_decap_8 FILLER_31_2291 ();
 sg13g2_decap_8 FILLER_31_2298 ();
 sg13g2_decap_8 FILLER_31_2305 ();
 sg13g2_decap_8 FILLER_31_2312 ();
 sg13g2_decap_8 FILLER_31_2319 ();
 sg13g2_decap_8 FILLER_31_2326 ();
 sg13g2_decap_8 FILLER_31_2333 ();
 sg13g2_decap_8 FILLER_31_2340 ();
 sg13g2_decap_8 FILLER_31_2347 ();
 sg13g2_decap_8 FILLER_31_2354 ();
 sg13g2_decap_8 FILLER_31_2361 ();
 sg13g2_decap_8 FILLER_31_2368 ();
 sg13g2_decap_8 FILLER_31_2375 ();
 sg13g2_decap_8 FILLER_31_2382 ();
 sg13g2_decap_8 FILLER_31_2389 ();
 sg13g2_decap_8 FILLER_31_2396 ();
 sg13g2_decap_8 FILLER_31_2403 ();
 sg13g2_decap_8 FILLER_31_2410 ();
 sg13g2_decap_8 FILLER_31_2417 ();
 sg13g2_decap_8 FILLER_31_2424 ();
 sg13g2_decap_8 FILLER_31_2431 ();
 sg13g2_decap_8 FILLER_31_2438 ();
 sg13g2_decap_8 FILLER_31_2445 ();
 sg13g2_decap_8 FILLER_31_2452 ();
 sg13g2_decap_8 FILLER_31_2459 ();
 sg13g2_decap_8 FILLER_31_2466 ();
 sg13g2_decap_8 FILLER_31_2473 ();
 sg13g2_decap_8 FILLER_31_2480 ();
 sg13g2_decap_8 FILLER_31_2487 ();
 sg13g2_decap_8 FILLER_31_2494 ();
 sg13g2_decap_8 FILLER_31_2501 ();
 sg13g2_decap_8 FILLER_31_2508 ();
 sg13g2_decap_8 FILLER_31_2515 ();
 sg13g2_decap_8 FILLER_31_2522 ();
 sg13g2_decap_8 FILLER_31_2529 ();
 sg13g2_decap_8 FILLER_31_2536 ();
 sg13g2_decap_8 FILLER_31_2543 ();
 sg13g2_decap_8 FILLER_31_2550 ();
 sg13g2_decap_8 FILLER_31_2557 ();
 sg13g2_decap_8 FILLER_31_2564 ();
 sg13g2_decap_8 FILLER_31_2571 ();
 sg13g2_decap_8 FILLER_31_2578 ();
 sg13g2_decap_8 FILLER_31_2585 ();
 sg13g2_decap_8 FILLER_31_2592 ();
 sg13g2_decap_8 FILLER_31_2599 ();
 sg13g2_decap_8 FILLER_31_2606 ();
 sg13g2_decap_8 FILLER_31_2613 ();
 sg13g2_decap_8 FILLER_31_2620 ();
 sg13g2_decap_8 FILLER_31_2627 ();
 sg13g2_decap_8 FILLER_31_2634 ();
 sg13g2_decap_8 FILLER_31_2641 ();
 sg13g2_decap_8 FILLER_31_2648 ();
 sg13g2_decap_8 FILLER_31_2655 ();
 sg13g2_decap_8 FILLER_31_2662 ();
 sg13g2_decap_4 FILLER_31_2669 ();
 sg13g2_fill_1 FILLER_31_2673 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_1 FILLER_32_34 ();
 sg13g2_decap_4 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_fill_1 FILLER_32_457 ();
 sg13g2_fill_2 FILLER_32_461 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_4 FILLER_32_490 ();
 sg13g2_fill_2 FILLER_32_494 ();
 sg13g2_decap_8 FILLER_32_529 ();
 sg13g2_decap_4 FILLER_32_536 ();
 sg13g2_fill_1 FILLER_32_540 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_fill_2 FILLER_32_564 ();
 sg13g2_fill_2 FILLER_32_614 ();
 sg13g2_fill_2 FILLER_32_635 ();
 sg13g2_decap_8 FILLER_32_645 ();
 sg13g2_decap_4 FILLER_32_652 ();
 sg13g2_fill_2 FILLER_32_656 ();
 sg13g2_fill_1 FILLER_32_676 ();
 sg13g2_fill_1 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_710 ();
 sg13g2_decap_4 FILLER_32_717 ();
 sg13g2_decap_8 FILLER_32_725 ();
 sg13g2_fill_1 FILLER_32_764 ();
 sg13g2_fill_2 FILLER_32_774 ();
 sg13g2_fill_2 FILLER_32_848 ();
 sg13g2_fill_2 FILLER_32_859 ();
 sg13g2_fill_2 FILLER_32_925 ();
 sg13g2_fill_1 FILLER_32_927 ();
 sg13g2_fill_2 FILLER_32_961 ();
 sg13g2_fill_1 FILLER_32_963 ();
 sg13g2_fill_1 FILLER_32_977 ();
 sg13g2_decap_8 FILLER_32_1006 ();
 sg13g2_fill_1 FILLER_32_1013 ();
 sg13g2_fill_1 FILLER_32_1025 ();
 sg13g2_decap_8 FILLER_32_1031 ();
 sg13g2_fill_1 FILLER_32_1038 ();
 sg13g2_decap_4 FILLER_32_1044 ();
 sg13g2_fill_1 FILLER_32_1048 ();
 sg13g2_fill_2 FILLER_32_1079 ();
 sg13g2_fill_1 FILLER_32_1094 ();
 sg13g2_fill_2 FILLER_32_1099 ();
 sg13g2_fill_1 FILLER_32_1101 ();
 sg13g2_decap_4 FILLER_32_1136 ();
 sg13g2_fill_1 FILLER_32_1140 ();
 sg13g2_decap_8 FILLER_32_1150 ();
 sg13g2_decap_8 FILLER_32_1157 ();
 sg13g2_decap_8 FILLER_32_1164 ();
 sg13g2_decap_4 FILLER_32_1171 ();
 sg13g2_fill_2 FILLER_32_1194 ();
 sg13g2_fill_2 FILLER_32_1211 ();
 sg13g2_fill_1 FILLER_32_1245 ();
 sg13g2_decap_8 FILLER_32_1336 ();
 sg13g2_decap_8 FILLER_32_1343 ();
 sg13g2_decap_8 FILLER_32_1350 ();
 sg13g2_fill_2 FILLER_32_1375 ();
 sg13g2_fill_1 FILLER_32_1377 ();
 sg13g2_fill_2 FILLER_32_1416 ();
 sg13g2_decap_8 FILLER_32_1431 ();
 sg13g2_decap_8 FILLER_32_1438 ();
 sg13g2_fill_2 FILLER_32_1445 ();
 sg13g2_fill_1 FILLER_32_1447 ();
 sg13g2_fill_1 FILLER_32_1457 ();
 sg13g2_fill_2 FILLER_32_1504 ();
 sg13g2_fill_1 FILLER_32_1506 ();
 sg13g2_fill_1 FILLER_32_1563 ();
 sg13g2_fill_2 FILLER_32_1573 ();
 sg13g2_fill_1 FILLER_32_1575 ();
 sg13g2_fill_1 FILLER_32_1631 ();
 sg13g2_fill_1 FILLER_32_1668 ();
 sg13g2_decap_4 FILLER_32_1714 ();
 sg13g2_fill_1 FILLER_32_1718 ();
 sg13g2_decap_8 FILLER_32_1737 ();
 sg13g2_decap_8 FILLER_32_1744 ();
 sg13g2_fill_1 FILLER_32_1751 ();
 sg13g2_fill_1 FILLER_32_1776 ();
 sg13g2_fill_1 FILLER_32_1850 ();
 sg13g2_decap_4 FILLER_32_1864 ();
 sg13g2_fill_2 FILLER_32_1901 ();
 sg13g2_fill_1 FILLER_32_1903 ();
 sg13g2_fill_2 FILLER_32_1981 ();
 sg13g2_fill_2 FILLER_32_2041 ();
 sg13g2_decap_8 FILLER_32_2049 ();
 sg13g2_decap_4 FILLER_32_2056 ();
 sg13g2_fill_1 FILLER_32_2060 ();
 sg13g2_decap_4 FILLER_32_2102 ();
 sg13g2_fill_2 FILLER_32_2219 ();
 sg13g2_decap_8 FILLER_32_2254 ();
 sg13g2_decap_8 FILLER_32_2261 ();
 sg13g2_decap_8 FILLER_32_2268 ();
 sg13g2_decap_8 FILLER_32_2275 ();
 sg13g2_decap_8 FILLER_32_2282 ();
 sg13g2_decap_8 FILLER_32_2289 ();
 sg13g2_decap_8 FILLER_32_2296 ();
 sg13g2_decap_8 FILLER_32_2303 ();
 sg13g2_decap_8 FILLER_32_2310 ();
 sg13g2_decap_8 FILLER_32_2317 ();
 sg13g2_decap_8 FILLER_32_2324 ();
 sg13g2_decap_8 FILLER_32_2331 ();
 sg13g2_decap_8 FILLER_32_2338 ();
 sg13g2_decap_8 FILLER_32_2345 ();
 sg13g2_decap_8 FILLER_32_2352 ();
 sg13g2_decap_8 FILLER_32_2359 ();
 sg13g2_decap_8 FILLER_32_2366 ();
 sg13g2_decap_8 FILLER_32_2373 ();
 sg13g2_decap_8 FILLER_32_2380 ();
 sg13g2_decap_8 FILLER_32_2387 ();
 sg13g2_decap_8 FILLER_32_2394 ();
 sg13g2_decap_8 FILLER_32_2401 ();
 sg13g2_decap_8 FILLER_32_2408 ();
 sg13g2_decap_8 FILLER_32_2415 ();
 sg13g2_decap_8 FILLER_32_2422 ();
 sg13g2_decap_8 FILLER_32_2429 ();
 sg13g2_decap_8 FILLER_32_2436 ();
 sg13g2_decap_8 FILLER_32_2443 ();
 sg13g2_decap_8 FILLER_32_2450 ();
 sg13g2_decap_8 FILLER_32_2457 ();
 sg13g2_decap_8 FILLER_32_2464 ();
 sg13g2_decap_8 FILLER_32_2471 ();
 sg13g2_decap_8 FILLER_32_2478 ();
 sg13g2_decap_8 FILLER_32_2485 ();
 sg13g2_decap_8 FILLER_32_2492 ();
 sg13g2_decap_8 FILLER_32_2499 ();
 sg13g2_decap_8 FILLER_32_2506 ();
 sg13g2_decap_8 FILLER_32_2513 ();
 sg13g2_decap_8 FILLER_32_2520 ();
 sg13g2_decap_8 FILLER_32_2527 ();
 sg13g2_decap_8 FILLER_32_2534 ();
 sg13g2_decap_8 FILLER_32_2541 ();
 sg13g2_decap_8 FILLER_32_2548 ();
 sg13g2_decap_8 FILLER_32_2555 ();
 sg13g2_decap_8 FILLER_32_2562 ();
 sg13g2_decap_8 FILLER_32_2569 ();
 sg13g2_decap_8 FILLER_32_2576 ();
 sg13g2_decap_8 FILLER_32_2583 ();
 sg13g2_decap_8 FILLER_32_2590 ();
 sg13g2_decap_8 FILLER_32_2597 ();
 sg13g2_decap_8 FILLER_32_2604 ();
 sg13g2_decap_8 FILLER_32_2611 ();
 sg13g2_decap_8 FILLER_32_2618 ();
 sg13g2_decap_8 FILLER_32_2625 ();
 sg13g2_decap_8 FILLER_32_2632 ();
 sg13g2_decap_8 FILLER_32_2639 ();
 sg13g2_decap_8 FILLER_32_2646 ();
 sg13g2_decap_8 FILLER_32_2653 ();
 sg13g2_decap_8 FILLER_32_2660 ();
 sg13g2_decap_8 FILLER_32_2667 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_decap_8 FILLER_33_127 ();
 sg13g2_decap_4 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_447 ();
 sg13g2_fill_2 FILLER_33_451 ();
 sg13g2_decap_8 FILLER_33_521 ();
 sg13g2_decap_8 FILLER_33_528 ();
 sg13g2_fill_2 FILLER_33_535 ();
 sg13g2_fill_1 FILLER_33_537 ();
 sg13g2_fill_1 FILLER_33_553 ();
 sg13g2_fill_1 FILLER_33_559 ();
 sg13g2_fill_1 FILLER_33_566 ();
 sg13g2_fill_2 FILLER_33_583 ();
 sg13g2_fill_1 FILLER_33_585 ();
 sg13g2_fill_1 FILLER_33_597 ();
 sg13g2_fill_2 FILLER_33_625 ();
 sg13g2_fill_2 FILLER_33_633 ();
 sg13g2_fill_1 FILLER_33_673 ();
 sg13g2_decap_4 FILLER_33_705 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_fill_1 FILLER_33_728 ();
 sg13g2_fill_1 FILLER_33_734 ();
 sg13g2_decap_8 FILLER_33_740 ();
 sg13g2_decap_8 FILLER_33_747 ();
 sg13g2_decap_4 FILLER_33_754 ();
 sg13g2_fill_1 FILLER_33_758 ();
 sg13g2_decap_8 FILLER_33_762 ();
 sg13g2_fill_1 FILLER_33_769 ();
 sg13g2_fill_1 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_858 ();
 sg13g2_decap_8 FILLER_33_865 ();
 sg13g2_fill_1 FILLER_33_872 ();
 sg13g2_fill_2 FILLER_33_877 ();
 sg13g2_fill_1 FILLER_33_884 ();
 sg13g2_decap_4 FILLER_33_920 ();
 sg13g2_decap_4 FILLER_33_928 ();
 sg13g2_fill_1 FILLER_33_932 ();
 sg13g2_fill_2 FILLER_33_942 ();
 sg13g2_decap_4 FILLER_33_948 ();
 sg13g2_fill_1 FILLER_33_952 ();
 sg13g2_fill_2 FILLER_33_962 ();
 sg13g2_fill_1 FILLER_33_964 ();
 sg13g2_fill_1 FILLER_33_983 ();
 sg13g2_decap_4 FILLER_33_1050 ();
 sg13g2_fill_2 FILLER_33_1054 ();
 sg13g2_fill_2 FILLER_33_1115 ();
 sg13g2_fill_2 FILLER_33_1134 ();
 sg13g2_decap_8 FILLER_33_1141 ();
 sg13g2_fill_1 FILLER_33_1148 ();
 sg13g2_decap_8 FILLER_33_1158 ();
 sg13g2_decap_4 FILLER_33_1165 ();
 sg13g2_fill_1 FILLER_33_1169 ();
 sg13g2_decap_4 FILLER_33_1208 ();
 sg13g2_fill_1 FILLER_33_1212 ();
 sg13g2_fill_1 FILLER_33_1234 ();
 sg13g2_fill_2 FILLER_33_1257 ();
 sg13g2_decap_8 FILLER_33_1332 ();
 sg13g2_decap_8 FILLER_33_1339 ();
 sg13g2_decap_4 FILLER_33_1375 ();
 sg13g2_decap_8 FILLER_33_1403 ();
 sg13g2_decap_4 FILLER_33_1410 ();
 sg13g2_fill_2 FILLER_33_1427 ();
 sg13g2_decap_4 FILLER_33_1485 ();
 sg13g2_fill_2 FILLER_33_1507 ();
 sg13g2_fill_2 FILLER_33_1518 ();
 sg13g2_fill_1 FILLER_33_1595 ();
 sg13g2_fill_2 FILLER_33_1607 ();
 sg13g2_fill_1 FILLER_33_1647 ();
 sg13g2_fill_1 FILLER_33_1750 ();
 sg13g2_fill_1 FILLER_33_1812 ();
 sg13g2_decap_8 FILLER_33_1858 ();
 sg13g2_fill_1 FILLER_33_1919 ();
 sg13g2_fill_2 FILLER_33_1971 ();
 sg13g2_fill_1 FILLER_33_2028 ();
 sg13g2_decap_8 FILLER_33_2051 ();
 sg13g2_decap_4 FILLER_33_2058 ();
 sg13g2_fill_2 FILLER_33_2123 ();
 sg13g2_decap_8 FILLER_33_2219 ();
 sg13g2_fill_2 FILLER_33_2226 ();
 sg13g2_fill_2 FILLER_33_2232 ();
 sg13g2_fill_1 FILLER_33_2234 ();
 sg13g2_decap_8 FILLER_33_2257 ();
 sg13g2_decap_8 FILLER_33_2264 ();
 sg13g2_decap_8 FILLER_33_2271 ();
 sg13g2_decap_8 FILLER_33_2278 ();
 sg13g2_decap_8 FILLER_33_2285 ();
 sg13g2_decap_8 FILLER_33_2292 ();
 sg13g2_decap_8 FILLER_33_2299 ();
 sg13g2_decap_8 FILLER_33_2306 ();
 sg13g2_decap_8 FILLER_33_2313 ();
 sg13g2_decap_8 FILLER_33_2320 ();
 sg13g2_decap_8 FILLER_33_2327 ();
 sg13g2_decap_8 FILLER_33_2334 ();
 sg13g2_decap_8 FILLER_33_2341 ();
 sg13g2_decap_4 FILLER_33_2348 ();
 sg13g2_fill_1 FILLER_33_2352 ();
 sg13g2_decap_8 FILLER_33_2357 ();
 sg13g2_decap_8 FILLER_33_2364 ();
 sg13g2_decap_8 FILLER_33_2371 ();
 sg13g2_decap_8 FILLER_33_2378 ();
 sg13g2_decap_8 FILLER_33_2385 ();
 sg13g2_decap_8 FILLER_33_2392 ();
 sg13g2_decap_8 FILLER_33_2399 ();
 sg13g2_decap_8 FILLER_33_2406 ();
 sg13g2_decap_8 FILLER_33_2413 ();
 sg13g2_decap_8 FILLER_33_2420 ();
 sg13g2_decap_8 FILLER_33_2427 ();
 sg13g2_decap_8 FILLER_33_2434 ();
 sg13g2_decap_8 FILLER_33_2441 ();
 sg13g2_decap_8 FILLER_33_2448 ();
 sg13g2_decap_8 FILLER_33_2455 ();
 sg13g2_decap_8 FILLER_33_2462 ();
 sg13g2_decap_8 FILLER_33_2469 ();
 sg13g2_decap_8 FILLER_33_2476 ();
 sg13g2_decap_8 FILLER_33_2483 ();
 sg13g2_decap_8 FILLER_33_2490 ();
 sg13g2_decap_8 FILLER_33_2497 ();
 sg13g2_decap_8 FILLER_33_2504 ();
 sg13g2_decap_8 FILLER_33_2511 ();
 sg13g2_decap_8 FILLER_33_2518 ();
 sg13g2_decap_8 FILLER_33_2525 ();
 sg13g2_decap_8 FILLER_33_2532 ();
 sg13g2_decap_8 FILLER_33_2539 ();
 sg13g2_decap_8 FILLER_33_2546 ();
 sg13g2_decap_8 FILLER_33_2553 ();
 sg13g2_decap_8 FILLER_33_2560 ();
 sg13g2_decap_8 FILLER_33_2567 ();
 sg13g2_decap_8 FILLER_33_2574 ();
 sg13g2_decap_8 FILLER_33_2581 ();
 sg13g2_decap_8 FILLER_33_2588 ();
 sg13g2_decap_8 FILLER_33_2595 ();
 sg13g2_decap_8 FILLER_33_2602 ();
 sg13g2_decap_8 FILLER_33_2609 ();
 sg13g2_decap_8 FILLER_33_2616 ();
 sg13g2_decap_8 FILLER_33_2623 ();
 sg13g2_decap_8 FILLER_33_2630 ();
 sg13g2_decap_8 FILLER_33_2637 ();
 sg13g2_decap_8 FILLER_33_2644 ();
 sg13g2_decap_8 FILLER_33_2651 ();
 sg13g2_decap_8 FILLER_33_2658 ();
 sg13g2_decap_8 FILLER_33_2665 ();
 sg13g2_fill_2 FILLER_33_2672 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_fill_1 FILLER_34_64 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_decap_4 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_478 ();
 sg13g2_decap_8 FILLER_34_496 ();
 sg13g2_fill_1 FILLER_34_503 ();
 sg13g2_decap_8 FILLER_34_509 ();
 sg13g2_decap_8 FILLER_34_516 ();
 sg13g2_fill_2 FILLER_34_523 ();
 sg13g2_fill_1 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_562 ();
 sg13g2_decap_8 FILLER_34_569 ();
 sg13g2_fill_2 FILLER_34_576 ();
 sg13g2_fill_2 FILLER_34_583 ();
 sg13g2_fill_1 FILLER_34_585 ();
 sg13g2_fill_2 FILLER_34_596 ();
 sg13g2_fill_1 FILLER_34_598 ();
 sg13g2_fill_2 FILLER_34_604 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_4 FILLER_34_651 ();
 sg13g2_fill_2 FILLER_34_665 ();
 sg13g2_fill_2 FILLER_34_676 ();
 sg13g2_fill_1 FILLER_34_678 ();
 sg13g2_decap_8 FILLER_34_702 ();
 sg13g2_fill_1 FILLER_34_709 ();
 sg13g2_fill_1 FILLER_34_720 ();
 sg13g2_fill_2 FILLER_34_740 ();
 sg13g2_fill_1 FILLER_34_748 ();
 sg13g2_fill_2 FILLER_34_786 ();
 sg13g2_decap_4 FILLER_34_819 ();
 sg13g2_fill_1 FILLER_34_823 ();
 sg13g2_fill_2 FILLER_34_833 ();
 sg13g2_decap_4 FILLER_34_857 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_34_899 ();
 sg13g2_decap_8 FILLER_34_906 ();
 sg13g2_decap_8 FILLER_34_913 ();
 sg13g2_decap_8 FILLER_34_920 ();
 sg13g2_decap_8 FILLER_34_927 ();
 sg13g2_decap_8 FILLER_34_934 ();
 sg13g2_fill_2 FILLER_34_941 ();
 sg13g2_decap_4 FILLER_34_970 ();
 sg13g2_decap_4 FILLER_34_1015 ();
 sg13g2_decap_4 FILLER_34_1047 ();
 sg13g2_fill_2 FILLER_34_1051 ();
 sg13g2_fill_1 FILLER_34_1067 ();
 sg13g2_fill_2 FILLER_34_1085 ();
 sg13g2_decap_8 FILLER_34_1092 ();
 sg13g2_decap_4 FILLER_34_1099 ();
 sg13g2_fill_1 FILLER_34_1103 ();
 sg13g2_fill_2 FILLER_34_1115 ();
 sg13g2_decap_4 FILLER_34_1176 ();
 sg13g2_fill_1 FILLER_34_1180 ();
 sg13g2_fill_2 FILLER_34_1208 ();
 sg13g2_fill_1 FILLER_34_1210 ();
 sg13g2_fill_1 FILLER_34_1263 ();
 sg13g2_fill_1 FILLER_34_1279 ();
 sg13g2_fill_2 FILLER_34_1294 ();
 sg13g2_fill_1 FILLER_34_1296 ();
 sg13g2_fill_1 FILLER_34_1310 ();
 sg13g2_fill_2 FILLER_34_1335 ();
 sg13g2_fill_2 FILLER_34_1365 ();
 sg13g2_fill_1 FILLER_34_1367 ();
 sg13g2_decap_4 FILLER_34_1413 ();
 sg13g2_fill_1 FILLER_34_1417 ();
 sg13g2_fill_1 FILLER_34_1446 ();
 sg13g2_fill_2 FILLER_34_1546 ();
 sg13g2_fill_2 FILLER_34_1598 ();
 sg13g2_fill_1 FILLER_34_1618 ();
 sg13g2_fill_2 FILLER_34_1655 ();
 sg13g2_decap_8 FILLER_34_1700 ();
 sg13g2_fill_1 FILLER_34_1784 ();
 sg13g2_fill_1 FILLER_34_1817 ();
 sg13g2_decap_4 FILLER_34_1857 ();
 sg13g2_fill_1 FILLER_34_1861 ();
 sg13g2_fill_2 FILLER_34_1951 ();
 sg13g2_fill_1 FILLER_34_2020 ();
 sg13g2_fill_2 FILLER_34_2054 ();
 sg13g2_fill_1 FILLER_34_2056 ();
 sg13g2_fill_2 FILLER_34_2173 ();
 sg13g2_fill_1 FILLER_34_2175 ();
 sg13g2_decap_8 FILLER_34_2224 ();
 sg13g2_decap_8 FILLER_34_2244 ();
 sg13g2_decap_8 FILLER_34_2251 ();
 sg13g2_decap_8 FILLER_34_2258 ();
 sg13g2_decap_8 FILLER_34_2265 ();
 sg13g2_decap_8 FILLER_34_2272 ();
 sg13g2_decap_8 FILLER_34_2279 ();
 sg13g2_decap_8 FILLER_34_2286 ();
 sg13g2_decap_8 FILLER_34_2293 ();
 sg13g2_decap_8 FILLER_34_2300 ();
 sg13g2_decap_8 FILLER_34_2307 ();
 sg13g2_decap_8 FILLER_34_2314 ();
 sg13g2_decap_8 FILLER_34_2321 ();
 sg13g2_decap_8 FILLER_34_2328 ();
 sg13g2_decap_8 FILLER_34_2335 ();
 sg13g2_fill_2 FILLER_34_2342 ();
 sg13g2_fill_2 FILLER_34_2352 ();
 sg13g2_decap_4 FILLER_34_2371 ();
 sg13g2_decap_8 FILLER_34_2378 ();
 sg13g2_fill_2 FILLER_34_2389 ();
 sg13g2_fill_2 FILLER_34_2395 ();
 sg13g2_fill_1 FILLER_34_2397 ();
 sg13g2_decap_4 FILLER_34_2402 ();
 sg13g2_fill_1 FILLER_34_2406 ();
 sg13g2_decap_8 FILLER_34_2411 ();
 sg13g2_decap_8 FILLER_34_2418 ();
 sg13g2_decap_8 FILLER_34_2425 ();
 sg13g2_decap_8 FILLER_34_2432 ();
 sg13g2_decap_8 FILLER_34_2439 ();
 sg13g2_decap_8 FILLER_34_2446 ();
 sg13g2_decap_8 FILLER_34_2453 ();
 sg13g2_decap_8 FILLER_34_2460 ();
 sg13g2_decap_8 FILLER_34_2467 ();
 sg13g2_decap_8 FILLER_34_2474 ();
 sg13g2_decap_8 FILLER_34_2481 ();
 sg13g2_decap_8 FILLER_34_2488 ();
 sg13g2_decap_8 FILLER_34_2495 ();
 sg13g2_decap_8 FILLER_34_2502 ();
 sg13g2_decap_8 FILLER_34_2509 ();
 sg13g2_decap_8 FILLER_34_2516 ();
 sg13g2_decap_8 FILLER_34_2523 ();
 sg13g2_decap_8 FILLER_34_2530 ();
 sg13g2_decap_8 FILLER_34_2537 ();
 sg13g2_decap_8 FILLER_34_2544 ();
 sg13g2_decap_8 FILLER_34_2551 ();
 sg13g2_decap_8 FILLER_34_2558 ();
 sg13g2_decap_8 FILLER_34_2565 ();
 sg13g2_decap_8 FILLER_34_2572 ();
 sg13g2_decap_8 FILLER_34_2579 ();
 sg13g2_decap_8 FILLER_34_2586 ();
 sg13g2_decap_8 FILLER_34_2593 ();
 sg13g2_decap_8 FILLER_34_2600 ();
 sg13g2_decap_8 FILLER_34_2607 ();
 sg13g2_decap_8 FILLER_34_2614 ();
 sg13g2_decap_8 FILLER_34_2621 ();
 sg13g2_decap_8 FILLER_34_2628 ();
 sg13g2_decap_8 FILLER_34_2635 ();
 sg13g2_decap_8 FILLER_34_2642 ();
 sg13g2_decap_8 FILLER_34_2649 ();
 sg13g2_decap_8 FILLER_34_2656 ();
 sg13g2_decap_8 FILLER_34_2663 ();
 sg13g2_decap_4 FILLER_34_2670 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_47 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_fill_1 FILLER_35_430 ();
 sg13g2_fill_2 FILLER_35_444 ();
 sg13g2_fill_1 FILLER_35_446 ();
 sg13g2_decap_8 FILLER_35_496 ();
 sg13g2_decap_8 FILLER_35_503 ();
 sg13g2_fill_2 FILLER_35_510 ();
 sg13g2_fill_1 FILLER_35_512 ();
 sg13g2_fill_2 FILLER_35_536 ();
 sg13g2_fill_2 FILLER_35_549 ();
 sg13g2_fill_1 FILLER_35_551 ();
 sg13g2_decap_8 FILLER_35_562 ();
 sg13g2_decap_8 FILLER_35_569 ();
 sg13g2_decap_4 FILLER_35_576 ();
 sg13g2_fill_2 FILLER_35_580 ();
 sg13g2_fill_1 FILLER_35_590 ();
 sg13g2_fill_2 FILLER_35_600 ();
 sg13g2_fill_1 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_631 ();
 sg13g2_decap_8 FILLER_35_638 ();
 sg13g2_decap_8 FILLER_35_671 ();
 sg13g2_decap_4 FILLER_35_678 ();
 sg13g2_fill_1 FILLER_35_682 ();
 sg13g2_decap_8 FILLER_35_688 ();
 sg13g2_decap_8 FILLER_35_695 ();
 sg13g2_decap_8 FILLER_35_702 ();
 sg13g2_fill_1 FILLER_35_733 ();
 sg13g2_fill_2 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_764 ();
 sg13g2_fill_2 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_814 ();
 sg13g2_fill_1 FILLER_35_821 ();
 sg13g2_decap_4 FILLER_35_835 ();
 sg13g2_fill_2 FILLER_35_877 ();
 sg13g2_decap_8 FILLER_35_912 ();
 sg13g2_decap_8 FILLER_35_919 ();
 sg13g2_decap_8 FILLER_35_926 ();
 sg13g2_decap_4 FILLER_35_933 ();
 sg13g2_decap_4 FILLER_35_1008 ();
 sg13g2_fill_1 FILLER_35_1012 ();
 sg13g2_fill_2 FILLER_35_1034 ();
 sg13g2_fill_2 FILLER_35_1063 ();
 sg13g2_fill_2 FILLER_35_1076 ();
 sg13g2_fill_1 FILLER_35_1078 ();
 sg13g2_decap_8 FILLER_35_1093 ();
 sg13g2_decap_4 FILLER_35_1100 ();
 sg13g2_decap_8 FILLER_35_1152 ();
 sg13g2_decap_4 FILLER_35_1159 ();
 sg13g2_fill_2 FILLER_35_1163 ();
 sg13g2_decap_4 FILLER_35_1181 ();
 sg13g2_fill_1 FILLER_35_1185 ();
 sg13g2_fill_1 FILLER_35_1249 ();
 sg13g2_fill_1 FILLER_35_1278 ();
 sg13g2_fill_1 FILLER_35_1283 ();
 sg13g2_decap_8 FILLER_35_1326 ();
 sg13g2_fill_1 FILLER_35_1333 ();
 sg13g2_fill_2 FILLER_35_1356 ();
 sg13g2_decap_4 FILLER_35_1382 ();
 sg13g2_fill_1 FILLER_35_1396 ();
 sg13g2_fill_2 FILLER_35_1424 ();
 sg13g2_fill_1 FILLER_35_1440 ();
 sg13g2_fill_2 FILLER_35_1459 ();
 sg13g2_fill_1 FILLER_35_1461 ();
 sg13g2_fill_2 FILLER_35_1515 ();
 sg13g2_fill_1 FILLER_35_1517 ();
 sg13g2_fill_2 FILLER_35_1541 ();
 sg13g2_fill_1 FILLER_35_1543 ();
 sg13g2_fill_2 FILLER_35_1587 ();
 sg13g2_fill_1 FILLER_35_1589 ();
 sg13g2_fill_1 FILLER_35_1643 ();
 sg13g2_decap_8 FILLER_35_1693 ();
 sg13g2_decap_4 FILLER_35_1700 ();
 sg13g2_fill_1 FILLER_35_1704 ();
 sg13g2_fill_2 FILLER_35_1730 ();
 sg13g2_fill_2 FILLER_35_1745 ();
 sg13g2_fill_1 FILLER_35_1747 ();
 sg13g2_fill_1 FILLER_35_1799 ();
 sg13g2_fill_2 FILLER_35_1818 ();
 sg13g2_fill_1 FILLER_35_1820 ();
 sg13g2_fill_1 FILLER_35_1849 ();
 sg13g2_fill_1 FILLER_35_1859 ();
 sg13g2_fill_2 FILLER_35_1970 ();
 sg13g2_fill_2 FILLER_35_2072 ();
 sg13g2_fill_1 FILLER_35_2079 ();
 sg13g2_decap_8 FILLER_35_2093 ();
 sg13g2_fill_1 FILLER_35_2100 ();
 sg13g2_fill_1 FILLER_35_2114 ();
 sg13g2_fill_1 FILLER_35_2135 ();
 sg13g2_fill_2 FILLER_35_2151 ();
 sg13g2_fill_1 FILLER_35_2153 ();
 sg13g2_decap_4 FILLER_35_2164 ();
 sg13g2_fill_1 FILLER_35_2168 ();
 sg13g2_fill_1 FILLER_35_2227 ();
 sg13g2_decap_8 FILLER_35_2233 ();
 sg13g2_decap_8 FILLER_35_2240 ();
 sg13g2_decap_8 FILLER_35_2247 ();
 sg13g2_decap_8 FILLER_35_2254 ();
 sg13g2_decap_8 FILLER_35_2261 ();
 sg13g2_decap_8 FILLER_35_2268 ();
 sg13g2_decap_8 FILLER_35_2275 ();
 sg13g2_decap_8 FILLER_35_2282 ();
 sg13g2_decap_8 FILLER_35_2289 ();
 sg13g2_decap_8 FILLER_35_2296 ();
 sg13g2_decap_8 FILLER_35_2303 ();
 sg13g2_decap_8 FILLER_35_2310 ();
 sg13g2_decap_8 FILLER_35_2317 ();
 sg13g2_decap_8 FILLER_35_2324 ();
 sg13g2_decap_8 FILLER_35_2331 ();
 sg13g2_fill_1 FILLER_35_2338 ();
 sg13g2_fill_2 FILLER_35_2348 ();
 sg13g2_decap_4 FILLER_35_2415 ();
 sg13g2_fill_1 FILLER_35_2419 ();
 sg13g2_decap_8 FILLER_35_2429 ();
 sg13g2_decap_8 FILLER_35_2436 ();
 sg13g2_decap_8 FILLER_35_2443 ();
 sg13g2_decap_8 FILLER_35_2450 ();
 sg13g2_decap_8 FILLER_35_2457 ();
 sg13g2_decap_8 FILLER_35_2464 ();
 sg13g2_decap_8 FILLER_35_2471 ();
 sg13g2_decap_8 FILLER_35_2478 ();
 sg13g2_decap_8 FILLER_35_2485 ();
 sg13g2_decap_8 FILLER_35_2492 ();
 sg13g2_decap_8 FILLER_35_2499 ();
 sg13g2_decap_8 FILLER_35_2506 ();
 sg13g2_decap_8 FILLER_35_2513 ();
 sg13g2_decap_8 FILLER_35_2520 ();
 sg13g2_decap_8 FILLER_35_2527 ();
 sg13g2_decap_8 FILLER_35_2534 ();
 sg13g2_decap_8 FILLER_35_2541 ();
 sg13g2_decap_8 FILLER_35_2548 ();
 sg13g2_decap_8 FILLER_35_2555 ();
 sg13g2_decap_8 FILLER_35_2562 ();
 sg13g2_decap_8 FILLER_35_2569 ();
 sg13g2_decap_8 FILLER_35_2576 ();
 sg13g2_decap_8 FILLER_35_2583 ();
 sg13g2_decap_8 FILLER_35_2590 ();
 sg13g2_decap_8 FILLER_35_2597 ();
 sg13g2_decap_8 FILLER_35_2604 ();
 sg13g2_decap_8 FILLER_35_2611 ();
 sg13g2_decap_8 FILLER_35_2618 ();
 sg13g2_decap_8 FILLER_35_2625 ();
 sg13g2_decap_8 FILLER_35_2632 ();
 sg13g2_decap_8 FILLER_35_2639 ();
 sg13g2_decap_8 FILLER_35_2646 ();
 sg13g2_decap_8 FILLER_35_2653 ();
 sg13g2_decap_8 FILLER_35_2660 ();
 sg13g2_decap_8 FILLER_35_2667 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_4 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_decap_4 FILLER_36_193 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_4 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_395 ();
 sg13g2_fill_1 FILLER_36_405 ();
 sg13g2_fill_1 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_36_442 ();
 sg13g2_fill_2 FILLER_36_449 ();
 sg13g2_fill_1 FILLER_36_482 ();
 sg13g2_decap_4 FILLER_36_509 ();
 sg13g2_fill_2 FILLER_36_513 ();
 sg13g2_fill_2 FILLER_36_527 ();
 sg13g2_fill_1 FILLER_36_529 ();
 sg13g2_decap_8 FILLER_36_565 ();
 sg13g2_decap_4 FILLER_36_572 ();
 sg13g2_fill_1 FILLER_36_588 ();
 sg13g2_fill_2 FILLER_36_625 ();
 sg13g2_decap_4 FILLER_36_635 ();
 sg13g2_fill_1 FILLER_36_639 ();
 sg13g2_decap_8 FILLER_36_668 ();
 sg13g2_decap_8 FILLER_36_675 ();
 sg13g2_fill_2 FILLER_36_682 ();
 sg13g2_fill_1 FILLER_36_684 ();
 sg13g2_decap_8 FILLER_36_691 ();
 sg13g2_decap_8 FILLER_36_698 ();
 sg13g2_decap_8 FILLER_36_705 ();
 sg13g2_decap_4 FILLER_36_712 ();
 sg13g2_fill_1 FILLER_36_716 ();
 sg13g2_fill_1 FILLER_36_738 ();
 sg13g2_decap_4 FILLER_36_746 ();
 sg13g2_fill_1 FILLER_36_750 ();
 sg13g2_decap_4 FILLER_36_764 ();
 sg13g2_decap_8 FILLER_36_794 ();
 sg13g2_fill_1 FILLER_36_801 ();
 sg13g2_decap_4 FILLER_36_828 ();
 sg13g2_fill_2 FILLER_36_862 ();
 sg13g2_fill_2 FILLER_36_872 ();
 sg13g2_fill_1 FILLER_36_880 ();
 sg13g2_fill_2 FILLER_36_959 ();
 sg13g2_fill_2 FILLER_36_1003 ();
 sg13g2_fill_2 FILLER_36_1045 ();
 sg13g2_fill_1 FILLER_36_1047 ();
 sg13g2_fill_2 FILLER_36_1053 ();
 sg13g2_fill_1 FILLER_36_1055 ();
 sg13g2_fill_2 FILLER_36_1079 ();
 sg13g2_fill_1 FILLER_36_1081 ();
 sg13g2_decap_8 FILLER_36_1098 ();
 sg13g2_fill_1 FILLER_36_1105 ();
 sg13g2_fill_2 FILLER_36_1154 ();
 sg13g2_fill_2 FILLER_36_1163 ();
 sg13g2_fill_2 FILLER_36_1294 ();
 sg13g2_fill_2 FILLER_36_1309 ();
 sg13g2_fill_1 FILLER_36_1311 ();
 sg13g2_decap_8 FILLER_36_1326 ();
 sg13g2_fill_2 FILLER_36_1333 ();
 sg13g2_fill_1 FILLER_36_1335 ();
 sg13g2_fill_1 FILLER_36_1363 ();
 sg13g2_decap_4 FILLER_36_1373 ();
 sg13g2_decap_4 FILLER_36_1412 ();
 sg13g2_fill_2 FILLER_36_1443 ();
 sg13g2_fill_1 FILLER_36_1445 ();
 sg13g2_fill_1 FILLER_36_1497 ();
 sg13g2_fill_2 FILLER_36_1511 ();
 sg13g2_fill_1 FILLER_36_1544 ();
 sg13g2_fill_2 FILLER_36_1564 ();
 sg13g2_fill_1 FILLER_36_1566 ();
 sg13g2_fill_2 FILLER_36_1576 ();
 sg13g2_fill_1 FILLER_36_1578 ();
 sg13g2_fill_2 FILLER_36_1615 ();
 sg13g2_fill_2 FILLER_36_1628 ();
 sg13g2_decap_8 FILLER_36_1689 ();
 sg13g2_decap_8 FILLER_36_1696 ();
 sg13g2_fill_2 FILLER_36_1703 ();
 sg13g2_fill_2 FILLER_36_1748 ();
 sg13g2_fill_1 FILLER_36_1750 ();
 sg13g2_fill_1 FILLER_36_1807 ();
 sg13g2_fill_2 FILLER_36_1853 ();
 sg13g2_fill_1 FILLER_36_1855 ();
 sg13g2_fill_1 FILLER_36_1884 ();
 sg13g2_decap_4 FILLER_36_1943 ();
 sg13g2_fill_1 FILLER_36_1960 ();
 sg13g2_decap_4 FILLER_36_1989 ();
 sg13g2_fill_2 FILLER_36_2036 ();
 sg13g2_fill_1 FILLER_36_2078 ();
 sg13g2_decap_8 FILLER_36_2091 ();
 sg13g2_decap_8 FILLER_36_2098 ();
 sg13g2_decap_8 FILLER_36_2105 ();
 sg13g2_fill_2 FILLER_36_2112 ();
 sg13g2_fill_1 FILLER_36_2114 ();
 sg13g2_fill_2 FILLER_36_2123 ();
 sg13g2_fill_1 FILLER_36_2162 ();
 sg13g2_decap_8 FILLER_36_2199 ();
 sg13g2_decap_8 FILLER_36_2247 ();
 sg13g2_decap_4 FILLER_36_2254 ();
 sg13g2_fill_1 FILLER_36_2258 ();
 sg13g2_decap_8 FILLER_36_2271 ();
 sg13g2_decap_8 FILLER_36_2278 ();
 sg13g2_decap_8 FILLER_36_2285 ();
 sg13g2_decap_8 FILLER_36_2292 ();
 sg13g2_decap_8 FILLER_36_2299 ();
 sg13g2_decap_8 FILLER_36_2306 ();
 sg13g2_decap_8 FILLER_36_2317 ();
 sg13g2_decap_8 FILLER_36_2324 ();
 sg13g2_fill_2 FILLER_36_2331 ();
 sg13g2_fill_2 FILLER_36_2343 ();
 sg13g2_fill_2 FILLER_36_2373 ();
 sg13g2_decap_8 FILLER_36_2434 ();
 sg13g2_decap_8 FILLER_36_2441 ();
 sg13g2_decap_8 FILLER_36_2448 ();
 sg13g2_decap_8 FILLER_36_2455 ();
 sg13g2_decap_8 FILLER_36_2462 ();
 sg13g2_decap_8 FILLER_36_2469 ();
 sg13g2_decap_8 FILLER_36_2476 ();
 sg13g2_decap_8 FILLER_36_2483 ();
 sg13g2_decap_8 FILLER_36_2490 ();
 sg13g2_decap_8 FILLER_36_2497 ();
 sg13g2_decap_8 FILLER_36_2504 ();
 sg13g2_decap_8 FILLER_36_2511 ();
 sg13g2_decap_8 FILLER_36_2518 ();
 sg13g2_decap_8 FILLER_36_2525 ();
 sg13g2_decap_8 FILLER_36_2532 ();
 sg13g2_decap_8 FILLER_36_2539 ();
 sg13g2_decap_8 FILLER_36_2546 ();
 sg13g2_decap_8 FILLER_36_2553 ();
 sg13g2_decap_8 FILLER_36_2560 ();
 sg13g2_decap_8 FILLER_36_2567 ();
 sg13g2_decap_8 FILLER_36_2574 ();
 sg13g2_decap_8 FILLER_36_2581 ();
 sg13g2_decap_8 FILLER_36_2588 ();
 sg13g2_decap_8 FILLER_36_2595 ();
 sg13g2_decap_8 FILLER_36_2602 ();
 sg13g2_decap_8 FILLER_36_2609 ();
 sg13g2_decap_8 FILLER_36_2616 ();
 sg13g2_decap_8 FILLER_36_2623 ();
 sg13g2_decap_8 FILLER_36_2630 ();
 sg13g2_decap_8 FILLER_36_2637 ();
 sg13g2_decap_8 FILLER_36_2644 ();
 sg13g2_decap_8 FILLER_36_2651 ();
 sg13g2_decap_8 FILLER_36_2658 ();
 sg13g2_decap_8 FILLER_36_2665 ();
 sg13g2_fill_2 FILLER_36_2672 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_30 ();
 sg13g2_fill_1 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_4 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_409 ();
 sg13g2_decap_8 FILLER_37_416 ();
 sg13g2_decap_8 FILLER_37_423 ();
 sg13g2_fill_2 FILLER_37_430 ();
 sg13g2_fill_2 FILLER_37_475 ();
 sg13g2_fill_2 FILLER_37_504 ();
 sg13g2_fill_1 FILLER_37_506 ();
 sg13g2_decap_8 FILLER_37_512 ();
 sg13g2_fill_2 FILLER_37_536 ();
 sg13g2_fill_1 FILLER_37_538 ();
 sg13g2_decap_8 FILLER_37_549 ();
 sg13g2_decap_4 FILLER_37_556 ();
 sg13g2_fill_1 FILLER_37_560 ();
 sg13g2_decap_4 FILLER_37_565 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_fill_1 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_fill_2 FILLER_37_672 ();
 sg13g2_fill_1 FILLER_37_674 ();
 sg13g2_decap_8 FILLER_37_697 ();
 sg13g2_fill_2 FILLER_37_704 ();
 sg13g2_decap_4 FILLER_37_723 ();
 sg13g2_fill_2 FILLER_37_727 ();
 sg13g2_fill_1 FILLER_37_736 ();
 sg13g2_fill_2 FILLER_37_752 ();
 sg13g2_fill_2 FILLER_37_760 ();
 sg13g2_decap_4 FILLER_37_795 ();
 sg13g2_fill_2 FILLER_37_799 ();
 sg13g2_fill_1 FILLER_37_920 ();
 sg13g2_decap_4 FILLER_37_941 ();
 sg13g2_fill_2 FILLER_37_971 ();
 sg13g2_fill_1 FILLER_37_978 ();
 sg13g2_fill_2 FILLER_37_1006 ();
 sg13g2_fill_1 FILLER_37_1008 ();
 sg13g2_fill_2 FILLER_37_1015 ();
 sg13g2_fill_1 FILLER_37_1017 ();
 sg13g2_fill_2 FILLER_37_1027 ();
 sg13g2_fill_2 FILLER_37_1063 ();
 sg13g2_fill_1 FILLER_37_1065 ();
 sg13g2_decap_8 FILLER_37_1087 ();
 sg13g2_decap_4 FILLER_37_1094 ();
 sg13g2_fill_2 FILLER_37_1098 ();
 sg13g2_decap_4 FILLER_37_1105 ();
 sg13g2_fill_2 FILLER_37_1109 ();
 sg13g2_decap_4 FILLER_37_1166 ();
 sg13g2_fill_2 FILLER_37_1170 ();
 sg13g2_fill_1 FILLER_37_1258 ();
 sg13g2_decap_8 FILLER_37_1322 ();
 sg13g2_decap_4 FILLER_37_1329 ();
 sg13g2_fill_2 FILLER_37_1333 ();
 sg13g2_decap_4 FILLER_37_1340 ();
 sg13g2_fill_2 FILLER_37_1344 ();
 sg13g2_decap_4 FILLER_37_1366 ();
 sg13g2_fill_2 FILLER_37_1375 ();
 sg13g2_fill_2 FILLER_37_1399 ();
 sg13g2_fill_1 FILLER_37_1401 ();
 sg13g2_fill_2 FILLER_37_1416 ();
 sg13g2_fill_1 FILLER_37_1418 ();
 sg13g2_fill_1 FILLER_37_1422 ();
 sg13g2_fill_2 FILLER_37_1449 ();
 sg13g2_fill_1 FILLER_37_1451 ();
 sg13g2_decap_4 FILLER_37_1479 ();
 sg13g2_fill_2 FILLER_37_1502 ();
 sg13g2_fill_1 FILLER_37_1504 ();
 sg13g2_fill_2 FILLER_37_1518 ();
 sg13g2_fill_2 FILLER_37_1551 ();
 sg13g2_fill_1 FILLER_37_1553 ();
 sg13g2_decap_8 FILLER_37_1584 ();
 sg13g2_fill_2 FILLER_37_1654 ();
 sg13g2_fill_1 FILLER_37_1656 ();
 sg13g2_decap_8 FILLER_37_1731 ();
 sg13g2_decap_8 FILLER_37_1738 ();
 sg13g2_decap_4 FILLER_37_1745 ();
 sg13g2_fill_2 FILLER_37_1749 ();
 sg13g2_fill_2 FILLER_37_1767 ();
 sg13g2_fill_1 FILLER_37_1769 ();
 sg13g2_fill_2 FILLER_37_1775 ();
 sg13g2_fill_1 FILLER_37_1777 ();
 sg13g2_decap_4 FILLER_37_1850 ();
 sg13g2_fill_1 FILLER_37_1854 ();
 sg13g2_fill_1 FILLER_37_1882 ();
 sg13g2_decap_4 FILLER_37_1935 ();
 sg13g2_fill_2 FILLER_37_1939 ();
 sg13g2_fill_2 FILLER_37_1946 ();
 sg13g2_fill_1 FILLER_37_1948 ();
 sg13g2_fill_1 FILLER_37_1965 ();
 sg13g2_fill_1 FILLER_37_1980 ();
 sg13g2_fill_2 FILLER_37_1990 ();
 sg13g2_fill_1 FILLER_37_2050 ();
 sg13g2_fill_2 FILLER_37_2074 ();
 sg13g2_decap_4 FILLER_37_2109 ();
 sg13g2_fill_1 FILLER_37_2113 ();
 sg13g2_fill_2 FILLER_37_2127 ();
 sg13g2_decap_8 FILLER_37_2183 ();
 sg13g2_decap_4 FILLER_37_2190 ();
 sg13g2_fill_1 FILLER_37_2194 ();
 sg13g2_fill_2 FILLER_37_2246 ();
 sg13g2_fill_1 FILLER_37_2248 ();
 sg13g2_decap_8 FILLER_37_2289 ();
 sg13g2_decap_8 FILLER_37_2296 ();
 sg13g2_decap_4 FILLER_37_2303 ();
 sg13g2_fill_1 FILLER_37_2307 ();
 sg13g2_fill_1 FILLER_37_2336 ();
 sg13g2_fill_1 FILLER_37_2405 ();
 sg13g2_decap_8 FILLER_37_2433 ();
 sg13g2_decap_8 FILLER_37_2440 ();
 sg13g2_decap_8 FILLER_37_2447 ();
 sg13g2_decap_8 FILLER_37_2454 ();
 sg13g2_decap_8 FILLER_37_2461 ();
 sg13g2_decap_8 FILLER_37_2468 ();
 sg13g2_decap_8 FILLER_37_2475 ();
 sg13g2_decap_8 FILLER_37_2482 ();
 sg13g2_decap_8 FILLER_37_2489 ();
 sg13g2_decap_8 FILLER_37_2496 ();
 sg13g2_decap_8 FILLER_37_2503 ();
 sg13g2_decap_8 FILLER_37_2510 ();
 sg13g2_decap_8 FILLER_37_2517 ();
 sg13g2_decap_8 FILLER_37_2524 ();
 sg13g2_decap_8 FILLER_37_2531 ();
 sg13g2_decap_8 FILLER_37_2538 ();
 sg13g2_decap_8 FILLER_37_2545 ();
 sg13g2_decap_8 FILLER_37_2552 ();
 sg13g2_decap_8 FILLER_37_2559 ();
 sg13g2_decap_8 FILLER_37_2566 ();
 sg13g2_decap_8 FILLER_37_2573 ();
 sg13g2_decap_8 FILLER_37_2580 ();
 sg13g2_decap_8 FILLER_37_2587 ();
 sg13g2_decap_8 FILLER_37_2594 ();
 sg13g2_decap_8 FILLER_37_2601 ();
 sg13g2_decap_8 FILLER_37_2608 ();
 sg13g2_decap_8 FILLER_37_2615 ();
 sg13g2_decap_8 FILLER_37_2622 ();
 sg13g2_decap_8 FILLER_37_2629 ();
 sg13g2_decap_8 FILLER_37_2636 ();
 sg13g2_decap_8 FILLER_37_2643 ();
 sg13g2_decap_8 FILLER_37_2650 ();
 sg13g2_decap_8 FILLER_37_2657 ();
 sg13g2_decap_8 FILLER_37_2664 ();
 sg13g2_fill_2 FILLER_37_2671 ();
 sg13g2_fill_1 FILLER_37_2673 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_120 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_318 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_38_443 ();
 sg13g2_fill_2 FILLER_38_486 ();
 sg13g2_fill_2 FILLER_38_507 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_fill_2 FILLER_38_525 ();
 sg13g2_fill_1 FILLER_38_527 ();
 sg13g2_fill_1 FILLER_38_537 ();
 sg13g2_decap_8 FILLER_38_542 ();
 sg13g2_decap_8 FILLER_38_549 ();
 sg13g2_fill_1 FILLER_38_556 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_fill_2 FILLER_38_626 ();
 sg13g2_decap_8 FILLER_38_638 ();
 sg13g2_decap_8 FILLER_38_645 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_2 FILLER_38_707 ();
 sg13g2_fill_1 FILLER_38_709 ();
 sg13g2_decap_8 FILLER_38_719 ();
 sg13g2_decap_4 FILLER_38_726 ();
 sg13g2_fill_2 FILLER_38_730 ();
 sg13g2_fill_1 FILLER_38_757 ();
 sg13g2_fill_1 FILLER_38_773 ();
 sg13g2_decap_8 FILLER_38_814 ();
 sg13g2_fill_2 FILLER_38_821 ();
 sg13g2_fill_1 FILLER_38_826 ();
 sg13g2_fill_2 FILLER_38_850 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_fill_1 FILLER_38_921 ();
 sg13g2_decap_4 FILLER_38_940 ();
 sg13g2_fill_1 FILLER_38_944 ();
 sg13g2_fill_2 FILLER_38_958 ();
 sg13g2_fill_2 FILLER_38_1043 ();
 sg13g2_fill_1 FILLER_38_1045 ();
 sg13g2_fill_2 FILLER_38_1060 ();
 sg13g2_fill_2 FILLER_38_1079 ();
 sg13g2_fill_1 FILLER_38_1081 ();
 sg13g2_fill_1 FILLER_38_1087 ();
 sg13g2_fill_1 FILLER_38_1093 ();
 sg13g2_decap_4 FILLER_38_1115 ();
 sg13g2_decap_8 FILLER_38_1140 ();
 sg13g2_decap_8 FILLER_38_1147 ();
 sg13g2_decap_8 FILLER_38_1154 ();
 sg13g2_decap_4 FILLER_38_1161 ();
 sg13g2_fill_2 FILLER_38_1165 ();
 sg13g2_fill_2 FILLER_38_1211 ();
 sg13g2_fill_2 FILLER_38_1246 ();
 sg13g2_decap_4 FILLER_38_1284 ();
 sg13g2_fill_2 FILLER_38_1345 ();
 sg13g2_fill_1 FILLER_38_1389 ();
 sg13g2_fill_2 FILLER_38_1400 ();
 sg13g2_decap_8 FILLER_38_1416 ();
 sg13g2_decap_4 FILLER_38_1423 ();
 sg13g2_fill_1 FILLER_38_1464 ();
 sg13g2_fill_2 FILLER_38_1505 ();
 sg13g2_decap_4 FILLER_38_1595 ();
 sg13g2_fill_2 FILLER_38_1599 ();
 sg13g2_fill_1 FILLER_38_1623 ();
 sg13g2_fill_1 FILLER_38_1661 ();
 sg13g2_fill_2 FILLER_38_1721 ();
 sg13g2_decap_4 FILLER_38_1750 ();
 sg13g2_fill_2 FILLER_38_1754 ();
 sg13g2_fill_1 FILLER_38_1778 ();
 sg13g2_decap_4 FILLER_38_1863 ();
 sg13g2_fill_2 FILLER_38_1867 ();
 sg13g2_fill_2 FILLER_38_1878 ();
 sg13g2_fill_1 FILLER_38_1880 ();
 sg13g2_fill_2 FILLER_38_1948 ();
 sg13g2_fill_1 FILLER_38_1950 ();
 sg13g2_fill_2 FILLER_38_1980 ();
 sg13g2_fill_1 FILLER_38_1982 ();
 sg13g2_fill_2 FILLER_38_2019 ();
 sg13g2_fill_2 FILLER_38_2030 ();
 sg13g2_fill_1 FILLER_38_2057 ();
 sg13g2_decap_8 FILLER_38_2119 ();
 sg13g2_decap_4 FILLER_38_2126 ();
 sg13g2_fill_1 FILLER_38_2130 ();
 sg13g2_decap_8 FILLER_38_2154 ();
 sg13g2_decap_4 FILLER_38_2161 ();
 sg13g2_decap_4 FILLER_38_2174 ();
 sg13g2_fill_1 FILLER_38_2178 ();
 sg13g2_fill_2 FILLER_38_2201 ();
 sg13g2_fill_1 FILLER_38_2203 ();
 sg13g2_fill_2 FILLER_38_2218 ();
 sg13g2_decap_8 FILLER_38_2299 ();
 sg13g2_decap_4 FILLER_38_2306 ();
 sg13g2_fill_1 FILLER_38_2374 ();
 sg13g2_decap_8 FILLER_38_2437 ();
 sg13g2_decap_8 FILLER_38_2444 ();
 sg13g2_decap_8 FILLER_38_2451 ();
 sg13g2_decap_8 FILLER_38_2458 ();
 sg13g2_decap_8 FILLER_38_2465 ();
 sg13g2_decap_8 FILLER_38_2472 ();
 sg13g2_decap_8 FILLER_38_2479 ();
 sg13g2_decap_8 FILLER_38_2486 ();
 sg13g2_decap_8 FILLER_38_2493 ();
 sg13g2_decap_8 FILLER_38_2500 ();
 sg13g2_decap_8 FILLER_38_2507 ();
 sg13g2_decap_8 FILLER_38_2514 ();
 sg13g2_decap_8 FILLER_38_2521 ();
 sg13g2_decap_8 FILLER_38_2528 ();
 sg13g2_decap_8 FILLER_38_2535 ();
 sg13g2_decap_8 FILLER_38_2542 ();
 sg13g2_decap_8 FILLER_38_2549 ();
 sg13g2_decap_8 FILLER_38_2556 ();
 sg13g2_decap_8 FILLER_38_2563 ();
 sg13g2_decap_8 FILLER_38_2570 ();
 sg13g2_decap_8 FILLER_38_2577 ();
 sg13g2_decap_8 FILLER_38_2584 ();
 sg13g2_decap_8 FILLER_38_2591 ();
 sg13g2_decap_8 FILLER_38_2598 ();
 sg13g2_decap_8 FILLER_38_2605 ();
 sg13g2_decap_8 FILLER_38_2612 ();
 sg13g2_decap_8 FILLER_38_2619 ();
 sg13g2_decap_8 FILLER_38_2626 ();
 sg13g2_decap_8 FILLER_38_2633 ();
 sg13g2_decap_8 FILLER_38_2640 ();
 sg13g2_decap_8 FILLER_38_2647 ();
 sg13g2_decap_8 FILLER_38_2654 ();
 sg13g2_decap_8 FILLER_38_2661 ();
 sg13g2_decap_4 FILLER_38_2668 ();
 sg13g2_fill_2 FILLER_38_2672 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_9 ();
 sg13g2_fill_2 FILLER_39_43 ();
 sg13g2_fill_1 FILLER_39_45 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_fill_2 FILLER_39_80 ();
 sg13g2_decap_4 FILLER_39_87 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_2 FILLER_39_166 ();
 sg13g2_fill_1 FILLER_39_168 ();
 sg13g2_fill_2 FILLER_39_232 ();
 sg13g2_fill_1 FILLER_39_234 ();
 sg13g2_fill_2 FILLER_39_285 ();
 sg13g2_fill_1 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_313 ();
 sg13g2_fill_2 FILLER_39_374 ();
 sg13g2_decap_8 FILLER_39_389 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_8 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_410 ();
 sg13g2_fill_2 FILLER_39_453 ();
 sg13g2_decap_8 FILLER_39_473 ();
 sg13g2_fill_2 FILLER_39_485 ();
 sg13g2_fill_1 FILLER_39_487 ();
 sg13g2_decap_8 FILLER_39_519 ();
 sg13g2_decap_4 FILLER_39_526 ();
 sg13g2_fill_2 FILLER_39_530 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_4 FILLER_39_543 ();
 sg13g2_fill_1 FILLER_39_547 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_4 FILLER_39_581 ();
 sg13g2_fill_2 FILLER_39_602 ();
 sg13g2_fill_1 FILLER_39_604 ();
 sg13g2_fill_1 FILLER_39_621 ();
 sg13g2_fill_1 FILLER_39_632 ();
 sg13g2_fill_2 FILLER_39_643 ();
 sg13g2_fill_1 FILLER_39_645 ();
 sg13g2_fill_2 FILLER_39_701 ();
 sg13g2_fill_1 FILLER_39_703 ();
 sg13g2_fill_2 FILLER_39_710 ();
 sg13g2_fill_1 FILLER_39_712 ();
 sg13g2_fill_2 FILLER_39_727 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_fill_1 FILLER_39_742 ();
 sg13g2_fill_1 FILLER_39_754 ();
 sg13g2_fill_1 FILLER_39_788 ();
 sg13g2_fill_2 FILLER_39_805 ();
 sg13g2_fill_2 FILLER_39_826 ();
 sg13g2_fill_1 FILLER_39_828 ();
 sg13g2_fill_2 FILLER_39_939 ();
 sg13g2_fill_1 FILLER_39_1024 ();
 sg13g2_decap_8 FILLER_39_1110 ();
 sg13g2_fill_1 FILLER_39_1117 ();
 sg13g2_decap_4 FILLER_39_1138 ();
 sg13g2_fill_2 FILLER_39_1142 ();
 sg13g2_decap_4 FILLER_39_1180 ();
 sg13g2_fill_1 FILLER_39_1276 ();
 sg13g2_decap_4 FILLER_39_1410 ();
 sg13g2_fill_2 FILLER_39_1414 ();
 sg13g2_fill_1 FILLER_39_1422 ();
 sg13g2_fill_1 FILLER_39_1446 ();
 sg13g2_fill_1 FILLER_39_1519 ();
 sg13g2_fill_1 FILLER_39_1549 ();
 sg13g2_decap_8 FILLER_39_1593 ();
 sg13g2_fill_2 FILLER_39_1605 ();
 sg13g2_fill_2 FILLER_39_1631 ();
 sg13g2_fill_1 FILLER_39_1633 ();
 sg13g2_fill_2 FILLER_39_1659 ();
 sg13g2_fill_2 FILLER_39_1677 ();
 sg13g2_fill_2 FILLER_39_1688 ();
 sg13g2_fill_1 FILLER_39_1751 ();
 sg13g2_fill_2 FILLER_39_1788 ();
 sg13g2_decap_8 FILLER_39_1876 ();
 sg13g2_decap_8 FILLER_39_1883 ();
 sg13g2_fill_2 FILLER_39_1890 ();
 sg13g2_fill_1 FILLER_39_1892 ();
 sg13g2_fill_1 FILLER_39_1947 ();
 sg13g2_fill_1 FILLER_39_1984 ();
 sg13g2_fill_1 FILLER_39_1997 ();
 sg13g2_fill_2 FILLER_39_2061 ();
 sg13g2_decap_8 FILLER_39_2119 ();
 sg13g2_decap_8 FILLER_39_2126 ();
 sg13g2_decap_4 FILLER_39_2143 ();
 sg13g2_decap_8 FILLER_39_2156 ();
 sg13g2_decap_4 FILLER_39_2163 ();
 sg13g2_fill_2 FILLER_39_2167 ();
 sg13g2_fill_2 FILLER_39_2216 ();
 sg13g2_fill_2 FILLER_39_2257 ();
 sg13g2_decap_4 FILLER_39_2303 ();
 sg13g2_fill_1 FILLER_39_2307 ();
 sg13g2_fill_2 FILLER_39_2340 ();
 sg13g2_fill_1 FILLER_39_2351 ();
 sg13g2_fill_2 FILLER_39_2384 ();
 sg13g2_decap_8 FILLER_39_2425 ();
 sg13g2_decap_8 FILLER_39_2432 ();
 sg13g2_decap_8 FILLER_39_2439 ();
 sg13g2_decap_8 FILLER_39_2446 ();
 sg13g2_decap_8 FILLER_39_2453 ();
 sg13g2_decap_8 FILLER_39_2460 ();
 sg13g2_decap_8 FILLER_39_2467 ();
 sg13g2_decap_8 FILLER_39_2474 ();
 sg13g2_decap_8 FILLER_39_2481 ();
 sg13g2_decap_8 FILLER_39_2488 ();
 sg13g2_decap_8 FILLER_39_2495 ();
 sg13g2_decap_8 FILLER_39_2502 ();
 sg13g2_decap_8 FILLER_39_2509 ();
 sg13g2_decap_8 FILLER_39_2516 ();
 sg13g2_decap_8 FILLER_39_2523 ();
 sg13g2_decap_8 FILLER_39_2530 ();
 sg13g2_decap_8 FILLER_39_2537 ();
 sg13g2_decap_8 FILLER_39_2544 ();
 sg13g2_decap_8 FILLER_39_2551 ();
 sg13g2_decap_8 FILLER_39_2558 ();
 sg13g2_decap_8 FILLER_39_2565 ();
 sg13g2_decap_8 FILLER_39_2572 ();
 sg13g2_decap_8 FILLER_39_2579 ();
 sg13g2_decap_8 FILLER_39_2586 ();
 sg13g2_decap_8 FILLER_39_2593 ();
 sg13g2_decap_8 FILLER_39_2600 ();
 sg13g2_decap_8 FILLER_39_2607 ();
 sg13g2_decap_8 FILLER_39_2614 ();
 sg13g2_decap_8 FILLER_39_2621 ();
 sg13g2_decap_8 FILLER_39_2628 ();
 sg13g2_decap_8 FILLER_39_2635 ();
 sg13g2_decap_8 FILLER_39_2642 ();
 sg13g2_decap_8 FILLER_39_2649 ();
 sg13g2_decap_8 FILLER_39_2656 ();
 sg13g2_decap_8 FILLER_39_2663 ();
 sg13g2_decap_4 FILLER_39_2670 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_25 ();
 sg13g2_fill_1 FILLER_40_40 ();
 sg13g2_decap_8 FILLER_40_51 ();
 sg13g2_fill_1 FILLER_40_58 ();
 sg13g2_decap_4 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_76 ();
 sg13g2_decap_8 FILLER_40_83 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_126 ();
 sg13g2_decap_4 FILLER_40_159 ();
 sg13g2_decap_8 FILLER_40_180 ();
 sg13g2_fill_1 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_228 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_fill_2 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_296 ();
 sg13g2_decap_4 FILLER_40_305 ();
 sg13g2_fill_2 FILLER_40_328 ();
 sg13g2_fill_1 FILLER_40_330 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_383 ();
 sg13g2_decap_4 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_decap_4 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_470 ();
 sg13g2_decap_8 FILLER_40_477 ();
 sg13g2_fill_2 FILLER_40_484 ();
 sg13g2_fill_1 FILLER_40_499 ();
 sg13g2_decap_4 FILLER_40_532 ();
 sg13g2_fill_2 FILLER_40_536 ();
 sg13g2_decap_8 FILLER_40_579 ();
 sg13g2_decap_8 FILLER_40_586 ();
 sg13g2_decap_4 FILLER_40_593 ();
 sg13g2_fill_2 FILLER_40_601 ();
 sg13g2_fill_2 FILLER_40_616 ();
 sg13g2_fill_1 FILLER_40_618 ();
 sg13g2_fill_2 FILLER_40_650 ();
 sg13g2_fill_1 FILLER_40_665 ();
 sg13g2_fill_2 FILLER_40_694 ();
 sg13g2_fill_1 FILLER_40_713 ();
 sg13g2_fill_1 FILLER_40_751 ();
 sg13g2_decap_8 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_fill_1 FILLER_40_794 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_fill_2 FILLER_40_830 ();
 sg13g2_fill_2 FILLER_40_840 ();
 sg13g2_fill_1 FILLER_40_868 ();
 sg13g2_fill_2 FILLER_40_884 ();
 sg13g2_fill_2 FILLER_40_901 ();
 sg13g2_fill_2 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_1059 ();
 sg13g2_decap_8 FILLER_40_1066 ();
 sg13g2_fill_1 FILLER_40_1090 ();
 sg13g2_decap_8 FILLER_40_1100 ();
 sg13g2_fill_2 FILLER_40_1107 ();
 sg13g2_decap_4 FILLER_40_1113 ();
 sg13g2_fill_1 FILLER_40_1125 ();
 sg13g2_decap_4 FILLER_40_1200 ();
 sg13g2_fill_2 FILLER_40_1204 ();
 sg13g2_fill_1 FILLER_40_1219 ();
 sg13g2_fill_2 FILLER_40_1266 ();
 sg13g2_fill_1 FILLER_40_1291 ();
 sg13g2_fill_2 FILLER_40_1300 ();
 sg13g2_fill_1 FILLER_40_1302 ();
 sg13g2_decap_4 FILLER_40_1322 ();
 sg13g2_decap_4 FILLER_40_1357 ();
 sg13g2_fill_1 FILLER_40_1407 ();
 sg13g2_fill_1 FILLER_40_1444 ();
 sg13g2_fill_2 FILLER_40_1464 ();
 sg13g2_fill_2 FILLER_40_1527 ();
 sg13g2_fill_1 FILLER_40_1545 ();
 sg13g2_fill_2 FILLER_40_1560 ();
 sg13g2_fill_1 FILLER_40_1562 ();
 sg13g2_decap_4 FILLER_40_1591 ();
 sg13g2_decap_4 FILLER_40_1724 ();
 sg13g2_fill_1 FILLER_40_1728 ();
 sg13g2_decap_4 FILLER_40_1738 ();
 sg13g2_fill_1 FILLER_40_1742 ();
 sg13g2_fill_2 FILLER_40_1788 ();
 sg13g2_fill_2 FILLER_40_1816 ();
 sg13g2_fill_1 FILLER_40_1818 ();
 sg13g2_fill_1 FILLER_40_1831 ();
 sg13g2_fill_2 FILLER_40_1847 ();
 sg13g2_decap_8 FILLER_40_1886 ();
 sg13g2_decap_8 FILLER_40_1893 ();
 sg13g2_fill_1 FILLER_40_1900 ();
 sg13g2_fill_1 FILLER_40_1989 ();
 sg13g2_fill_1 FILLER_40_2081 ();
 sg13g2_decap_8 FILLER_40_2129 ();
 sg13g2_decap_8 FILLER_40_2136 ();
 sg13g2_fill_1 FILLER_40_2143 ();
 sg13g2_decap_8 FILLER_40_2153 ();
 sg13g2_decap_4 FILLER_40_2160 ();
 sg13g2_fill_1 FILLER_40_2164 ();
 sg13g2_fill_1 FILLER_40_2175 ();
 sg13g2_decap_8 FILLER_40_2305 ();
 sg13g2_decap_4 FILLER_40_2312 ();
 sg13g2_fill_1 FILLER_40_2316 ();
 sg13g2_fill_2 FILLER_40_2333 ();
 sg13g2_fill_2 FILLER_40_2368 ();
 sg13g2_decap_8 FILLER_40_2419 ();
 sg13g2_decap_8 FILLER_40_2426 ();
 sg13g2_decap_8 FILLER_40_2433 ();
 sg13g2_decap_8 FILLER_40_2440 ();
 sg13g2_decap_8 FILLER_40_2447 ();
 sg13g2_decap_8 FILLER_40_2454 ();
 sg13g2_decap_8 FILLER_40_2461 ();
 sg13g2_decap_8 FILLER_40_2468 ();
 sg13g2_decap_8 FILLER_40_2475 ();
 sg13g2_decap_8 FILLER_40_2482 ();
 sg13g2_decap_8 FILLER_40_2489 ();
 sg13g2_decap_8 FILLER_40_2496 ();
 sg13g2_decap_8 FILLER_40_2503 ();
 sg13g2_decap_8 FILLER_40_2510 ();
 sg13g2_decap_8 FILLER_40_2517 ();
 sg13g2_decap_8 FILLER_40_2524 ();
 sg13g2_decap_8 FILLER_40_2531 ();
 sg13g2_decap_8 FILLER_40_2538 ();
 sg13g2_decap_8 FILLER_40_2545 ();
 sg13g2_decap_8 FILLER_40_2552 ();
 sg13g2_decap_8 FILLER_40_2559 ();
 sg13g2_decap_8 FILLER_40_2566 ();
 sg13g2_decap_8 FILLER_40_2573 ();
 sg13g2_decap_8 FILLER_40_2580 ();
 sg13g2_decap_8 FILLER_40_2587 ();
 sg13g2_decap_8 FILLER_40_2594 ();
 sg13g2_decap_8 FILLER_40_2601 ();
 sg13g2_decap_8 FILLER_40_2608 ();
 sg13g2_decap_8 FILLER_40_2615 ();
 sg13g2_decap_8 FILLER_40_2622 ();
 sg13g2_decap_8 FILLER_40_2629 ();
 sg13g2_decap_8 FILLER_40_2636 ();
 sg13g2_decap_8 FILLER_40_2643 ();
 sg13g2_decap_8 FILLER_40_2650 ();
 sg13g2_decap_8 FILLER_40_2657 ();
 sg13g2_decap_8 FILLER_40_2664 ();
 sg13g2_fill_2 FILLER_40_2671 ();
 sg13g2_fill_1 FILLER_40_2673 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_4 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_46 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_fill_2 FILLER_41_92 ();
 sg13g2_fill_1 FILLER_41_94 ();
 sg13g2_decap_8 FILLER_41_99 ();
 sg13g2_decap_8 FILLER_41_106 ();
 sg13g2_decap_8 FILLER_41_113 ();
 sg13g2_fill_1 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_4 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_185 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_fill_1 FILLER_41_233 ();
 sg13g2_fill_2 FILLER_41_251 ();
 sg13g2_fill_2 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_298 ();
 sg13g2_decap_4 FILLER_41_305 ();
 sg13g2_fill_2 FILLER_41_309 ();
 sg13g2_decap_4 FILLER_41_373 ();
 sg13g2_fill_1 FILLER_41_377 ();
 sg13g2_fill_2 FILLER_41_383 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_decap_8 FILLER_41_472 ();
 sg13g2_decap_4 FILLER_41_483 ();
 sg13g2_fill_2 FILLER_41_487 ();
 sg13g2_decap_8 FILLER_41_493 ();
 sg13g2_decap_4 FILLER_41_500 ();
 sg13g2_fill_2 FILLER_41_504 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_fill_1 FILLER_41_585 ();
 sg13g2_decap_8 FILLER_41_605 ();
 sg13g2_decap_4 FILLER_41_612 ();
 sg13g2_fill_2 FILLER_41_616 ();
 sg13g2_decap_4 FILLER_41_622 ();
 sg13g2_fill_2 FILLER_41_635 ();
 sg13g2_decap_8 FILLER_41_642 ();
 sg13g2_decap_4 FILLER_41_649 ();
 sg13g2_fill_2 FILLER_41_653 ();
 sg13g2_decap_8 FILLER_41_661 ();
 sg13g2_decap_4 FILLER_41_668 ();
 sg13g2_fill_1 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_fill_2 FILLER_41_696 ();
 sg13g2_fill_1 FILLER_41_698 ();
 sg13g2_fill_1 FILLER_41_706 ();
 sg13g2_decap_8 FILLER_41_753 ();
 sg13g2_decap_4 FILLER_41_760 ();
 sg13g2_fill_1 FILLER_41_764 ();
 sg13g2_decap_4 FILLER_41_768 ();
 sg13g2_fill_2 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_790 ();
 sg13g2_fill_1 FILLER_41_797 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_fill_2 FILLER_41_821 ();
 sg13g2_fill_1 FILLER_41_823 ();
 sg13g2_fill_2 FILLER_41_852 ();
 sg13g2_decap_8 FILLER_41_867 ();
 sg13g2_fill_2 FILLER_41_874 ();
 sg13g2_fill_2 FILLER_41_1006 ();
 sg13g2_fill_1 FILLER_41_1036 ();
 sg13g2_fill_2 FILLER_41_1050 ();
 sg13g2_fill_1 FILLER_41_1073 ();
 sg13g2_decap_8 FILLER_41_1087 ();
 sg13g2_decap_8 FILLER_41_1094 ();
 sg13g2_decap_4 FILLER_41_1101 ();
 sg13g2_fill_2 FILLER_41_1105 ();
 sg13g2_fill_1 FILLER_41_1146 ();
 sg13g2_fill_1 FILLER_41_1165 ();
 sg13g2_fill_1 FILLER_41_1176 ();
 sg13g2_fill_1 FILLER_41_1193 ();
 sg13g2_decap_4 FILLER_41_1224 ();
 sg13g2_fill_1 FILLER_41_1238 ();
 sg13g2_decap_4 FILLER_41_1263 ();
 sg13g2_fill_2 FILLER_41_1267 ();
 sg13g2_fill_2 FILLER_41_1279 ();
 sg13g2_fill_2 FILLER_41_1293 ();
 sg13g2_fill_2 FILLER_41_1305 ();
 sg13g2_fill_2 FILLER_41_1316 ();
 sg13g2_fill_1 FILLER_41_1367 ();
 sg13g2_fill_2 FILLER_41_1377 ();
 sg13g2_fill_1 FILLER_41_1449 ();
 sg13g2_fill_2 FILLER_41_1461 ();
 sg13g2_fill_2 FILLER_41_1489 ();
 sg13g2_decap_4 FILLER_41_1538 ();
 sg13g2_fill_2 FILLER_41_1549 ();
 sg13g2_fill_2 FILLER_41_1585 ();
 sg13g2_fill_1 FILLER_41_1587 ();
 sg13g2_fill_2 FILLER_41_1675 ();
 sg13g2_fill_2 FILLER_41_1713 ();
 sg13g2_fill_2 FILLER_41_1731 ();
 sg13g2_fill_1 FILLER_41_1733 ();
 sg13g2_decap_4 FILLER_41_1812 ();
 sg13g2_fill_1 FILLER_41_1816 ();
 sg13g2_decap_8 FILLER_41_1826 ();
 sg13g2_decap_4 FILLER_41_1833 ();
 sg13g2_fill_2 FILLER_41_1870 ();
 sg13g2_decap_4 FILLER_41_1900 ();
 sg13g2_fill_2 FILLER_41_1917 ();
 sg13g2_decap_4 FILLER_41_1927 ();
 sg13g2_fill_1 FILLER_41_1939 ();
 sg13g2_decap_4 FILLER_41_1954 ();
 sg13g2_fill_2 FILLER_41_1958 ();
 sg13g2_fill_1 FILLER_41_2036 ();
 sg13g2_fill_2 FILLER_41_2048 ();
 sg13g2_fill_1 FILLER_41_2062 ();
 sg13g2_fill_2 FILLER_41_2068 ();
 sg13g2_fill_1 FILLER_41_2090 ();
 sg13g2_decap_8 FILLER_41_2133 ();
 sg13g2_fill_2 FILLER_41_2140 ();
 sg13g2_fill_1 FILLER_41_2142 ();
 sg13g2_fill_1 FILLER_41_2170 ();
 sg13g2_fill_1 FILLER_41_2180 ();
 sg13g2_fill_2 FILLER_41_2190 ();
 sg13g2_fill_2 FILLER_41_2205 ();
 sg13g2_fill_2 FILLER_41_2216 ();
 sg13g2_fill_1 FILLER_41_2230 ();
 sg13g2_fill_2 FILLER_41_2262 ();
 sg13g2_fill_2 FILLER_41_2295 ();
 sg13g2_decap_8 FILLER_41_2313 ();
 sg13g2_decap_4 FILLER_41_2320 ();
 sg13g2_fill_2 FILLER_41_2328 ();
 sg13g2_fill_1 FILLER_41_2330 ();
 sg13g2_fill_2 FILLER_41_2364 ();
 sg13g2_fill_1 FILLER_41_2407 ();
 sg13g2_decap_8 FILLER_41_2430 ();
 sg13g2_decap_8 FILLER_41_2437 ();
 sg13g2_decap_8 FILLER_41_2444 ();
 sg13g2_decap_8 FILLER_41_2451 ();
 sg13g2_decap_8 FILLER_41_2458 ();
 sg13g2_decap_8 FILLER_41_2465 ();
 sg13g2_decap_8 FILLER_41_2472 ();
 sg13g2_decap_8 FILLER_41_2479 ();
 sg13g2_decap_8 FILLER_41_2486 ();
 sg13g2_decap_8 FILLER_41_2493 ();
 sg13g2_decap_8 FILLER_41_2500 ();
 sg13g2_decap_8 FILLER_41_2507 ();
 sg13g2_decap_8 FILLER_41_2514 ();
 sg13g2_decap_8 FILLER_41_2521 ();
 sg13g2_decap_8 FILLER_41_2528 ();
 sg13g2_decap_8 FILLER_41_2535 ();
 sg13g2_decap_8 FILLER_41_2542 ();
 sg13g2_decap_8 FILLER_41_2549 ();
 sg13g2_decap_8 FILLER_41_2556 ();
 sg13g2_decap_8 FILLER_41_2563 ();
 sg13g2_decap_8 FILLER_41_2570 ();
 sg13g2_decap_8 FILLER_41_2577 ();
 sg13g2_decap_8 FILLER_41_2584 ();
 sg13g2_decap_8 FILLER_41_2591 ();
 sg13g2_decap_8 FILLER_41_2598 ();
 sg13g2_decap_8 FILLER_41_2605 ();
 sg13g2_decap_8 FILLER_41_2612 ();
 sg13g2_decap_8 FILLER_41_2619 ();
 sg13g2_decap_8 FILLER_41_2626 ();
 sg13g2_decap_8 FILLER_41_2633 ();
 sg13g2_decap_8 FILLER_41_2640 ();
 sg13g2_decap_8 FILLER_41_2647 ();
 sg13g2_decap_8 FILLER_41_2654 ();
 sg13g2_decap_8 FILLER_41_2661 ();
 sg13g2_decap_4 FILLER_41_2668 ();
 sg13g2_fill_2 FILLER_41_2672 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_decap_8 FILLER_42_30 ();
 sg13g2_decap_4 FILLER_42_37 ();
 sg13g2_fill_2 FILLER_42_112 ();
 sg13g2_decap_4 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_fill_1 FILLER_42_201 ();
 sg13g2_fill_2 FILLER_42_223 ();
 sg13g2_fill_2 FILLER_42_278 ();
 sg13g2_fill_2 FILLER_42_293 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_fill_2 FILLER_42_368 ();
 sg13g2_fill_1 FILLER_42_397 ();
 sg13g2_fill_2 FILLER_42_489 ();
 sg13g2_decap_8 FILLER_42_500 ();
 sg13g2_fill_2 FILLER_42_507 ();
 sg13g2_fill_2 FILLER_42_568 ();
 sg13g2_decap_4 FILLER_42_616 ();
 sg13g2_fill_2 FILLER_42_620 ();
 sg13g2_fill_2 FILLER_42_629 ();
 sg13g2_fill_2 FILLER_42_655 ();
 sg13g2_fill_2 FILLER_42_675 ();
 sg13g2_fill_1 FILLER_42_677 ();
 sg13g2_decap_8 FILLER_42_684 ();
 sg13g2_decap_8 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_698 ();
 sg13g2_decap_8 FILLER_42_705 ();
 sg13g2_fill_1 FILLER_42_712 ();
 sg13g2_decap_8 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_fill_2 FILLER_42_810 ();
 sg13g2_fill_1 FILLER_42_825 ();
 sg13g2_decap_4 FILLER_42_869 ();
 sg13g2_fill_1 FILLER_42_917 ();
 sg13g2_fill_2 FILLER_42_927 ();
 sg13g2_fill_1 FILLER_42_929 ();
 sg13g2_fill_1 FILLER_42_967 ();
 sg13g2_fill_2 FILLER_42_1029 ();
 sg13g2_fill_1 FILLER_42_1031 ();
 sg13g2_fill_1 FILLER_42_1075 ();
 sg13g2_decap_8 FILLER_42_1085 ();
 sg13g2_decap_4 FILLER_42_1092 ();
 sg13g2_fill_2 FILLER_42_1096 ();
 sg13g2_fill_2 FILLER_42_1136 ();
 sg13g2_decap_4 FILLER_42_1179 ();
 sg13g2_fill_1 FILLER_42_1183 ();
 sg13g2_fill_2 FILLER_42_1205 ();
 sg13g2_decap_8 FILLER_42_1234 ();
 sg13g2_decap_4 FILLER_42_1241 ();
 sg13g2_fill_1 FILLER_42_1272 ();
 sg13g2_fill_1 FILLER_42_1304 ();
 sg13g2_fill_1 FILLER_42_1309 ();
 sg13g2_fill_1 FILLER_42_1325 ();
 sg13g2_fill_2 FILLER_42_1330 ();
 sg13g2_fill_2 FILLER_42_1338 ();
 sg13g2_fill_2 FILLER_42_1421 ();
 sg13g2_fill_2 FILLER_42_1446 ();
 sg13g2_decap_8 FILLER_42_1453 ();
 sg13g2_decap_8 FILLER_42_1460 ();
 sg13g2_fill_2 FILLER_42_1473 ();
 sg13g2_fill_2 FILLER_42_1498 ();
 sg13g2_decap_4 FILLER_42_1521 ();
 sg13g2_decap_8 FILLER_42_1532 ();
 sg13g2_decap_8 FILLER_42_1539 ();
 sg13g2_fill_1 FILLER_42_1546 ();
 sg13g2_fill_2 FILLER_42_1565 ();
 sg13g2_decap_4 FILLER_42_1580 ();
 sg13g2_fill_1 FILLER_42_1584 ();
 sg13g2_fill_2 FILLER_42_1675 ();
 sg13g2_fill_1 FILLER_42_1677 ();
 sg13g2_fill_1 FILLER_42_1687 ();
 sg13g2_fill_1 FILLER_42_1697 ();
 sg13g2_fill_2 FILLER_42_1711 ();
 sg13g2_fill_1 FILLER_42_1721 ();
 sg13g2_fill_2 FILLER_42_1738 ();
 sg13g2_fill_1 FILLER_42_1740 ();
 sg13g2_fill_1 FILLER_42_1754 ();
 sg13g2_fill_2 FILLER_42_1786 ();
 sg13g2_decap_8 FILLER_42_1804 ();
 sg13g2_fill_1 FILLER_42_1811 ();
 sg13g2_fill_2 FILLER_42_1816 ();
 sg13g2_decap_8 FILLER_42_1831 ();
 sg13g2_fill_1 FILLER_42_1838 ();
 sg13g2_fill_2 FILLER_42_1857 ();
 sg13g2_fill_1 FILLER_42_1871 ();
 sg13g2_decap_4 FILLER_42_1915 ();
 sg13g2_decap_4 FILLER_42_1927 ();
 sg13g2_fill_1 FILLER_42_1954 ();
 sg13g2_fill_1 FILLER_42_1992 ();
 sg13g2_fill_2 FILLER_42_2005 ();
 sg13g2_fill_1 FILLER_42_2030 ();
 sg13g2_decap_8 FILLER_42_2040 ();
 sg13g2_fill_2 FILLER_42_2061 ();
 sg13g2_fill_2 FILLER_42_2078 ();
 sg13g2_fill_1 FILLER_42_2080 ();
 sg13g2_decap_4 FILLER_42_2084 ();
 sg13g2_fill_2 FILLER_42_2088 ();
 sg13g2_fill_1 FILLER_42_2105 ();
 sg13g2_decap_8 FILLER_42_2124 ();
 sg13g2_decap_4 FILLER_42_2131 ();
 sg13g2_fill_1 FILLER_42_2135 ();
 sg13g2_decap_4 FILLER_42_2154 ();
 sg13g2_fill_1 FILLER_42_2158 ();
 sg13g2_fill_2 FILLER_42_2208 ();
 sg13g2_fill_1 FILLER_42_2318 ();
 sg13g2_fill_2 FILLER_42_2368 ();
 sg13g2_fill_1 FILLER_42_2397 ();
 sg13g2_decap_8 FILLER_42_2435 ();
 sg13g2_decap_8 FILLER_42_2442 ();
 sg13g2_decap_8 FILLER_42_2449 ();
 sg13g2_decap_8 FILLER_42_2456 ();
 sg13g2_decap_8 FILLER_42_2463 ();
 sg13g2_decap_8 FILLER_42_2470 ();
 sg13g2_decap_8 FILLER_42_2477 ();
 sg13g2_decap_8 FILLER_42_2484 ();
 sg13g2_decap_8 FILLER_42_2491 ();
 sg13g2_decap_8 FILLER_42_2498 ();
 sg13g2_decap_8 FILLER_42_2505 ();
 sg13g2_decap_8 FILLER_42_2512 ();
 sg13g2_decap_8 FILLER_42_2519 ();
 sg13g2_decap_8 FILLER_42_2526 ();
 sg13g2_decap_8 FILLER_42_2533 ();
 sg13g2_decap_8 FILLER_42_2540 ();
 sg13g2_decap_8 FILLER_42_2547 ();
 sg13g2_decap_8 FILLER_42_2554 ();
 sg13g2_decap_8 FILLER_42_2561 ();
 sg13g2_decap_8 FILLER_42_2568 ();
 sg13g2_decap_8 FILLER_42_2575 ();
 sg13g2_decap_8 FILLER_42_2582 ();
 sg13g2_decap_8 FILLER_42_2589 ();
 sg13g2_decap_8 FILLER_42_2596 ();
 sg13g2_decap_8 FILLER_42_2603 ();
 sg13g2_decap_8 FILLER_42_2610 ();
 sg13g2_decap_8 FILLER_42_2617 ();
 sg13g2_decap_8 FILLER_42_2624 ();
 sg13g2_decap_8 FILLER_42_2631 ();
 sg13g2_decap_8 FILLER_42_2638 ();
 sg13g2_decap_8 FILLER_42_2645 ();
 sg13g2_decap_8 FILLER_42_2652 ();
 sg13g2_decap_8 FILLER_42_2659 ();
 sg13g2_decap_8 FILLER_42_2666 ();
 sg13g2_fill_1 FILLER_42_2673 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_33 ();
 sg13g2_fill_1 FILLER_43_106 ();
 sg13g2_fill_1 FILLER_43_139 ();
 sg13g2_decap_4 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_197 ();
 sg13g2_decap_4 FILLER_43_212 ();
 sg13g2_decap_8 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_227 ();
 sg13g2_decap_4 FILLER_43_284 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_360 ();
 sg13g2_fill_2 FILLER_43_415 ();
 sg13g2_fill_1 FILLER_43_417 ();
 sg13g2_fill_1 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_fill_1 FILLER_43_516 ();
 sg13g2_decap_4 FILLER_43_522 ();
 sg13g2_fill_2 FILLER_43_535 ();
 sg13g2_fill_2 FILLER_43_560 ();
 sg13g2_fill_2 FILLER_43_580 ();
 sg13g2_fill_1 FILLER_43_648 ();
 sg13g2_decap_8 FILLER_43_689 ();
 sg13g2_decap_4 FILLER_43_696 ();
 sg13g2_fill_1 FILLER_43_700 ();
 sg13g2_decap_4 FILLER_43_748 ();
 sg13g2_fill_2 FILLER_43_759 ();
 sg13g2_decap_8 FILLER_43_816 ();
 sg13g2_fill_2 FILLER_43_823 ();
 sg13g2_fill_2 FILLER_43_843 ();
 sg13g2_fill_1 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_860 ();
 sg13g2_fill_2 FILLER_43_867 ();
 sg13g2_fill_1 FILLER_43_897 ();
 sg13g2_fill_2 FILLER_43_959 ();
 sg13g2_decap_4 FILLER_43_1021 ();
 sg13g2_fill_2 FILLER_43_1030 ();
 sg13g2_fill_1 FILLER_43_1032 ();
 sg13g2_decap_4 FILLER_43_1037 ();
 sg13g2_decap_8 FILLER_43_1079 ();
 sg13g2_fill_1 FILLER_43_1086 ();
 sg13g2_decap_4 FILLER_43_1095 ();
 sg13g2_fill_2 FILLER_43_1099 ();
 sg13g2_fill_2 FILLER_43_1127 ();
 sg13g2_fill_1 FILLER_43_1133 ();
 sg13g2_decap_8 FILLER_43_1149 ();
 sg13g2_fill_2 FILLER_43_1156 ();
 sg13g2_fill_1 FILLER_43_1158 ();
 sg13g2_fill_2 FILLER_43_1308 ();
 sg13g2_fill_1 FILLER_43_1310 ();
 sg13g2_decap_8 FILLER_43_1333 ();
 sg13g2_fill_1 FILLER_43_1367 ();
 sg13g2_decap_4 FILLER_43_1452 ();
 sg13g2_fill_1 FILLER_43_1459 ();
 sg13g2_fill_2 FILLER_43_1475 ();
 sg13g2_fill_1 FILLER_43_1477 ();
 sg13g2_fill_1 FILLER_43_1483 ();
 sg13g2_fill_1 FILLER_43_1493 ();
 sg13g2_fill_1 FILLER_43_1542 ();
 sg13g2_fill_2 FILLER_43_1592 ();
 sg13g2_fill_1 FILLER_43_1594 ();
 sg13g2_fill_2 FILLER_43_1686 ();
 sg13g2_fill_2 FILLER_43_1715 ();
 sg13g2_fill_1 FILLER_43_1717 ();
 sg13g2_fill_2 FILLER_43_1746 ();
 sg13g2_fill_2 FILLER_43_1784 ();
 sg13g2_decap_4 FILLER_43_1804 ();
 sg13g2_fill_2 FILLER_43_1813 ();
 sg13g2_fill_1 FILLER_43_1842 ();
 sg13g2_decap_4 FILLER_43_1913 ();
 sg13g2_fill_1 FILLER_43_1917 ();
 sg13g2_decap_4 FILLER_43_1944 ();
 sg13g2_fill_1 FILLER_43_1957 ();
 sg13g2_decap_8 FILLER_43_1986 ();
 sg13g2_fill_2 FILLER_43_1993 ();
 sg13g2_fill_1 FILLER_43_1995 ();
 sg13g2_fill_2 FILLER_43_2026 ();
 sg13g2_fill_2 FILLER_43_2035 ();
 sg13g2_fill_1 FILLER_43_2041 ();
 sg13g2_fill_1 FILLER_43_2060 ();
 sg13g2_decap_4 FILLER_43_2084 ();
 sg13g2_fill_1 FILLER_43_2088 ();
 sg13g2_decap_8 FILLER_43_2121 ();
 sg13g2_fill_2 FILLER_43_2137 ();
 sg13g2_fill_1 FILLER_43_2139 ();
 sg13g2_decap_8 FILLER_43_2157 ();
 sg13g2_fill_2 FILLER_43_2164 ();
 sg13g2_fill_1 FILLER_43_2166 ();
 sg13g2_fill_2 FILLER_43_2199 ();
 sg13g2_fill_2 FILLER_43_2229 ();
 sg13g2_fill_1 FILLER_43_2231 ();
 sg13g2_fill_1 FILLER_43_2274 ();
 sg13g2_fill_1 FILLER_43_2333 ();
 sg13g2_fill_1 FILLER_43_2366 ();
 sg13g2_fill_1 FILLER_43_2386 ();
 sg13g2_decap_8 FILLER_43_2427 ();
 sg13g2_decap_8 FILLER_43_2434 ();
 sg13g2_decap_8 FILLER_43_2441 ();
 sg13g2_decap_8 FILLER_43_2448 ();
 sg13g2_decap_8 FILLER_43_2455 ();
 sg13g2_decap_8 FILLER_43_2462 ();
 sg13g2_decap_8 FILLER_43_2469 ();
 sg13g2_decap_8 FILLER_43_2476 ();
 sg13g2_decap_8 FILLER_43_2483 ();
 sg13g2_decap_8 FILLER_43_2490 ();
 sg13g2_decap_8 FILLER_43_2497 ();
 sg13g2_decap_8 FILLER_43_2504 ();
 sg13g2_decap_8 FILLER_43_2511 ();
 sg13g2_decap_8 FILLER_43_2518 ();
 sg13g2_decap_8 FILLER_43_2525 ();
 sg13g2_decap_8 FILLER_43_2532 ();
 sg13g2_decap_8 FILLER_43_2539 ();
 sg13g2_decap_8 FILLER_43_2546 ();
 sg13g2_decap_8 FILLER_43_2553 ();
 sg13g2_decap_8 FILLER_43_2560 ();
 sg13g2_decap_8 FILLER_43_2567 ();
 sg13g2_decap_8 FILLER_43_2574 ();
 sg13g2_decap_8 FILLER_43_2581 ();
 sg13g2_decap_8 FILLER_43_2588 ();
 sg13g2_decap_8 FILLER_43_2595 ();
 sg13g2_decap_8 FILLER_43_2602 ();
 sg13g2_decap_8 FILLER_43_2609 ();
 sg13g2_decap_8 FILLER_43_2616 ();
 sg13g2_decap_8 FILLER_43_2623 ();
 sg13g2_decap_8 FILLER_43_2630 ();
 sg13g2_decap_8 FILLER_43_2637 ();
 sg13g2_decap_8 FILLER_43_2644 ();
 sg13g2_decap_8 FILLER_43_2651 ();
 sg13g2_decap_8 FILLER_43_2658 ();
 sg13g2_decap_8 FILLER_43_2665 ();
 sg13g2_fill_2 FILLER_43_2672 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_97 ();
 sg13g2_fill_1 FILLER_44_99 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_143 ();
 sg13g2_fill_1 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_decap_4 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_282 ();
 sg13g2_fill_2 FILLER_44_305 ();
 sg13g2_fill_1 FILLER_44_370 ();
 sg13g2_fill_2 FILLER_44_403 ();
 sg13g2_fill_1 FILLER_44_405 ();
 sg13g2_fill_1 FILLER_44_438 ();
 sg13g2_fill_1 FILLER_44_450 ();
 sg13g2_decap_4 FILLER_44_510 ();
 sg13g2_decap_8 FILLER_44_527 ();
 sg13g2_decap_4 FILLER_44_534 ();
 sg13g2_fill_2 FILLER_44_538 ();
 sg13g2_fill_2 FILLER_44_592 ();
 sg13g2_decap_4 FILLER_44_613 ();
 sg13g2_decap_4 FILLER_44_686 ();
 sg13g2_fill_1 FILLER_44_729 ();
 sg13g2_fill_2 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_818 ();
 sg13g2_decap_4 FILLER_44_825 ();
 sg13g2_fill_2 FILLER_44_829 ();
 sg13g2_fill_2 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_4 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_858 ();
 sg13g2_fill_1 FILLER_44_872 ();
 sg13g2_fill_1 FILLER_44_901 ();
 sg13g2_fill_1 FILLER_44_984 ();
 sg13g2_fill_2 FILLER_44_1040 ();
 sg13g2_fill_2 FILLER_44_1050 ();
 sg13g2_fill_1 FILLER_44_1052 ();
 sg13g2_decap_8 FILLER_44_1067 ();
 sg13g2_fill_1 FILLER_44_1074 ();
 sg13g2_decap_8 FILLER_44_1096 ();
 sg13g2_decap_4 FILLER_44_1103 ();
 sg13g2_fill_1 FILLER_44_1107 ();
 sg13g2_fill_1 FILLER_44_1121 ();
 sg13g2_decap_4 FILLER_44_1139 ();
 sg13g2_fill_1 FILLER_44_1143 ();
 sg13g2_fill_2 FILLER_44_1154 ();
 sg13g2_fill_1 FILLER_44_1191 ();
 sg13g2_fill_2 FILLER_44_1284 ();
 sg13g2_fill_2 FILLER_44_1314 ();
 sg13g2_fill_1 FILLER_44_1347 ();
 sg13g2_decap_4 FILLER_44_1354 ();
 sg13g2_decap_4 FILLER_44_1364 ();
 sg13g2_fill_1 FILLER_44_1396 ();
 sg13g2_decap_4 FILLER_44_1409 ();
 sg13g2_fill_1 FILLER_44_1413 ();
 sg13g2_fill_2 FILLER_44_1454 ();
 sg13g2_fill_2 FILLER_44_1479 ();
 sg13g2_fill_1 FILLER_44_1481 ();
 sg13g2_decap_4 FILLER_44_1509 ();
 sg13g2_fill_2 FILLER_44_1513 ();
 sg13g2_fill_1 FILLER_44_1543 ();
 sg13g2_fill_2 FILLER_44_1554 ();
 sg13g2_fill_2 FILLER_44_1605 ();
 sg13g2_fill_1 FILLER_44_1654 ();
 sg13g2_fill_2 FILLER_44_1682 ();
 sg13g2_fill_1 FILLER_44_1684 ();
 sg13g2_decap_8 FILLER_44_1783 ();
 sg13g2_decap_4 FILLER_44_1790 ();
 sg13g2_fill_2 FILLER_44_1799 ();
 sg13g2_fill_1 FILLER_44_1823 ();
 sg13g2_fill_1 FILLER_44_1848 ();
 sg13g2_fill_1 FILLER_44_1862 ();
 sg13g2_fill_2 FILLER_44_1918 ();
 sg13g2_fill_2 FILLER_44_1970 ();
 sg13g2_decap_8 FILLER_44_1981 ();
 sg13g2_fill_2 FILLER_44_1992 ();
 sg13g2_fill_2 FILLER_44_2021 ();
 sg13g2_fill_1 FILLER_44_2023 ();
 sg13g2_fill_1 FILLER_44_2037 ();
 sg13g2_fill_2 FILLER_44_2050 ();
 sg13g2_fill_1 FILLER_44_2062 ();
 sg13g2_fill_2 FILLER_44_2069 ();
 sg13g2_fill_1 FILLER_44_2081 ();
 sg13g2_fill_2 FILLER_44_2142 ();
 sg13g2_fill_1 FILLER_44_2150 ();
 sg13g2_fill_1 FILLER_44_2164 ();
 sg13g2_fill_2 FILLER_44_2232 ();
 sg13g2_fill_1 FILLER_44_2234 ();
 sg13g2_fill_2 FILLER_44_2272 ();
 sg13g2_fill_2 FILLER_44_2297 ();
 sg13g2_decap_4 FILLER_44_2326 ();
 sg13g2_decap_8 FILLER_44_2424 ();
 sg13g2_decap_8 FILLER_44_2431 ();
 sg13g2_decap_8 FILLER_44_2438 ();
 sg13g2_decap_8 FILLER_44_2445 ();
 sg13g2_decap_8 FILLER_44_2452 ();
 sg13g2_decap_8 FILLER_44_2459 ();
 sg13g2_decap_8 FILLER_44_2466 ();
 sg13g2_decap_8 FILLER_44_2473 ();
 sg13g2_decap_8 FILLER_44_2480 ();
 sg13g2_decap_8 FILLER_44_2487 ();
 sg13g2_decap_8 FILLER_44_2494 ();
 sg13g2_decap_8 FILLER_44_2501 ();
 sg13g2_decap_8 FILLER_44_2508 ();
 sg13g2_decap_8 FILLER_44_2515 ();
 sg13g2_decap_8 FILLER_44_2522 ();
 sg13g2_decap_8 FILLER_44_2529 ();
 sg13g2_decap_8 FILLER_44_2536 ();
 sg13g2_decap_8 FILLER_44_2543 ();
 sg13g2_decap_8 FILLER_44_2550 ();
 sg13g2_decap_8 FILLER_44_2557 ();
 sg13g2_decap_8 FILLER_44_2564 ();
 sg13g2_decap_8 FILLER_44_2571 ();
 sg13g2_decap_8 FILLER_44_2578 ();
 sg13g2_decap_8 FILLER_44_2585 ();
 sg13g2_decap_8 FILLER_44_2592 ();
 sg13g2_decap_8 FILLER_44_2599 ();
 sg13g2_decap_8 FILLER_44_2606 ();
 sg13g2_decap_8 FILLER_44_2613 ();
 sg13g2_decap_8 FILLER_44_2620 ();
 sg13g2_decap_8 FILLER_44_2627 ();
 sg13g2_decap_8 FILLER_44_2634 ();
 sg13g2_decap_8 FILLER_44_2641 ();
 sg13g2_decap_8 FILLER_44_2648 ();
 sg13g2_decap_8 FILLER_44_2655 ();
 sg13g2_decap_8 FILLER_44_2662 ();
 sg13g2_decap_4 FILLER_44_2669 ();
 sg13g2_fill_1 FILLER_44_2673 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_68 ();
 sg13g2_fill_1 FILLER_45_70 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_decap_4 FILLER_45_102 ();
 sg13g2_decap_8 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_222 ();
 sg13g2_fill_2 FILLER_45_229 ();
 sg13g2_fill_1 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_256 ();
 sg13g2_fill_2 FILLER_45_263 ();
 sg13g2_fill_1 FILLER_45_265 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_fill_1 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_328 ();
 sg13g2_fill_1 FILLER_45_338 ();
 sg13g2_fill_1 FILLER_45_353 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_fill_2 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_380 ();
 sg13g2_fill_1 FILLER_45_410 ();
 sg13g2_fill_2 FILLER_45_426 ();
 sg13g2_fill_2 FILLER_45_447 ();
 sg13g2_fill_1 FILLER_45_449 ();
 sg13g2_fill_2 FILLER_45_475 ();
 sg13g2_fill_1 FILLER_45_477 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_fill_2 FILLER_45_497 ();
 sg13g2_fill_1 FILLER_45_499 ();
 sg13g2_fill_1 FILLER_45_527 ();
 sg13g2_fill_2 FILLER_45_537 ();
 sg13g2_fill_2 FILLER_45_566 ();
 sg13g2_fill_1 FILLER_45_586 ();
 sg13g2_decap_4 FILLER_45_600 ();
 sg13g2_fill_2 FILLER_45_604 ();
 sg13g2_fill_1 FILLER_45_622 ();
 sg13g2_decap_4 FILLER_45_632 ();
 sg13g2_decap_4 FILLER_45_650 ();
 sg13g2_fill_2 FILLER_45_654 ();
 sg13g2_fill_1 FILLER_45_689 ();
 sg13g2_fill_1 FILLER_45_721 ();
 sg13g2_decap_4 FILLER_45_746 ();
 sg13g2_fill_2 FILLER_45_750 ();
 sg13g2_decap_4 FILLER_45_796 ();
 sg13g2_decap_4 FILLER_45_809 ();
 sg13g2_decap_4 FILLER_45_826 ();
 sg13g2_fill_1 FILLER_45_830 ();
 sg13g2_fill_2 FILLER_45_867 ();
 sg13g2_fill_1 FILLER_45_869 ();
 sg13g2_fill_2 FILLER_45_902 ();
 sg13g2_fill_2 FILLER_45_948 ();
 sg13g2_fill_2 FILLER_45_959 ();
 sg13g2_fill_1 FILLER_45_974 ();
 sg13g2_fill_1 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1032 ();
 sg13g2_fill_1 FILLER_45_1042 ();
 sg13g2_decap_8 FILLER_45_1053 ();
 sg13g2_decap_8 FILLER_45_1060 ();
 sg13g2_decap_8 FILLER_45_1067 ();
 sg13g2_fill_1 FILLER_45_1074 ();
 sg13g2_fill_2 FILLER_45_1097 ();
 sg13g2_fill_2 FILLER_45_1104 ();
 sg13g2_fill_1 FILLER_45_1106 ();
 sg13g2_fill_2 FILLER_45_1121 ();
 sg13g2_fill_1 FILLER_45_1129 ();
 sg13g2_fill_1 FILLER_45_1204 ();
 sg13g2_fill_1 FILLER_45_1268 ();
 sg13g2_fill_2 FILLER_45_1294 ();
 sg13g2_fill_1 FILLER_45_1296 ();
 sg13g2_fill_1 FILLER_45_1329 ();
 sg13g2_decap_8 FILLER_45_1335 ();
 sg13g2_fill_2 FILLER_45_1342 ();
 sg13g2_fill_1 FILLER_45_1400 ();
 sg13g2_fill_2 FILLER_45_1406 ();
 sg13g2_decap_4 FILLER_45_1421 ();
 sg13g2_fill_1 FILLER_45_1425 ();
 sg13g2_fill_2 FILLER_45_1466 ();
 sg13g2_fill_2 FILLER_45_1504 ();
 sg13g2_fill_2 FILLER_45_1521 ();
 sg13g2_fill_2 FILLER_45_1608 ();
 sg13g2_fill_1 FILLER_45_1615 ();
 sg13g2_fill_2 FILLER_45_1652 ();
 sg13g2_fill_1 FILLER_45_1707 ();
 sg13g2_decap_4 FILLER_45_1748 ();
 sg13g2_decap_8 FILLER_45_1779 ();
 sg13g2_fill_1 FILLER_45_1786 ();
 sg13g2_fill_1 FILLER_45_1815 ();
 sg13g2_fill_2 FILLER_45_1883 ();
 sg13g2_fill_1 FILLER_45_1907 ();
 sg13g2_fill_1 FILLER_45_1925 ();
 sg13g2_decap_8 FILLER_45_1974 ();
 sg13g2_fill_1 FILLER_45_1981 ();
 sg13g2_fill_2 FILLER_45_1991 ();
 sg13g2_fill_2 FILLER_45_2039 ();
 sg13g2_fill_1 FILLER_45_2041 ();
 sg13g2_fill_2 FILLER_45_2047 ();
 sg13g2_decap_4 FILLER_45_2054 ();
 sg13g2_fill_2 FILLER_45_2062 ();
 sg13g2_fill_1 FILLER_45_2064 ();
 sg13g2_fill_2 FILLER_45_2074 ();
 sg13g2_fill_1 FILLER_45_2076 ();
 sg13g2_decap_8 FILLER_45_2114 ();
 sg13g2_decap_4 FILLER_45_2121 ();
 sg13g2_decap_4 FILLER_45_2179 ();
 sg13g2_fill_2 FILLER_45_2272 ();
 sg13g2_fill_2 FILLER_45_2310 ();
 sg13g2_decap_8 FILLER_45_2325 ();
 sg13g2_decap_4 FILLER_45_2332 ();
 sg13g2_decap_8 FILLER_45_2418 ();
 sg13g2_decap_8 FILLER_45_2425 ();
 sg13g2_decap_8 FILLER_45_2432 ();
 sg13g2_decap_8 FILLER_45_2439 ();
 sg13g2_decap_8 FILLER_45_2446 ();
 sg13g2_decap_8 FILLER_45_2453 ();
 sg13g2_decap_8 FILLER_45_2460 ();
 sg13g2_decap_8 FILLER_45_2467 ();
 sg13g2_decap_8 FILLER_45_2474 ();
 sg13g2_decap_8 FILLER_45_2481 ();
 sg13g2_decap_8 FILLER_45_2488 ();
 sg13g2_decap_8 FILLER_45_2495 ();
 sg13g2_decap_8 FILLER_45_2502 ();
 sg13g2_decap_8 FILLER_45_2509 ();
 sg13g2_decap_8 FILLER_45_2516 ();
 sg13g2_decap_8 FILLER_45_2523 ();
 sg13g2_decap_8 FILLER_45_2530 ();
 sg13g2_decap_8 FILLER_45_2537 ();
 sg13g2_decap_8 FILLER_45_2544 ();
 sg13g2_decap_8 FILLER_45_2551 ();
 sg13g2_decap_8 FILLER_45_2558 ();
 sg13g2_decap_8 FILLER_45_2565 ();
 sg13g2_decap_8 FILLER_45_2572 ();
 sg13g2_decap_8 FILLER_45_2579 ();
 sg13g2_decap_8 FILLER_45_2586 ();
 sg13g2_decap_8 FILLER_45_2593 ();
 sg13g2_decap_8 FILLER_45_2600 ();
 sg13g2_decap_8 FILLER_45_2607 ();
 sg13g2_decap_8 FILLER_45_2614 ();
 sg13g2_decap_8 FILLER_45_2621 ();
 sg13g2_decap_8 FILLER_45_2628 ();
 sg13g2_decap_8 FILLER_45_2635 ();
 sg13g2_decap_8 FILLER_45_2642 ();
 sg13g2_decap_8 FILLER_45_2649 ();
 sg13g2_decap_8 FILLER_45_2656 ();
 sg13g2_decap_8 FILLER_45_2663 ();
 sg13g2_decap_4 FILLER_45_2670 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_23 ();
 sg13g2_fill_2 FILLER_46_52 ();
 sg13g2_fill_1 FILLER_46_54 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_fill_2 FILLER_46_105 ();
 sg13g2_fill_1 FILLER_46_107 ();
 sg13g2_fill_1 FILLER_46_122 ();
 sg13g2_decap_8 FILLER_46_207 ();
 sg13g2_fill_2 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_340 ();
 sg13g2_fill_1 FILLER_46_382 ();
 sg13g2_fill_2 FILLER_46_411 ();
 sg13g2_decap_8 FILLER_46_429 ();
 sg13g2_decap_4 FILLER_46_436 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_fill_2 FILLER_46_490 ();
 sg13g2_fill_1 FILLER_46_492 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_fill_2 FILLER_46_658 ();
 sg13g2_fill_2 FILLER_46_711 ();
 sg13g2_fill_2 FILLER_46_722 ();
 sg13g2_fill_2 FILLER_46_751 ();
 sg13g2_decap_8 FILLER_46_781 ();
 sg13g2_fill_1 FILLER_46_788 ();
 sg13g2_fill_2 FILLER_46_830 ();
 sg13g2_fill_1 FILLER_46_942 ();
 sg13g2_fill_1 FILLER_46_987 ();
 sg13g2_fill_1 FILLER_46_994 ();
 sg13g2_fill_2 FILLER_46_1004 ();
 sg13g2_fill_1 FILLER_46_1006 ();
 sg13g2_fill_2 FILLER_46_1016 ();
 sg13g2_fill_1 FILLER_46_1018 ();
 sg13g2_fill_1 FILLER_46_1037 ();
 sg13g2_decap_8 FILLER_46_1053 ();
 sg13g2_fill_1 FILLER_46_1060 ();
 sg13g2_fill_1 FILLER_46_1090 ();
 sg13g2_decap_8 FILLER_46_1140 ();
 sg13g2_decap_8 FILLER_46_1204 ();
 sg13g2_fill_2 FILLER_46_1211 ();
 sg13g2_fill_1 FILLER_46_1213 ();
 sg13g2_fill_2 FILLER_46_1234 ();
 sg13g2_fill_2 FILLER_46_1272 ();
 sg13g2_fill_2 FILLER_46_1283 ();
 sg13g2_fill_2 FILLER_46_1301 ();
 sg13g2_decap_8 FILLER_46_1328 ();
 sg13g2_decap_8 FILLER_46_1335 ();
 sg13g2_decap_8 FILLER_46_1342 ();
 sg13g2_decap_8 FILLER_46_1349 ();
 sg13g2_decap_8 FILLER_46_1356 ();
 sg13g2_decap_4 FILLER_46_1363 ();
 sg13g2_fill_1 FILLER_46_1408 ();
 sg13g2_decap_4 FILLER_46_1417 ();
 sg13g2_fill_1 FILLER_46_1421 ();
 sg13g2_decap_4 FILLER_46_1427 ();
 sg13g2_fill_2 FILLER_46_1431 ();
 sg13g2_decap_4 FILLER_46_1444 ();
 sg13g2_fill_2 FILLER_46_1480 ();
 sg13g2_decap_8 FILLER_46_1517 ();
 sg13g2_fill_2 FILLER_46_1629 ();
 sg13g2_fill_1 FILLER_46_1631 ();
 sg13g2_fill_2 FILLER_46_1655 ();
 sg13g2_fill_2 FILLER_46_1683 ();
 sg13g2_fill_1 FILLER_46_1685 ();
 sg13g2_decap_8 FILLER_46_1720 ();
 sg13g2_decap_8 FILLER_46_1736 ();
 sg13g2_decap_8 FILLER_46_1743 ();
 sg13g2_decap_4 FILLER_46_1750 ();
 sg13g2_fill_1 FILLER_46_1754 ();
 sg13g2_decap_8 FILLER_46_1764 ();
 sg13g2_fill_2 FILLER_46_1771 ();
 sg13g2_fill_1 FILLER_46_1773 ();
 sg13g2_fill_2 FILLER_46_1778 ();
 sg13g2_fill_1 FILLER_46_1780 ();
 sg13g2_fill_1 FILLER_46_1789 ();
 sg13g2_decap_4 FILLER_46_1832 ();
 sg13g2_fill_2 FILLER_46_1836 ();
 sg13g2_fill_1 FILLER_46_1841 ();
 sg13g2_decap_8 FILLER_46_1911 ();
 sg13g2_fill_2 FILLER_46_1918 ();
 sg13g2_fill_1 FILLER_46_1920 ();
 sg13g2_decap_8 FILLER_46_1924 ();
 sg13g2_fill_1 FILLER_46_1931 ();
 sg13g2_fill_2 FILLER_46_2001 ();
 sg13g2_fill_1 FILLER_46_2042 ();
 sg13g2_decap_8 FILLER_46_2060 ();
 sg13g2_decap_4 FILLER_46_2067 ();
 sg13g2_fill_2 FILLER_46_2112 ();
 sg13g2_fill_1 FILLER_46_2114 ();
 sg13g2_fill_2 FILLER_46_2304 ();
 sg13g2_decap_8 FILLER_46_2319 ();
 sg13g2_decap_4 FILLER_46_2326 ();
 sg13g2_fill_1 FILLER_46_2343 ();
 sg13g2_decap_8 FILLER_46_2405 ();
 sg13g2_decap_8 FILLER_46_2412 ();
 sg13g2_decap_8 FILLER_46_2419 ();
 sg13g2_decap_8 FILLER_46_2426 ();
 sg13g2_decap_8 FILLER_46_2433 ();
 sg13g2_decap_8 FILLER_46_2440 ();
 sg13g2_decap_8 FILLER_46_2447 ();
 sg13g2_decap_8 FILLER_46_2454 ();
 sg13g2_decap_8 FILLER_46_2461 ();
 sg13g2_decap_8 FILLER_46_2468 ();
 sg13g2_decap_8 FILLER_46_2475 ();
 sg13g2_decap_8 FILLER_46_2482 ();
 sg13g2_decap_8 FILLER_46_2489 ();
 sg13g2_decap_8 FILLER_46_2496 ();
 sg13g2_decap_8 FILLER_46_2503 ();
 sg13g2_decap_8 FILLER_46_2510 ();
 sg13g2_decap_8 FILLER_46_2517 ();
 sg13g2_decap_8 FILLER_46_2524 ();
 sg13g2_decap_8 FILLER_46_2531 ();
 sg13g2_decap_8 FILLER_46_2538 ();
 sg13g2_decap_8 FILLER_46_2545 ();
 sg13g2_decap_8 FILLER_46_2552 ();
 sg13g2_decap_8 FILLER_46_2559 ();
 sg13g2_decap_8 FILLER_46_2566 ();
 sg13g2_decap_8 FILLER_46_2573 ();
 sg13g2_decap_8 FILLER_46_2580 ();
 sg13g2_decap_8 FILLER_46_2587 ();
 sg13g2_decap_8 FILLER_46_2594 ();
 sg13g2_decap_8 FILLER_46_2601 ();
 sg13g2_decap_8 FILLER_46_2608 ();
 sg13g2_decap_8 FILLER_46_2615 ();
 sg13g2_decap_8 FILLER_46_2622 ();
 sg13g2_decap_8 FILLER_46_2629 ();
 sg13g2_decap_8 FILLER_46_2636 ();
 sg13g2_decap_8 FILLER_46_2643 ();
 sg13g2_decap_8 FILLER_46_2650 ();
 sg13g2_decap_8 FILLER_46_2657 ();
 sg13g2_decap_8 FILLER_46_2664 ();
 sg13g2_fill_2 FILLER_46_2671 ();
 sg13g2_fill_1 FILLER_46_2673 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_fill_2 FILLER_47_74 ();
 sg13g2_fill_1 FILLER_47_76 ();
 sg13g2_decap_8 FILLER_47_95 ();
 sg13g2_decap_4 FILLER_47_102 ();
 sg13g2_fill_2 FILLER_47_106 ();
 sg13g2_fill_1 FILLER_47_200 ();
 sg13g2_decap_4 FILLER_47_214 ();
 sg13g2_fill_2 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_229 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_299 ();
 sg13g2_fill_2 FILLER_47_350 ();
 sg13g2_decap_4 FILLER_47_426 ();
 sg13g2_fill_1 FILLER_47_430 ();
 sg13g2_fill_1 FILLER_47_435 ();
 sg13g2_decap_8 FILLER_47_449 ();
 sg13g2_fill_1 FILLER_47_456 ();
 sg13g2_decap_4 FILLER_47_493 ();
 sg13g2_fill_2 FILLER_47_497 ();
 sg13g2_decap_4 FILLER_47_537 ();
 sg13g2_fill_2 FILLER_47_541 ();
 sg13g2_fill_1 FILLER_47_638 ();
 sg13g2_decap_4 FILLER_47_652 ();
 sg13g2_fill_2 FILLER_47_656 ();
 sg13g2_fill_1 FILLER_47_663 ();
 sg13g2_decap_4 FILLER_47_687 ();
 sg13g2_fill_1 FILLER_47_691 ();
 sg13g2_fill_2 FILLER_47_699 ();
 sg13g2_decap_8 FILLER_47_718 ();
 sg13g2_fill_1 FILLER_47_737 ();
 sg13g2_decap_4 FILLER_47_751 ();
 sg13g2_fill_1 FILLER_47_755 ();
 sg13g2_decap_4 FILLER_47_784 ();
 sg13g2_fill_1 FILLER_47_805 ();
 sg13g2_fill_1 FILLER_47_843 ();
 sg13g2_fill_2 FILLER_47_857 ();
 sg13g2_fill_1 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_878 ();
 sg13g2_fill_1 FILLER_47_910 ();
 sg13g2_fill_1 FILLER_47_917 ();
 sg13g2_fill_1 FILLER_47_1046 ();
 sg13g2_fill_1 FILLER_47_1062 ();
 sg13g2_decap_4 FILLER_47_1087 ();
 sg13g2_fill_1 FILLER_47_1091 ();
 sg13g2_decap_8 FILLER_47_1144 ();
 sg13g2_decap_8 FILLER_47_1151 ();
 sg13g2_fill_2 FILLER_47_1158 ();
 sg13g2_fill_1 FILLER_47_1160 ();
 sg13g2_decap_8 FILLER_47_1201 ();
 sg13g2_decap_8 FILLER_47_1208 ();
 sg13g2_decap_8 FILLER_47_1215 ();
 sg13g2_decap_8 FILLER_47_1222 ();
 sg13g2_fill_2 FILLER_47_1245 ();
 sg13g2_fill_2 FILLER_47_1252 ();
 sg13g2_fill_1 FILLER_47_1279 ();
 sg13g2_fill_1 FILLER_47_1304 ();
 sg13g2_decap_8 FILLER_47_1323 ();
 sg13g2_decap_8 FILLER_47_1339 ();
 sg13g2_decap_8 FILLER_47_1346 ();
 sg13g2_decap_4 FILLER_47_1353 ();
 sg13g2_decap_8 FILLER_47_1360 ();
 sg13g2_decap_8 FILLER_47_1367 ();
 sg13g2_decap_8 FILLER_47_1374 ();
 sg13g2_fill_1 FILLER_47_1381 ();
 sg13g2_fill_1 FILLER_47_1413 ();
 sg13g2_decap_4 FILLER_47_1427 ();
 sg13g2_decap_8 FILLER_47_1463 ();
 sg13g2_fill_1 FILLER_47_1470 ();
 sg13g2_decap_8 FILLER_47_1509 ();
 sg13g2_fill_2 FILLER_47_1516 ();
 sg13g2_fill_2 FILLER_47_1523 ();
 sg13g2_fill_1 FILLER_47_1525 ();
 sg13g2_fill_2 FILLER_47_1579 ();
 sg13g2_fill_1 FILLER_47_1621 ();
 sg13g2_fill_2 FILLER_47_1660 ();
 sg13g2_fill_1 FILLER_47_1662 ();
 sg13g2_fill_2 FILLER_47_1712 ();
 sg13g2_fill_1 FILLER_47_1714 ();
 sg13g2_decap_4 FILLER_47_1723 ();
 sg13g2_fill_1 FILLER_47_1727 ();
 sg13g2_decap_8 FILLER_47_1735 ();
 sg13g2_decap_4 FILLER_47_1742 ();
 sg13g2_fill_1 FILLER_47_1746 ();
 sg13g2_decap_8 FILLER_47_1752 ();
 sg13g2_decap_4 FILLER_47_1759 ();
 sg13g2_fill_1 FILLER_47_1767 ();
 sg13g2_fill_1 FILLER_47_1796 ();
 sg13g2_decap_8 FILLER_47_1817 ();
 sg13g2_fill_1 FILLER_47_1837 ();
 sg13g2_fill_1 FILLER_47_1850 ();
 sg13g2_fill_1 FILLER_47_1877 ();
 sg13g2_fill_1 FILLER_47_1888 ();
 sg13g2_fill_2 FILLER_47_1916 ();
 sg13g2_fill_1 FILLER_47_1930 ();
 sg13g2_decap_4 FILLER_47_1939 ();
 sg13g2_fill_1 FILLER_47_1943 ();
 sg13g2_fill_1 FILLER_47_1953 ();
 sg13g2_fill_1 FILLER_47_2014 ();
 sg13g2_decap_4 FILLER_47_2121 ();
 sg13g2_fill_1 FILLER_47_2125 ();
 sg13g2_decap_8 FILLER_47_2184 ();
 sg13g2_decap_8 FILLER_47_2191 ();
 sg13g2_fill_1 FILLER_47_2225 ();
 sg13g2_fill_1 FILLER_47_2316 ();
 sg13g2_fill_2 FILLER_47_2387 ();
 sg13g2_decap_8 FILLER_47_2392 ();
 sg13g2_decap_8 FILLER_47_2399 ();
 sg13g2_decap_8 FILLER_47_2406 ();
 sg13g2_decap_8 FILLER_47_2413 ();
 sg13g2_decap_8 FILLER_47_2420 ();
 sg13g2_decap_8 FILLER_47_2427 ();
 sg13g2_decap_8 FILLER_47_2434 ();
 sg13g2_decap_8 FILLER_47_2441 ();
 sg13g2_decap_8 FILLER_47_2448 ();
 sg13g2_decap_8 FILLER_47_2455 ();
 sg13g2_decap_8 FILLER_47_2462 ();
 sg13g2_decap_8 FILLER_47_2469 ();
 sg13g2_decap_8 FILLER_47_2476 ();
 sg13g2_decap_8 FILLER_47_2483 ();
 sg13g2_decap_8 FILLER_47_2490 ();
 sg13g2_decap_8 FILLER_47_2497 ();
 sg13g2_decap_8 FILLER_47_2504 ();
 sg13g2_decap_8 FILLER_47_2511 ();
 sg13g2_decap_8 FILLER_47_2518 ();
 sg13g2_decap_8 FILLER_47_2525 ();
 sg13g2_decap_8 FILLER_47_2532 ();
 sg13g2_decap_8 FILLER_47_2539 ();
 sg13g2_decap_8 FILLER_47_2546 ();
 sg13g2_decap_8 FILLER_47_2553 ();
 sg13g2_decap_8 FILLER_47_2560 ();
 sg13g2_decap_8 FILLER_47_2567 ();
 sg13g2_decap_8 FILLER_47_2574 ();
 sg13g2_decap_8 FILLER_47_2581 ();
 sg13g2_decap_8 FILLER_47_2588 ();
 sg13g2_decap_8 FILLER_47_2595 ();
 sg13g2_decap_8 FILLER_47_2602 ();
 sg13g2_decap_8 FILLER_47_2609 ();
 sg13g2_decap_8 FILLER_47_2616 ();
 sg13g2_decap_8 FILLER_47_2623 ();
 sg13g2_decap_8 FILLER_47_2630 ();
 sg13g2_decap_8 FILLER_47_2637 ();
 sg13g2_decap_8 FILLER_47_2644 ();
 sg13g2_decap_8 FILLER_47_2651 ();
 sg13g2_decap_8 FILLER_47_2658 ();
 sg13g2_decap_8 FILLER_47_2665 ();
 sg13g2_fill_2 FILLER_47_2672 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_fill_2 FILLER_48_77 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_fill_1 FILLER_48_157 ();
 sg13g2_fill_2 FILLER_48_247 ();
 sg13g2_fill_2 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_323 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_fill_1 FILLER_48_358 ();
 sg13g2_fill_2 FILLER_48_421 ();
 sg13g2_decap_4 FILLER_48_427 ();
 sg13g2_fill_2 FILLER_48_453 ();
 sg13g2_fill_1 FILLER_48_466 ();
 sg13g2_decap_8 FILLER_48_494 ();
 sg13g2_fill_1 FILLER_48_547 ();
 sg13g2_fill_1 FILLER_48_570 ();
 sg13g2_fill_2 FILLER_48_583 ();
 sg13g2_fill_1 FILLER_48_600 ();
 sg13g2_fill_1 FILLER_48_614 ();
 sg13g2_fill_1 FILLER_48_620 ();
 sg13g2_fill_1 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_677 ();
 sg13g2_decap_4 FILLER_48_684 ();
 sg13g2_fill_2 FILLER_48_688 ();
 sg13g2_decap_8 FILLER_48_712 ();
 sg13g2_decap_8 FILLER_48_719 ();
 sg13g2_fill_1 FILLER_48_726 ();
 sg13g2_fill_2 FILLER_48_747 ();
 sg13g2_decap_4 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_fill_2 FILLER_48_787 ();
 sg13g2_fill_2 FILLER_48_817 ();
 sg13g2_fill_2 FILLER_48_836 ();
 sg13g2_fill_2 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_fill_2 FILLER_48_856 ();
 sg13g2_fill_1 FILLER_48_858 ();
 sg13g2_fill_2 FILLER_48_873 ();
 sg13g2_fill_1 FILLER_48_875 ();
 sg13g2_fill_2 FILLER_48_880 ();
 sg13g2_fill_1 FILLER_48_882 ();
 sg13g2_fill_1 FILLER_48_902 ();
 sg13g2_fill_2 FILLER_48_913 ();
 sg13g2_fill_1 FILLER_48_998 ();
 sg13g2_fill_1 FILLER_48_1034 ();
 sg13g2_fill_2 FILLER_48_1041 ();
 sg13g2_fill_1 FILLER_48_1073 ();
 sg13g2_fill_2 FILLER_48_1108 ();
 sg13g2_fill_1 FILLER_48_1110 ();
 sg13g2_fill_2 FILLER_48_1119 ();
 sg13g2_fill_1 FILLER_48_1121 ();
 sg13g2_decap_8 FILLER_48_1140 ();
 sg13g2_decap_8 FILLER_48_1147 ();
 sg13g2_decap_4 FILLER_48_1217 ();
 sg13g2_fill_1 FILLER_48_1221 ();
 sg13g2_fill_2 FILLER_48_1260 ();
 sg13g2_fill_2 FILLER_48_1289 ();
 sg13g2_fill_1 FILLER_48_1300 ();
 sg13g2_fill_2 FILLER_48_1318 ();
 sg13g2_fill_1 FILLER_48_1350 ();
 sg13g2_decap_8 FILLER_48_1372 ();
 sg13g2_decap_8 FILLER_48_1379 ();
 sg13g2_decap_8 FILLER_48_1386 ();
 sg13g2_decap_4 FILLER_48_1393 ();
 sg13g2_fill_2 FILLER_48_1397 ();
 sg13g2_decap_4 FILLER_48_1404 ();
 sg13g2_fill_2 FILLER_48_1408 ();
 sg13g2_fill_1 FILLER_48_1415 ();
 sg13g2_fill_2 FILLER_48_1442 ();
 sg13g2_fill_1 FILLER_48_1444 ();
 sg13g2_decap_8 FILLER_48_1463 ();
 sg13g2_decap_8 FILLER_48_1470 ();
 sg13g2_decap_4 FILLER_48_1477 ();
 sg13g2_fill_2 FILLER_48_1500 ();
 sg13g2_fill_2 FILLER_48_1507 ();
 sg13g2_fill_1 FILLER_48_1509 ();
 sg13g2_fill_1 FILLER_48_1522 ();
 sg13g2_fill_2 FILLER_48_1559 ();
 sg13g2_fill_1 FILLER_48_1561 ();
 sg13g2_fill_2 FILLER_48_1595 ();
 sg13g2_fill_1 FILLER_48_1597 ();
 sg13g2_fill_1 FILLER_48_1686 ();
 sg13g2_fill_1 FILLER_48_1700 ();
 sg13g2_fill_1 FILLER_48_1728 ();
 sg13g2_fill_2 FILLER_48_1734 ();
 sg13g2_fill_1 FILLER_48_1736 ();
 sg13g2_fill_1 FILLER_48_1812 ();
 sg13g2_decap_8 FILLER_48_1822 ();
 sg13g2_decap_4 FILLER_48_1829 ();
 sg13g2_fill_1 FILLER_48_1896 ();
 sg13g2_decap_8 FILLER_48_1963 ();
 sg13g2_fill_1 FILLER_48_1970 ();
 sg13g2_decap_4 FILLER_48_1976 ();
 sg13g2_fill_1 FILLER_48_1993 ();
 sg13g2_decap_4 FILLER_48_2000 ();
 sg13g2_fill_2 FILLER_48_2004 ();
 sg13g2_decap_4 FILLER_48_2019 ();
 sg13g2_fill_1 FILLER_48_2071 ();
 sg13g2_fill_2 FILLER_48_2123 ();
 sg13g2_fill_2 FILLER_48_2152 ();
 sg13g2_fill_1 FILLER_48_2154 ();
 sg13g2_decap_8 FILLER_48_2182 ();
 sg13g2_fill_1 FILLER_48_2189 ();
 sg13g2_fill_2 FILLER_48_2225 ();
 sg13g2_fill_1 FILLER_48_2227 ();
 sg13g2_fill_1 FILLER_48_2265 ();
 sg13g2_fill_2 FILLER_48_2271 ();
 sg13g2_fill_1 FILLER_48_2273 ();
 sg13g2_fill_2 FILLER_48_2330 ();
 sg13g2_fill_1 FILLER_48_2361 ();
 sg13g2_decap_8 FILLER_48_2374 ();
 sg13g2_decap_8 FILLER_48_2381 ();
 sg13g2_decap_8 FILLER_48_2388 ();
 sg13g2_decap_8 FILLER_48_2395 ();
 sg13g2_decap_8 FILLER_48_2402 ();
 sg13g2_decap_8 FILLER_48_2409 ();
 sg13g2_decap_8 FILLER_48_2416 ();
 sg13g2_decap_8 FILLER_48_2423 ();
 sg13g2_decap_8 FILLER_48_2430 ();
 sg13g2_decap_8 FILLER_48_2437 ();
 sg13g2_decap_8 FILLER_48_2444 ();
 sg13g2_decap_8 FILLER_48_2451 ();
 sg13g2_decap_8 FILLER_48_2458 ();
 sg13g2_decap_8 FILLER_48_2465 ();
 sg13g2_decap_8 FILLER_48_2472 ();
 sg13g2_decap_8 FILLER_48_2479 ();
 sg13g2_decap_8 FILLER_48_2486 ();
 sg13g2_decap_8 FILLER_48_2493 ();
 sg13g2_decap_8 FILLER_48_2500 ();
 sg13g2_decap_8 FILLER_48_2507 ();
 sg13g2_decap_8 FILLER_48_2514 ();
 sg13g2_decap_8 FILLER_48_2521 ();
 sg13g2_decap_8 FILLER_48_2528 ();
 sg13g2_decap_8 FILLER_48_2535 ();
 sg13g2_decap_8 FILLER_48_2542 ();
 sg13g2_decap_8 FILLER_48_2549 ();
 sg13g2_decap_8 FILLER_48_2556 ();
 sg13g2_decap_8 FILLER_48_2563 ();
 sg13g2_decap_8 FILLER_48_2570 ();
 sg13g2_decap_8 FILLER_48_2577 ();
 sg13g2_decap_8 FILLER_48_2584 ();
 sg13g2_decap_8 FILLER_48_2591 ();
 sg13g2_decap_8 FILLER_48_2598 ();
 sg13g2_decap_8 FILLER_48_2605 ();
 sg13g2_decap_8 FILLER_48_2612 ();
 sg13g2_decap_8 FILLER_48_2619 ();
 sg13g2_decap_8 FILLER_48_2626 ();
 sg13g2_decap_8 FILLER_48_2633 ();
 sg13g2_decap_8 FILLER_48_2640 ();
 sg13g2_decap_8 FILLER_48_2647 ();
 sg13g2_decap_8 FILLER_48_2654 ();
 sg13g2_decap_8 FILLER_48_2661 ();
 sg13g2_decap_4 FILLER_48_2668 ();
 sg13g2_fill_2 FILLER_48_2672 ();
 sg13g2_fill_2 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_68 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_107 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_195 ();
 sg13g2_fill_2 FILLER_49_277 ();
 sg13g2_fill_2 FILLER_49_318 ();
 sg13g2_fill_1 FILLER_49_320 ();
 sg13g2_fill_1 FILLER_49_342 ();
 sg13g2_decap_8 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_359 ();
 sg13g2_fill_2 FILLER_49_421 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_461 ();
 sg13g2_decap_8 FILLER_49_498 ();
 sg13g2_decap_8 FILLER_49_505 ();
 sg13g2_decap_8 FILLER_49_512 ();
 sg13g2_fill_2 FILLER_49_519 ();
 sg13g2_fill_2 FILLER_49_556 ();
 sg13g2_fill_2 FILLER_49_606 ();
 sg13g2_fill_2 FILLER_49_634 ();
 sg13g2_decap_4 FILLER_49_726 ();
 sg13g2_fill_2 FILLER_49_730 ();
 sg13g2_fill_2 FILLER_49_789 ();
 sg13g2_fill_1 FILLER_49_791 ();
 sg13g2_fill_1 FILLER_49_806 ();
 sg13g2_fill_2 FILLER_49_816 ();
 sg13g2_fill_1 FILLER_49_848 ();
 sg13g2_fill_1 FILLER_49_904 ();
 sg13g2_decap_8 FILLER_49_914 ();
 sg13g2_decap_8 FILLER_49_921 ();
 sg13g2_fill_2 FILLER_49_980 ();
 sg13g2_fill_1 FILLER_49_1010 ();
 sg13g2_fill_2 FILLER_49_1041 ();
 sg13g2_fill_1 FILLER_49_1043 ();
 sg13g2_fill_1 FILLER_49_1057 ();
 sg13g2_fill_1 FILLER_49_1068 ();
 sg13g2_decap_8 FILLER_49_1073 ();
 sg13g2_fill_1 FILLER_49_1080 ();
 sg13g2_fill_2 FILLER_49_1094 ();
 sg13g2_decap_8 FILLER_49_1101 ();
 sg13g2_fill_2 FILLER_49_1133 ();
 sg13g2_fill_1 FILLER_49_1135 ();
 sg13g2_decap_8 FILLER_49_1145 ();
 sg13g2_fill_1 FILLER_49_1175 ();
 sg13g2_fill_2 FILLER_49_1231 ();
 sg13g2_fill_2 FILLER_49_1251 ();
 sg13g2_fill_1 FILLER_49_1312 ();
 sg13g2_fill_1 FILLER_49_1336 ();
 sg13g2_decap_8 FILLER_49_1396 ();
 sg13g2_fill_2 FILLER_49_1403 ();
 sg13g2_fill_1 FILLER_49_1410 ();
 sg13g2_fill_2 FILLER_49_1415 ();
 sg13g2_fill_1 FILLER_49_1417 ();
 sg13g2_decap_4 FILLER_49_1469 ();
 sg13g2_fill_2 FILLER_49_1473 ();
 sg13g2_fill_2 FILLER_49_1491 ();
 sg13g2_fill_1 FILLER_49_1502 ();
 sg13g2_fill_1 FILLER_49_1520 ();
 sg13g2_decap_8 FILLER_49_1526 ();
 sg13g2_decap_8 FILLER_49_1533 ();
 sg13g2_fill_2 FILLER_49_1540 ();
 sg13g2_fill_1 FILLER_49_1542 ();
 sg13g2_decap_8 FILLER_49_1557 ();
 sg13g2_decap_4 FILLER_49_1564 ();
 sg13g2_fill_1 FILLER_49_1577 ();
 sg13g2_decap_4 FILLER_49_1596 ();
 sg13g2_fill_1 FILLER_49_1674 ();
 sg13g2_fill_2 FILLER_49_1690 ();
 sg13g2_fill_1 FILLER_49_1692 ();
 sg13g2_decap_4 FILLER_49_1734 ();
 sg13g2_fill_2 FILLER_49_1783 ();
 sg13g2_fill_1 FILLER_49_1785 ();
 sg13g2_fill_1 FILLER_49_1829 ();
 sg13g2_decap_8 FILLER_49_1839 ();
 sg13g2_fill_2 FILLER_49_1846 ();
 sg13g2_fill_1 FILLER_49_1848 ();
 sg13g2_fill_2 FILLER_49_1898 ();
 sg13g2_decap_8 FILLER_49_1959 ();
 sg13g2_decap_8 FILLER_49_1966 ();
 sg13g2_decap_8 FILLER_49_1973 ();
 sg13g2_decap_8 FILLER_49_1980 ();
 sg13g2_decap_8 FILLER_49_1987 ();
 sg13g2_decap_8 FILLER_49_1994 ();
 sg13g2_decap_8 FILLER_49_2001 ();
 sg13g2_decap_8 FILLER_49_2012 ();
 sg13g2_decap_8 FILLER_49_2019 ();
 sg13g2_decap_8 FILLER_49_2054 ();
 sg13g2_fill_1 FILLER_49_2061 ();
 sg13g2_decap_8 FILLER_49_2075 ();
 sg13g2_decap_4 FILLER_49_2082 ();
 sg13g2_fill_2 FILLER_49_2086 ();
 sg13g2_decap_8 FILLER_49_2117 ();
 sg13g2_decap_8 FILLER_49_2127 ();
 sg13g2_fill_2 FILLER_49_2134 ();
 sg13g2_fill_1 FILLER_49_2136 ();
 sg13g2_decap_4 FILLER_49_2179 ();
 sg13g2_fill_2 FILLER_49_2183 ();
 sg13g2_fill_2 FILLER_49_2217 ();
 sg13g2_fill_2 FILLER_49_2228 ();
 sg13g2_fill_1 FILLER_49_2230 ();
 sg13g2_decap_8 FILLER_49_2304 ();
 sg13g2_decap_8 FILLER_49_2311 ();
 sg13g2_decap_4 FILLER_49_2318 ();
 sg13g2_fill_1 FILLER_49_2322 ();
 sg13g2_decap_8 FILLER_49_2382 ();
 sg13g2_decap_8 FILLER_49_2389 ();
 sg13g2_decap_8 FILLER_49_2396 ();
 sg13g2_decap_8 FILLER_49_2403 ();
 sg13g2_decap_8 FILLER_49_2410 ();
 sg13g2_decap_8 FILLER_49_2417 ();
 sg13g2_decap_8 FILLER_49_2424 ();
 sg13g2_decap_8 FILLER_49_2431 ();
 sg13g2_decap_8 FILLER_49_2438 ();
 sg13g2_decap_8 FILLER_49_2445 ();
 sg13g2_decap_8 FILLER_49_2452 ();
 sg13g2_decap_8 FILLER_49_2459 ();
 sg13g2_decap_8 FILLER_49_2466 ();
 sg13g2_decap_8 FILLER_49_2473 ();
 sg13g2_decap_8 FILLER_49_2480 ();
 sg13g2_decap_8 FILLER_49_2487 ();
 sg13g2_decap_8 FILLER_49_2494 ();
 sg13g2_decap_8 FILLER_49_2501 ();
 sg13g2_decap_8 FILLER_49_2508 ();
 sg13g2_decap_8 FILLER_49_2515 ();
 sg13g2_decap_8 FILLER_49_2522 ();
 sg13g2_decap_8 FILLER_49_2529 ();
 sg13g2_decap_8 FILLER_49_2536 ();
 sg13g2_decap_8 FILLER_49_2543 ();
 sg13g2_decap_8 FILLER_49_2550 ();
 sg13g2_decap_8 FILLER_49_2557 ();
 sg13g2_decap_8 FILLER_49_2564 ();
 sg13g2_decap_8 FILLER_49_2571 ();
 sg13g2_decap_8 FILLER_49_2578 ();
 sg13g2_decap_8 FILLER_49_2585 ();
 sg13g2_decap_8 FILLER_49_2592 ();
 sg13g2_decap_8 FILLER_49_2599 ();
 sg13g2_decap_8 FILLER_49_2606 ();
 sg13g2_decap_8 FILLER_49_2613 ();
 sg13g2_decap_8 FILLER_49_2620 ();
 sg13g2_decap_8 FILLER_49_2627 ();
 sg13g2_decap_8 FILLER_49_2634 ();
 sg13g2_decap_8 FILLER_49_2641 ();
 sg13g2_decap_8 FILLER_49_2648 ();
 sg13g2_decap_8 FILLER_49_2655 ();
 sg13g2_decap_8 FILLER_49_2662 ();
 sg13g2_decap_4 FILLER_49_2669 ();
 sg13g2_fill_1 FILLER_49_2673 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_2 FILLER_50_47 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_fill_1 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_288 ();
 sg13g2_fill_2 FILLER_50_349 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_fill_1 FILLER_50_421 ();
 sg13g2_fill_1 FILLER_50_469 ();
 sg13g2_fill_2 FILLER_50_484 ();
 sg13g2_fill_1 FILLER_50_486 ();
 sg13g2_decap_8 FILLER_50_514 ();
 sg13g2_decap_4 FILLER_50_521 ();
 sg13g2_fill_1 FILLER_50_525 ();
 sg13g2_fill_2 FILLER_50_539 ();
 sg13g2_fill_1 FILLER_50_577 ();
 sg13g2_decap_4 FILLER_50_606 ();
 sg13g2_fill_1 FILLER_50_610 ();
 sg13g2_fill_1 FILLER_50_639 ();
 sg13g2_fill_2 FILLER_50_684 ();
 sg13g2_fill_1 FILLER_50_686 ();
 sg13g2_decap_4 FILLER_50_700 ();
 sg13g2_fill_1 FILLER_50_704 ();
 sg13g2_fill_1 FILLER_50_746 ();
 sg13g2_fill_2 FILLER_50_819 ();
 sg13g2_fill_1 FILLER_50_874 ();
 sg13g2_fill_1 FILLER_50_879 ();
 sg13g2_decap_8 FILLER_50_916 ();
 sg13g2_fill_2 FILLER_50_923 ();
 sg13g2_fill_1 FILLER_50_938 ();
 sg13g2_decap_4 FILLER_50_1003 ();
 sg13g2_fill_2 FILLER_50_1007 ();
 sg13g2_fill_2 FILLER_50_1031 ();
 sg13g2_fill_2 FILLER_50_1038 ();
 sg13g2_decap_8 FILLER_50_1048 ();
 sg13g2_fill_2 FILLER_50_1055 ();
 sg13g2_fill_1 FILLER_50_1082 ();
 sg13g2_decap_4 FILLER_50_1096 ();
 sg13g2_decap_8 FILLER_50_1109 ();
 sg13g2_decap_8 FILLER_50_1116 ();
 sg13g2_fill_1 FILLER_50_1123 ();
 sg13g2_fill_1 FILLER_50_1191 ();
 sg13g2_fill_1 FILLER_50_1335 ();
 sg13g2_fill_1 FILLER_50_1405 ();
 sg13g2_fill_1 FILLER_50_1423 ();
 sg13g2_fill_2 FILLER_50_1438 ();
 sg13g2_fill_2 FILLER_50_1463 ();
 sg13g2_fill_1 FILLER_50_1465 ();
 sg13g2_fill_2 FILLER_50_1473 ();
 sg13g2_fill_2 FILLER_50_1510 ();
 sg13g2_fill_1 FILLER_50_1512 ();
 sg13g2_decap_4 FILLER_50_1541 ();
 sg13g2_fill_2 FILLER_50_1557 ();
 sg13g2_fill_1 FILLER_50_1559 ();
 sg13g2_fill_2 FILLER_50_1569 ();
 sg13g2_fill_2 FILLER_50_1582 ();
 sg13g2_fill_2 FILLER_50_1607 ();
 sg13g2_fill_1 FILLER_50_1609 ();
 sg13g2_fill_1 FILLER_50_1631 ();
 sg13g2_fill_2 FILLER_50_1699 ();
 sg13g2_fill_1 FILLER_50_1701 ();
 sg13g2_decap_4 FILLER_50_1725 ();
 sg13g2_fill_1 FILLER_50_1729 ();
 sg13g2_decap_8 FILLER_50_1738 ();
 sg13g2_fill_2 FILLER_50_1859 ();
 sg13g2_fill_1 FILLER_50_1906 ();
 sg13g2_fill_2 FILLER_50_1937 ();
 sg13g2_decap_4 FILLER_50_1978 ();
 sg13g2_fill_2 FILLER_50_1982 ();
 sg13g2_fill_1 FILLER_50_1991 ();
 sg13g2_fill_1 FILLER_50_2041 ();
 sg13g2_fill_2 FILLER_50_2061 ();
 sg13g2_decap_8 FILLER_50_2069 ();
 sg13g2_fill_2 FILLER_50_2076 ();
 sg13g2_fill_1 FILLER_50_2078 ();
 sg13g2_decap_8 FILLER_50_2083 ();
 sg13g2_decap_4 FILLER_50_2090 ();
 sg13g2_fill_1 FILLER_50_2094 ();
 sg13g2_fill_1 FILLER_50_2109 ();
 sg13g2_decap_8 FILLER_50_2113 ();
 sg13g2_fill_2 FILLER_50_2120 ();
 sg13g2_fill_1 FILLER_50_2122 ();
 sg13g2_fill_2 FILLER_50_2151 ();
 sg13g2_fill_1 FILLER_50_2153 ();
 sg13g2_decap_4 FILLER_50_2162 ();
 sg13g2_fill_2 FILLER_50_2166 ();
 sg13g2_decap_4 FILLER_50_2174 ();
 sg13g2_fill_1 FILLER_50_2178 ();
 sg13g2_fill_2 FILLER_50_2228 ();
 sg13g2_fill_1 FILLER_50_2230 ();
 sg13g2_fill_2 FILLER_50_2261 ();
 sg13g2_fill_2 FILLER_50_2277 ();
 sg13g2_fill_1 FILLER_50_2279 ();
 sg13g2_fill_2 FILLER_50_2301 ();
 sg13g2_fill_1 FILLER_50_2303 ();
 sg13g2_decap_4 FILLER_50_2317 ();
 sg13g2_fill_1 FILLER_50_2321 ();
 sg13g2_decap_4 FILLER_50_2326 ();
 sg13g2_decap_8 FILLER_50_2374 ();
 sg13g2_decap_8 FILLER_50_2381 ();
 sg13g2_decap_8 FILLER_50_2388 ();
 sg13g2_decap_8 FILLER_50_2395 ();
 sg13g2_decap_8 FILLER_50_2402 ();
 sg13g2_decap_8 FILLER_50_2409 ();
 sg13g2_decap_8 FILLER_50_2416 ();
 sg13g2_decap_8 FILLER_50_2423 ();
 sg13g2_decap_8 FILLER_50_2430 ();
 sg13g2_decap_8 FILLER_50_2437 ();
 sg13g2_decap_8 FILLER_50_2444 ();
 sg13g2_decap_8 FILLER_50_2451 ();
 sg13g2_decap_8 FILLER_50_2458 ();
 sg13g2_decap_8 FILLER_50_2465 ();
 sg13g2_decap_8 FILLER_50_2472 ();
 sg13g2_decap_8 FILLER_50_2479 ();
 sg13g2_decap_8 FILLER_50_2486 ();
 sg13g2_decap_8 FILLER_50_2493 ();
 sg13g2_decap_8 FILLER_50_2500 ();
 sg13g2_decap_8 FILLER_50_2507 ();
 sg13g2_decap_8 FILLER_50_2514 ();
 sg13g2_decap_8 FILLER_50_2521 ();
 sg13g2_decap_8 FILLER_50_2528 ();
 sg13g2_decap_8 FILLER_50_2535 ();
 sg13g2_decap_8 FILLER_50_2542 ();
 sg13g2_decap_8 FILLER_50_2549 ();
 sg13g2_decap_8 FILLER_50_2556 ();
 sg13g2_decap_8 FILLER_50_2563 ();
 sg13g2_decap_8 FILLER_50_2570 ();
 sg13g2_decap_8 FILLER_50_2577 ();
 sg13g2_decap_8 FILLER_50_2584 ();
 sg13g2_decap_8 FILLER_50_2591 ();
 sg13g2_decap_8 FILLER_50_2598 ();
 sg13g2_decap_8 FILLER_50_2605 ();
 sg13g2_decap_8 FILLER_50_2612 ();
 sg13g2_decap_8 FILLER_50_2619 ();
 sg13g2_decap_8 FILLER_50_2626 ();
 sg13g2_decap_8 FILLER_50_2633 ();
 sg13g2_decap_8 FILLER_50_2640 ();
 sg13g2_decap_8 FILLER_50_2647 ();
 sg13g2_decap_8 FILLER_50_2654 ();
 sg13g2_decap_8 FILLER_50_2661 ();
 sg13g2_decap_4 FILLER_50_2668 ();
 sg13g2_fill_2 FILLER_50_2672 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_fill_1 FILLER_51_34 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_fill_2 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_107 ();
 sg13g2_fill_2 FILLER_51_135 ();
 sg13g2_decap_8 FILLER_51_196 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_fill_2 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_fill_2 FILLER_51_312 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_384 ();
 sg13g2_fill_1 FILLER_51_460 ();
 sg13g2_fill_2 FILLER_51_507 ();
 sg13g2_decap_4 FILLER_51_536 ();
 sg13g2_fill_2 FILLER_51_540 ();
 sg13g2_fill_1 FILLER_51_578 ();
 sg13g2_fill_2 FILLER_51_614 ();
 sg13g2_fill_2 FILLER_51_644 ();
 sg13g2_fill_1 FILLER_51_646 ();
 sg13g2_decap_8 FILLER_51_682 ();
 sg13g2_decap_4 FILLER_51_689 ();
 sg13g2_fill_2 FILLER_51_693 ();
 sg13g2_fill_2 FILLER_51_709 ();
 sg13g2_fill_1 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_740 ();
 sg13g2_fill_1 FILLER_51_809 ();
 sg13g2_fill_2 FILLER_51_869 ();
 sg13g2_fill_1 FILLER_51_871 ();
 sg13g2_fill_2 FILLER_51_948 ();
 sg13g2_fill_1 FILLER_51_950 ();
 sg13g2_fill_1 FILLER_51_1001 ();
 sg13g2_decap_8 FILLER_51_1014 ();
 sg13g2_fill_1 FILLER_51_1021 ();
 sg13g2_fill_2 FILLER_51_1032 ();
 sg13g2_fill_1 FILLER_51_1034 ();
 sg13g2_decap_8 FILLER_51_1057 ();
 sg13g2_decap_8 FILLER_51_1064 ();
 sg13g2_decap_4 FILLER_51_1071 ();
 sg13g2_fill_1 FILLER_51_1075 ();
 sg13g2_fill_1 FILLER_51_1083 ();
 sg13g2_fill_2 FILLER_51_1112 ();
 sg13g2_fill_1 FILLER_51_1114 ();
 sg13g2_fill_1 FILLER_51_1194 ();
 sg13g2_fill_2 FILLER_51_1208 ();
 sg13g2_fill_1 FILLER_51_1247 ();
 sg13g2_fill_1 FILLER_51_1272 ();
 sg13g2_fill_2 FILLER_51_1292 ();
 sg13g2_fill_1 FILLER_51_1368 ();
 sg13g2_fill_1 FILLER_51_1439 ();
 sg13g2_fill_2 FILLER_51_1446 ();
 sg13g2_fill_2 FILLER_51_1453 ();
 sg13g2_fill_2 FILLER_51_1468 ();
 sg13g2_fill_1 FILLER_51_1470 ();
 sg13g2_fill_1 FILLER_51_1499 ();
 sg13g2_fill_1 FILLER_51_1579 ();
 sg13g2_fill_2 FILLER_51_1599 ();
 sg13g2_fill_1 FILLER_51_1601 ();
 sg13g2_fill_2 FILLER_51_1639 ();
 sg13g2_fill_1 FILLER_51_1699 ();
 sg13g2_fill_1 FILLER_51_1754 ();
 sg13g2_decap_4 FILLER_51_1880 ();
 sg13g2_fill_2 FILLER_51_1935 ();
 sg13g2_fill_2 FILLER_51_1968 ();
 sg13g2_decap_4 FILLER_51_2065 ();
 sg13g2_decap_4 FILLER_51_2082 ();
 sg13g2_fill_1 FILLER_51_2086 ();
 sg13g2_decap_8 FILLER_51_2118 ();
 sg13g2_decap_8 FILLER_51_2125 ();
 sg13g2_decap_4 FILLER_51_2132 ();
 sg13g2_fill_1 FILLER_51_2136 ();
 sg13g2_fill_1 FILLER_51_2155 ();
 sg13g2_decap_8 FILLER_51_2170 ();
 sg13g2_fill_1 FILLER_51_2177 ();
 sg13g2_fill_2 FILLER_51_2205 ();
 sg13g2_fill_2 FILLER_51_2234 ();
 sg13g2_fill_1 FILLER_51_2236 ();
 sg13g2_fill_2 FILLER_51_2246 ();
 sg13g2_fill_2 FILLER_51_2279 ();
 sg13g2_fill_1 FILLER_51_2281 ();
 sg13g2_fill_2 FILLER_51_2297 ();
 sg13g2_fill_1 FILLER_51_2299 ();
 sg13g2_decap_8 FILLER_51_2328 ();
 sg13g2_decap_4 FILLER_51_2335 ();
 sg13g2_fill_1 FILLER_51_2339 ();
 sg13g2_fill_2 FILLER_51_2349 ();
 sg13g2_fill_2 FILLER_51_2372 ();
 sg13g2_decap_8 FILLER_51_2377 ();
 sg13g2_decap_8 FILLER_51_2384 ();
 sg13g2_decap_8 FILLER_51_2391 ();
 sg13g2_decap_8 FILLER_51_2398 ();
 sg13g2_decap_8 FILLER_51_2405 ();
 sg13g2_decap_8 FILLER_51_2412 ();
 sg13g2_decap_8 FILLER_51_2419 ();
 sg13g2_decap_8 FILLER_51_2426 ();
 sg13g2_decap_8 FILLER_51_2433 ();
 sg13g2_decap_8 FILLER_51_2440 ();
 sg13g2_decap_8 FILLER_51_2447 ();
 sg13g2_decap_8 FILLER_51_2454 ();
 sg13g2_decap_8 FILLER_51_2461 ();
 sg13g2_decap_8 FILLER_51_2468 ();
 sg13g2_decap_8 FILLER_51_2475 ();
 sg13g2_decap_8 FILLER_51_2482 ();
 sg13g2_decap_8 FILLER_51_2489 ();
 sg13g2_decap_8 FILLER_51_2496 ();
 sg13g2_decap_8 FILLER_51_2503 ();
 sg13g2_decap_8 FILLER_51_2510 ();
 sg13g2_decap_8 FILLER_51_2517 ();
 sg13g2_decap_8 FILLER_51_2524 ();
 sg13g2_decap_8 FILLER_51_2531 ();
 sg13g2_decap_8 FILLER_51_2538 ();
 sg13g2_decap_8 FILLER_51_2545 ();
 sg13g2_decap_8 FILLER_51_2552 ();
 sg13g2_decap_8 FILLER_51_2559 ();
 sg13g2_decap_8 FILLER_51_2566 ();
 sg13g2_decap_8 FILLER_51_2573 ();
 sg13g2_decap_8 FILLER_51_2580 ();
 sg13g2_decap_8 FILLER_51_2587 ();
 sg13g2_decap_8 FILLER_51_2594 ();
 sg13g2_decap_8 FILLER_51_2601 ();
 sg13g2_decap_8 FILLER_51_2608 ();
 sg13g2_decap_8 FILLER_51_2615 ();
 sg13g2_decap_8 FILLER_51_2622 ();
 sg13g2_decap_8 FILLER_51_2629 ();
 sg13g2_decap_8 FILLER_51_2636 ();
 sg13g2_decap_8 FILLER_51_2643 ();
 sg13g2_decap_8 FILLER_51_2650 ();
 sg13g2_decap_8 FILLER_51_2657 ();
 sg13g2_decap_8 FILLER_51_2664 ();
 sg13g2_fill_2 FILLER_51_2671 ();
 sg13g2_fill_1 FILLER_51_2673 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_2 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_42 ();
 sg13g2_fill_2 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_92 ();
 sg13g2_decap_8 FILLER_52_102 ();
 sg13g2_decap_8 FILLER_52_109 ();
 sg13g2_fill_2 FILLER_52_134 ();
 sg13g2_fill_2 FILLER_52_149 ();
 sg13g2_fill_1 FILLER_52_179 ();
 sg13g2_decap_8 FILLER_52_193 ();
 sg13g2_decap_4 FILLER_52_200 ();
 sg13g2_decap_8 FILLER_52_213 ();
 sg13g2_fill_2 FILLER_52_220 ();
 sg13g2_fill_1 FILLER_52_222 ();
 sg13g2_fill_2 FILLER_52_249 ();
 sg13g2_fill_1 FILLER_52_295 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_2 FILLER_52_319 ();
 sg13g2_fill_2 FILLER_52_340 ();
 sg13g2_fill_2 FILLER_52_360 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_fill_2 FILLER_52_382 ();
 sg13g2_decap_8 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_52_435 ();
 sg13g2_fill_2 FILLER_52_440 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_fill_1 FILLER_52_452 ();
 sg13g2_fill_2 FILLER_52_466 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_fill_2 FILLER_52_501 ();
 sg13g2_fill_1 FILLER_52_503 ();
 sg13g2_decap_8 FILLER_52_539 ();
 sg13g2_decap_8 FILLER_52_564 ();
 sg13g2_decap_4 FILLER_52_571 ();
 sg13g2_decap_8 FILLER_52_580 ();
 sg13g2_fill_1 FILLER_52_587 ();
 sg13g2_decap_4 FILLER_52_613 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_fill_1 FILLER_52_626 ();
 sg13g2_decap_8 FILLER_52_636 ();
 sg13g2_decap_8 FILLER_52_643 ();
 sg13g2_decap_4 FILLER_52_650 ();
 sg13g2_fill_1 FILLER_52_654 ();
 sg13g2_decap_8 FILLER_52_683 ();
 sg13g2_fill_1 FILLER_52_690 ();
 sg13g2_fill_2 FILLER_52_741 ();
 sg13g2_fill_1 FILLER_52_743 ();
 sg13g2_fill_2 FILLER_52_765 ();
 sg13g2_fill_1 FILLER_52_767 ();
 sg13g2_fill_2 FILLER_52_915 ();
 sg13g2_fill_1 FILLER_52_917 ();
 sg13g2_fill_1 FILLER_52_931 ();
 sg13g2_fill_2 FILLER_52_980 ();
 sg13g2_fill_2 FILLER_52_991 ();
 sg13g2_fill_1 FILLER_52_1021 ();
 sg13g2_decap_8 FILLER_52_1054 ();
 sg13g2_decap_4 FILLER_52_1102 ();
 sg13g2_fill_1 FILLER_52_1106 ();
 sg13g2_fill_1 FILLER_52_1134 ();
 sg13g2_fill_2 FILLER_52_1166 ();
 sg13g2_fill_2 FILLER_52_1268 ();
 sg13g2_fill_1 FILLER_52_1270 ();
 sg13g2_fill_1 FILLER_52_1323 ();
 sg13g2_fill_2 FILLER_52_1399 ();
 sg13g2_fill_1 FILLER_52_1401 ();
 sg13g2_fill_2 FILLER_52_1448 ();
 sg13g2_fill_2 FILLER_52_1496 ();
 sg13g2_fill_1 FILLER_52_1498 ();
 sg13g2_fill_1 FILLER_52_1507 ();
 sg13g2_decap_4 FILLER_52_1561 ();
 sg13g2_fill_1 FILLER_52_1565 ();
 sg13g2_fill_1 FILLER_52_1587 ();
 sg13g2_decap_8 FILLER_52_1593 ();
 sg13g2_decap_4 FILLER_52_1600 ();
 sg13g2_fill_1 FILLER_52_1612 ();
 sg13g2_fill_1 FILLER_52_1671 ();
 sg13g2_decap_8 FILLER_52_1731 ();
 sg13g2_decap_4 FILLER_52_1738 ();
 sg13g2_fill_1 FILLER_52_1742 ();
 sg13g2_fill_2 FILLER_52_1756 ();
 sg13g2_fill_2 FILLER_52_1800 ();
 sg13g2_fill_1 FILLER_52_1842 ();
 sg13g2_fill_1 FILLER_52_1898 ();
 sg13g2_fill_2 FILLER_52_1941 ();
 sg13g2_fill_2 FILLER_52_1983 ();
 sg13g2_fill_2 FILLER_52_1990 ();
 sg13g2_fill_1 FILLER_52_1992 ();
 sg13g2_fill_2 FILLER_52_2006 ();
 sg13g2_fill_1 FILLER_52_2029 ();
 sg13g2_fill_2 FILLER_52_2036 ();
 sg13g2_fill_1 FILLER_52_2038 ();
 sg13g2_fill_2 FILLER_52_2077 ();
 sg13g2_fill_1 FILLER_52_2079 ();
 sg13g2_fill_2 FILLER_52_2174 ();
 sg13g2_fill_1 FILLER_52_2176 ();
 sg13g2_fill_2 FILLER_52_2183 ();
 sg13g2_fill_1 FILLER_52_2203 ();
 sg13g2_fill_1 FILLER_52_2241 ();
 sg13g2_fill_2 FILLER_52_2269 ();
 sg13g2_decap_8 FILLER_52_2331 ();
 sg13g2_decap_8 FILLER_52_2338 ();
 sg13g2_decap_4 FILLER_52_2345 ();
 sg13g2_fill_2 FILLER_52_2358 ();
 sg13g2_fill_1 FILLER_52_2360 ();
 sg13g2_fill_1 FILLER_52_2385 ();
 sg13g2_decap_8 FILLER_52_2390 ();
 sg13g2_decap_8 FILLER_52_2397 ();
 sg13g2_decap_8 FILLER_52_2404 ();
 sg13g2_decap_8 FILLER_52_2411 ();
 sg13g2_decap_8 FILLER_52_2418 ();
 sg13g2_decap_8 FILLER_52_2425 ();
 sg13g2_decap_8 FILLER_52_2432 ();
 sg13g2_decap_8 FILLER_52_2439 ();
 sg13g2_decap_8 FILLER_52_2446 ();
 sg13g2_decap_8 FILLER_52_2453 ();
 sg13g2_decap_8 FILLER_52_2460 ();
 sg13g2_decap_8 FILLER_52_2467 ();
 sg13g2_decap_8 FILLER_52_2474 ();
 sg13g2_decap_8 FILLER_52_2481 ();
 sg13g2_decap_8 FILLER_52_2488 ();
 sg13g2_decap_8 FILLER_52_2495 ();
 sg13g2_decap_8 FILLER_52_2502 ();
 sg13g2_decap_8 FILLER_52_2509 ();
 sg13g2_decap_8 FILLER_52_2516 ();
 sg13g2_decap_8 FILLER_52_2523 ();
 sg13g2_decap_8 FILLER_52_2530 ();
 sg13g2_decap_8 FILLER_52_2537 ();
 sg13g2_decap_8 FILLER_52_2544 ();
 sg13g2_decap_8 FILLER_52_2551 ();
 sg13g2_decap_8 FILLER_52_2558 ();
 sg13g2_decap_8 FILLER_52_2565 ();
 sg13g2_decap_8 FILLER_52_2572 ();
 sg13g2_decap_8 FILLER_52_2579 ();
 sg13g2_decap_8 FILLER_52_2586 ();
 sg13g2_decap_8 FILLER_52_2593 ();
 sg13g2_decap_8 FILLER_52_2600 ();
 sg13g2_decap_8 FILLER_52_2607 ();
 sg13g2_decap_8 FILLER_52_2614 ();
 sg13g2_decap_8 FILLER_52_2621 ();
 sg13g2_decap_8 FILLER_52_2628 ();
 sg13g2_decap_8 FILLER_52_2635 ();
 sg13g2_decap_8 FILLER_52_2642 ();
 sg13g2_decap_8 FILLER_52_2649 ();
 sg13g2_decap_8 FILLER_52_2656 ();
 sg13g2_decap_8 FILLER_52_2663 ();
 sg13g2_decap_4 FILLER_52_2670 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_34 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_70 ();
 sg13g2_fill_1 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_123 ();
 sg13g2_fill_2 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_289 ();
 sg13g2_fill_2 FILLER_53_322 ();
 sg13g2_fill_1 FILLER_53_384 ();
 sg13g2_fill_2 FILLER_53_425 ();
 sg13g2_fill_2 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_440 ();
 sg13g2_decap_4 FILLER_53_446 ();
 sg13g2_fill_1 FILLER_53_450 ();
 sg13g2_fill_1 FILLER_53_468 ();
 sg13g2_fill_1 FILLER_53_495 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_fill_1 FILLER_53_545 ();
 sg13g2_decap_8 FILLER_53_559 ();
 sg13g2_decap_8 FILLER_53_566 ();
 sg13g2_fill_1 FILLER_53_573 ();
 sg13g2_decap_8 FILLER_53_622 ();
 sg13g2_decap_8 FILLER_53_629 ();
 sg13g2_decap_8 FILLER_53_636 ();
 sg13g2_decap_8 FILLER_53_643 ();
 sg13g2_decap_8 FILLER_53_650 ();
 sg13g2_decap_8 FILLER_53_657 ();
 sg13g2_fill_1 FILLER_53_690 ();
 sg13g2_decap_4 FILLER_53_704 ();
 sg13g2_fill_1 FILLER_53_708 ();
 sg13g2_fill_1 FILLER_53_718 ();
 sg13g2_decap_8 FILLER_53_730 ();
 sg13g2_fill_2 FILLER_53_737 ();
 sg13g2_fill_2 FILLER_53_776 ();
 sg13g2_fill_2 FILLER_53_863 ();
 sg13g2_fill_1 FILLER_53_874 ();
 sg13g2_decap_8 FILLER_53_889 ();
 sg13g2_fill_1 FILLER_53_896 ();
 sg13g2_fill_1 FILLER_53_948 ();
 sg13g2_decap_8 FILLER_53_987 ();
 sg13g2_decap_8 FILLER_53_994 ();
 sg13g2_fill_2 FILLER_53_1020 ();
 sg13g2_decap_4 FILLER_53_1060 ();
 sg13g2_decap_8 FILLER_53_1105 ();
 sg13g2_decap_4 FILLER_53_1112 ();
 sg13g2_fill_1 FILLER_53_1170 ();
 sg13g2_fill_1 FILLER_53_1180 ();
 sg13g2_fill_1 FILLER_53_1202 ();
 sg13g2_fill_1 FILLER_53_1227 ();
 sg13g2_decap_4 FILLER_53_1263 ();
 sg13g2_fill_1 FILLER_53_1330 ();
 sg13g2_fill_2 FILLER_53_1468 ();
 sg13g2_decap_4 FILLER_53_1497 ();
 sg13g2_fill_1 FILLER_53_1501 ();
 sg13g2_fill_2 FILLER_53_1540 ();
 sg13g2_fill_2 FILLER_53_1557 ();
 sg13g2_fill_1 FILLER_53_1559 ();
 sg13g2_fill_1 FILLER_53_1599 ();
 sg13g2_fill_2 FILLER_53_1664 ();
 sg13g2_fill_1 FILLER_53_1708 ();
 sg13g2_decap_4 FILLER_53_1743 ();
 sg13g2_fill_2 FILLER_53_1747 ();
 sg13g2_decap_8 FILLER_53_1786 ();
 sg13g2_decap_8 FILLER_53_1793 ();
 sg13g2_decap_4 FILLER_53_1800 ();
 sg13g2_fill_2 FILLER_53_1804 ();
 sg13g2_decap_8 FILLER_53_1836 ();
 sg13g2_decap_8 FILLER_53_1843 ();
 sg13g2_fill_1 FILLER_53_1850 ();
 sg13g2_fill_1 FILLER_53_1887 ();
 sg13g2_fill_2 FILLER_53_1933 ();
 sg13g2_fill_2 FILLER_53_1962 ();
 sg13g2_decap_8 FILLER_53_1989 ();
 sg13g2_fill_1 FILLER_53_2021 ();
 sg13g2_fill_2 FILLER_53_2042 ();
 sg13g2_fill_1 FILLER_53_2044 ();
 sg13g2_decap_4 FILLER_53_2057 ();
 sg13g2_fill_1 FILLER_53_2067 ();
 sg13g2_decap_4 FILLER_53_2133 ();
 sg13g2_fill_1 FILLER_53_2137 ();
 sg13g2_fill_1 FILLER_53_2168 ();
 sg13g2_fill_2 FILLER_53_2222 ();
 sg13g2_fill_1 FILLER_53_2291 ();
 sg13g2_decap_8 FILLER_53_2417 ();
 sg13g2_decap_8 FILLER_53_2424 ();
 sg13g2_decap_8 FILLER_53_2431 ();
 sg13g2_decap_8 FILLER_53_2438 ();
 sg13g2_decap_8 FILLER_53_2445 ();
 sg13g2_decap_8 FILLER_53_2452 ();
 sg13g2_decap_8 FILLER_53_2459 ();
 sg13g2_decap_8 FILLER_53_2466 ();
 sg13g2_decap_8 FILLER_53_2473 ();
 sg13g2_decap_8 FILLER_53_2480 ();
 sg13g2_decap_8 FILLER_53_2487 ();
 sg13g2_decap_8 FILLER_53_2494 ();
 sg13g2_decap_8 FILLER_53_2501 ();
 sg13g2_decap_8 FILLER_53_2508 ();
 sg13g2_decap_8 FILLER_53_2515 ();
 sg13g2_decap_8 FILLER_53_2522 ();
 sg13g2_decap_8 FILLER_53_2529 ();
 sg13g2_decap_8 FILLER_53_2536 ();
 sg13g2_decap_8 FILLER_53_2543 ();
 sg13g2_decap_8 FILLER_53_2550 ();
 sg13g2_decap_8 FILLER_53_2557 ();
 sg13g2_decap_8 FILLER_53_2564 ();
 sg13g2_decap_8 FILLER_53_2571 ();
 sg13g2_decap_8 FILLER_53_2578 ();
 sg13g2_decap_8 FILLER_53_2585 ();
 sg13g2_decap_8 FILLER_53_2592 ();
 sg13g2_decap_8 FILLER_53_2599 ();
 sg13g2_decap_8 FILLER_53_2606 ();
 sg13g2_decap_8 FILLER_53_2613 ();
 sg13g2_decap_8 FILLER_53_2620 ();
 sg13g2_decap_8 FILLER_53_2627 ();
 sg13g2_decap_8 FILLER_53_2634 ();
 sg13g2_decap_8 FILLER_53_2641 ();
 sg13g2_decap_8 FILLER_53_2648 ();
 sg13g2_decap_8 FILLER_53_2655 ();
 sg13g2_decap_8 FILLER_53_2662 ();
 sg13g2_decap_4 FILLER_53_2669 ();
 sg13g2_fill_1 FILLER_53_2673 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_fill_1 FILLER_54_37 ();
 sg13g2_fill_2 FILLER_54_47 ();
 sg13g2_fill_2 FILLER_54_68 ();
 sg13g2_fill_1 FILLER_54_90 ();
 sg13g2_fill_2 FILLER_54_118 ();
 sg13g2_fill_1 FILLER_54_120 ();
 sg13g2_fill_2 FILLER_54_188 ();
 sg13g2_fill_1 FILLER_54_249 ();
 sg13g2_fill_2 FILLER_54_254 ();
 sg13g2_fill_1 FILLER_54_332 ();
 sg13g2_decap_8 FILLER_54_355 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_fill_1 FILLER_54_411 ();
 sg13g2_fill_1 FILLER_54_466 ();
 sg13g2_fill_1 FILLER_54_512 ();
 sg13g2_decap_8 FILLER_54_545 ();
 sg13g2_decap_8 FILLER_54_552 ();
 sg13g2_decap_8 FILLER_54_559 ();
 sg13g2_decap_4 FILLER_54_566 ();
 sg13g2_fill_1 FILLER_54_570 ();
 sg13g2_fill_2 FILLER_54_604 ();
 sg13g2_decap_4 FILLER_54_703 ();
 sg13g2_fill_1 FILLER_54_707 ();
 sg13g2_fill_2 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_fill_2 FILLER_54_810 ();
 sg13g2_fill_2 FILLER_54_817 ();
 sg13g2_fill_1 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_892 ();
 sg13g2_decap_4 FILLER_54_899 ();
 sg13g2_fill_2 FILLER_54_903 ();
 sg13g2_decap_4 FILLER_54_918 ();
 sg13g2_fill_2 FILLER_54_999 ();
 sg13g2_fill_1 FILLER_54_1052 ();
 sg13g2_fill_2 FILLER_54_1057 ();
 sg13g2_decap_8 FILLER_54_1100 ();
 sg13g2_decap_8 FILLER_54_1107 ();
 sg13g2_fill_2 FILLER_54_1114 ();
 sg13g2_fill_1 FILLER_54_1116 ();
 sg13g2_fill_1 FILLER_54_1166 ();
 sg13g2_fill_2 FILLER_54_1286 ();
 sg13g2_fill_2 FILLER_54_1306 ();
 sg13g2_fill_2 FILLER_54_1325 ();
 sg13g2_fill_1 FILLER_54_1379 ();
 sg13g2_fill_2 FILLER_54_1393 ();
 sg13g2_fill_1 FILLER_54_1448 ();
 sg13g2_fill_2 FILLER_54_1462 ();
 sg13g2_fill_1 FILLER_54_1469 ();
 sg13g2_fill_2 FILLER_54_1483 ();
 sg13g2_decap_4 FILLER_54_1509 ();
 sg13g2_decap_8 FILLER_54_1530 ();
 sg13g2_decap_8 FILLER_54_1537 ();
 sg13g2_fill_2 FILLER_54_1583 ();
 sg13g2_fill_2 FILLER_54_1615 ();
 sg13g2_fill_2 FILLER_54_1663 ();
 sg13g2_fill_1 FILLER_54_1665 ();
 sg13g2_fill_2 FILLER_54_1679 ();
 sg13g2_fill_1 FILLER_54_1681 ();
 sg13g2_fill_2 FILLER_54_1686 ();
 sg13g2_fill_1 FILLER_54_1688 ();
 sg13g2_fill_2 FILLER_54_1778 ();
 sg13g2_fill_2 FILLER_54_1802 ();
 sg13g2_fill_1 FILLER_54_1804 ();
 sg13g2_fill_1 FILLER_54_1810 ();
 sg13g2_decap_8 FILLER_54_1834 ();
 sg13g2_decap_8 FILLER_54_1841 ();
 sg13g2_fill_2 FILLER_54_1848 ();
 sg13g2_fill_1 FILLER_54_1850 ();
 sg13g2_fill_2 FILLER_54_1867 ();
 sg13g2_fill_1 FILLER_54_1878 ();
 sg13g2_fill_2 FILLER_54_1926 ();
 sg13g2_fill_1 FILLER_54_1940 ();
 sg13g2_fill_1 FILLER_54_1958 ();
 sg13g2_fill_1 FILLER_54_1985 ();
 sg13g2_decap_8 FILLER_54_1999 ();
 sg13g2_decap_8 FILLER_54_2006 ();
 sg13g2_decap_4 FILLER_54_2013 ();
 sg13g2_decap_4 FILLER_54_2025 ();
 sg13g2_fill_2 FILLER_54_2029 ();
 sg13g2_fill_2 FILLER_54_2044 ();
 sg13g2_decap_4 FILLER_54_2052 ();
 sg13g2_fill_2 FILLER_54_2056 ();
 sg13g2_fill_2 FILLER_54_2082 ();
 sg13g2_fill_1 FILLER_54_2084 ();
 sg13g2_fill_2 FILLER_54_2091 ();
 sg13g2_fill_1 FILLER_54_2093 ();
 sg13g2_decap_4 FILLER_54_2132 ();
 sg13g2_fill_2 FILLER_54_2136 ();
 sg13g2_fill_2 FILLER_54_2143 ();
 sg13g2_fill_2 FILLER_54_2160 ();
 sg13g2_fill_1 FILLER_54_2162 ();
 sg13g2_fill_2 FILLER_54_2185 ();
 sg13g2_fill_1 FILLER_54_2375 ();
 sg13g2_decap_8 FILLER_54_2421 ();
 sg13g2_decap_8 FILLER_54_2428 ();
 sg13g2_decap_8 FILLER_54_2435 ();
 sg13g2_decap_8 FILLER_54_2442 ();
 sg13g2_decap_8 FILLER_54_2449 ();
 sg13g2_decap_8 FILLER_54_2456 ();
 sg13g2_decap_8 FILLER_54_2463 ();
 sg13g2_decap_8 FILLER_54_2470 ();
 sg13g2_decap_8 FILLER_54_2477 ();
 sg13g2_decap_8 FILLER_54_2484 ();
 sg13g2_decap_8 FILLER_54_2491 ();
 sg13g2_decap_8 FILLER_54_2498 ();
 sg13g2_decap_8 FILLER_54_2505 ();
 sg13g2_decap_8 FILLER_54_2512 ();
 sg13g2_decap_8 FILLER_54_2519 ();
 sg13g2_decap_8 FILLER_54_2526 ();
 sg13g2_decap_8 FILLER_54_2533 ();
 sg13g2_decap_8 FILLER_54_2540 ();
 sg13g2_decap_8 FILLER_54_2547 ();
 sg13g2_decap_8 FILLER_54_2554 ();
 sg13g2_decap_8 FILLER_54_2561 ();
 sg13g2_decap_8 FILLER_54_2568 ();
 sg13g2_decap_8 FILLER_54_2575 ();
 sg13g2_decap_8 FILLER_54_2582 ();
 sg13g2_decap_8 FILLER_54_2589 ();
 sg13g2_decap_8 FILLER_54_2596 ();
 sg13g2_decap_8 FILLER_54_2603 ();
 sg13g2_decap_8 FILLER_54_2610 ();
 sg13g2_decap_8 FILLER_54_2617 ();
 sg13g2_decap_8 FILLER_54_2624 ();
 sg13g2_decap_8 FILLER_54_2631 ();
 sg13g2_decap_8 FILLER_54_2638 ();
 sg13g2_decap_8 FILLER_54_2645 ();
 sg13g2_decap_8 FILLER_54_2652 ();
 sg13g2_decap_8 FILLER_54_2659 ();
 sg13g2_decap_8 FILLER_54_2666 ();
 sg13g2_fill_1 FILLER_54_2673 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_fill_2 FILLER_55_43 ();
 sg13g2_fill_1 FILLER_55_45 ();
 sg13g2_fill_2 FILLER_55_68 ();
 sg13g2_fill_1 FILLER_55_80 ();
 sg13g2_decap_4 FILLER_55_120 ();
 sg13g2_fill_1 FILLER_55_157 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_fill_2 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_272 ();
 sg13g2_fill_1 FILLER_55_274 ();
 sg13g2_fill_2 FILLER_55_288 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_decap_8 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_fill_1 FILLER_55_398 ();
 sg13g2_fill_1 FILLER_55_447 ();
 sg13g2_fill_1 FILLER_55_478 ();
 sg13g2_fill_2 FILLER_55_493 ();
 sg13g2_decap_8 FILLER_55_538 ();
 sg13g2_fill_2 FILLER_55_545 ();
 sg13g2_fill_1 FILLER_55_547 ();
 sg13g2_fill_2 FILLER_55_588 ();
 sg13g2_fill_1 FILLER_55_590 ();
 sg13g2_fill_2 FILLER_55_611 ();
 sg13g2_fill_1 FILLER_55_694 ();
 sg13g2_fill_2 FILLER_55_796 ();
 sg13g2_fill_1 FILLER_55_798 ();
 sg13g2_fill_1 FILLER_55_833 ();
 sg13g2_decap_4 FILLER_55_915 ();
 sg13g2_fill_1 FILLER_55_919 ();
 sg13g2_fill_2 FILLER_55_948 ();
 sg13g2_fill_1 FILLER_55_968 ();
 sg13g2_fill_2 FILLER_55_997 ();
 sg13g2_fill_1 FILLER_55_1037 ();
 sg13g2_fill_2 FILLER_55_1043 ();
 sg13g2_decap_4 FILLER_55_1049 ();
 sg13g2_fill_2 FILLER_55_1076 ();
 sg13g2_fill_1 FILLER_55_1078 ();
 sg13g2_decap_4 FILLER_55_1089 ();
 sg13g2_fill_1 FILLER_55_1121 ();
 sg13g2_decap_8 FILLER_55_1128 ();
 sg13g2_fill_1 FILLER_55_1135 ();
 sg13g2_fill_1 FILLER_55_1168 ();
 sg13g2_fill_1 FILLER_55_1188 ();
 sg13g2_fill_2 FILLER_55_1243 ();
 sg13g2_fill_1 FILLER_55_1245 ();
 sg13g2_fill_2 FILLER_55_1287 ();
 sg13g2_fill_1 FILLER_55_1370 ();
 sg13g2_fill_2 FILLER_55_1391 ();
 sg13g2_fill_1 FILLER_55_1393 ();
 sg13g2_fill_1 FILLER_55_1450 ();
 sg13g2_decap_8 FILLER_55_1457 ();
 sg13g2_fill_2 FILLER_55_1464 ();
 sg13g2_fill_1 FILLER_55_1499 ();
 sg13g2_fill_1 FILLER_55_1505 ();
 sg13g2_fill_2 FILLER_55_1551 ();
 sg13g2_fill_1 FILLER_55_1553 ();
 sg13g2_fill_2 FILLER_55_1575 ();
 sg13g2_fill_1 FILLER_55_1604 ();
 sg13g2_fill_2 FILLER_55_1642 ();
 sg13g2_fill_1 FILLER_55_1644 ();
 sg13g2_fill_1 FILLER_55_1688 ();
 sg13g2_fill_2 FILLER_55_1758 ();
 sg13g2_fill_1 FILLER_55_1773 ();
 sg13g2_fill_2 FILLER_55_1814 ();
 sg13g2_decap_4 FILLER_55_1841 ();
 sg13g2_fill_1 FILLER_55_1845 ();
 sg13g2_fill_1 FILLER_55_1864 ();
 sg13g2_fill_1 FILLER_55_2010 ();
 sg13g2_decap_4 FILLER_55_2042 ();
 sg13g2_fill_2 FILLER_55_2046 ();
 sg13g2_decap_8 FILLER_55_2052 ();
 sg13g2_fill_1 FILLER_55_2059 ();
 sg13g2_fill_2 FILLER_55_2091 ();
 sg13g2_fill_1 FILLER_55_2093 ();
 sg13g2_decap_4 FILLER_55_2105 ();
 sg13g2_fill_1 FILLER_55_2109 ();
 sg13g2_fill_2 FILLER_55_2151 ();
 sg13g2_fill_1 FILLER_55_2153 ();
 sg13g2_fill_2 FILLER_55_2162 ();
 sg13g2_fill_1 FILLER_55_2164 ();
 sg13g2_fill_2 FILLER_55_2170 ();
 sg13g2_fill_1 FILLER_55_2172 ();
 sg13g2_fill_2 FILLER_55_2190 ();
 sg13g2_fill_2 FILLER_55_2255 ();
 sg13g2_fill_1 FILLER_55_2257 ();
 sg13g2_fill_2 FILLER_55_2295 ();
 sg13g2_fill_1 FILLER_55_2297 ();
 sg13g2_fill_2 FILLER_55_2311 ();
 sg13g2_fill_1 FILLER_55_2313 ();
 sg13g2_fill_2 FILLER_55_2344 ();
 sg13g2_fill_2 FILLER_55_2373 ();
 sg13g2_fill_1 FILLER_55_2389 ();
 sg13g2_decap_8 FILLER_55_2430 ();
 sg13g2_decap_8 FILLER_55_2437 ();
 sg13g2_decap_8 FILLER_55_2444 ();
 sg13g2_decap_8 FILLER_55_2451 ();
 sg13g2_decap_8 FILLER_55_2458 ();
 sg13g2_decap_8 FILLER_55_2465 ();
 sg13g2_decap_8 FILLER_55_2472 ();
 sg13g2_decap_8 FILLER_55_2479 ();
 sg13g2_decap_8 FILLER_55_2486 ();
 sg13g2_decap_8 FILLER_55_2493 ();
 sg13g2_decap_8 FILLER_55_2500 ();
 sg13g2_decap_8 FILLER_55_2507 ();
 sg13g2_decap_8 FILLER_55_2514 ();
 sg13g2_decap_8 FILLER_55_2521 ();
 sg13g2_decap_8 FILLER_55_2528 ();
 sg13g2_decap_8 FILLER_55_2535 ();
 sg13g2_decap_8 FILLER_55_2542 ();
 sg13g2_decap_8 FILLER_55_2549 ();
 sg13g2_decap_8 FILLER_55_2556 ();
 sg13g2_decap_8 FILLER_55_2563 ();
 sg13g2_decap_8 FILLER_55_2570 ();
 sg13g2_decap_8 FILLER_55_2577 ();
 sg13g2_decap_8 FILLER_55_2584 ();
 sg13g2_decap_8 FILLER_55_2591 ();
 sg13g2_decap_8 FILLER_55_2598 ();
 sg13g2_decap_8 FILLER_55_2605 ();
 sg13g2_decap_8 FILLER_55_2612 ();
 sg13g2_decap_8 FILLER_55_2619 ();
 sg13g2_decap_8 FILLER_55_2626 ();
 sg13g2_decap_8 FILLER_55_2633 ();
 sg13g2_decap_8 FILLER_55_2640 ();
 sg13g2_decap_8 FILLER_55_2647 ();
 sg13g2_decap_8 FILLER_55_2654 ();
 sg13g2_decap_8 FILLER_55_2661 ();
 sg13g2_decap_4 FILLER_55_2668 ();
 sg13g2_fill_2 FILLER_55_2672 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_9 ();
 sg13g2_fill_2 FILLER_56_42 ();
 sg13g2_fill_1 FILLER_56_44 ();
 sg13g2_fill_2 FILLER_56_107 ();
 sg13g2_fill_1 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_fill_1 FILLER_56_121 ();
 sg13g2_fill_1 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_206 ();
 sg13g2_fill_2 FILLER_56_220 ();
 sg13g2_fill_1 FILLER_56_222 ();
 sg13g2_fill_1 FILLER_56_232 ();
 sg13g2_fill_1 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_332 ();
 sg13g2_fill_1 FILLER_56_339 ();
 sg13g2_fill_1 FILLER_56_345 ();
 sg13g2_decap_8 FILLER_56_363 ();
 sg13g2_fill_2 FILLER_56_387 ();
 sg13g2_fill_1 FILLER_56_389 ();
 sg13g2_fill_2 FILLER_56_399 ();
 sg13g2_fill_1 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_417 ();
 sg13g2_fill_2 FILLER_56_457 ();
 sg13g2_fill_1 FILLER_56_459 ();
 sg13g2_fill_2 FILLER_56_496 ();
 sg13g2_fill_2 FILLER_56_539 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_fill_2 FILLER_56_603 ();
 sg13g2_fill_1 FILLER_56_605 ();
 sg13g2_fill_2 FILLER_56_622 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_2 FILLER_56_709 ();
 sg13g2_fill_2 FILLER_56_718 ();
 sg13g2_fill_1 FILLER_56_720 ();
 sg13g2_fill_1 FILLER_56_737 ();
 sg13g2_fill_2 FILLER_56_791 ();
 sg13g2_fill_1 FILLER_56_793 ();
 sg13g2_fill_2 FILLER_56_821 ();
 sg13g2_fill_2 FILLER_56_888 ();
 sg13g2_fill_2 FILLER_56_912 ();
 sg13g2_fill_1 FILLER_56_914 ();
 sg13g2_fill_2 FILLER_56_959 ();
 sg13g2_fill_2 FILLER_56_977 ();
 sg13g2_decap_8 FILLER_56_1026 ();
 sg13g2_decap_8 FILLER_56_1033 ();
 sg13g2_decap_8 FILLER_56_1040 ();
 sg13g2_decap_8 FILLER_56_1047 ();
 sg13g2_fill_2 FILLER_56_1054 ();
 sg13g2_decap_4 FILLER_56_1083 ();
 sg13g2_decap_4 FILLER_56_1124 ();
 sg13g2_fill_2 FILLER_56_1128 ();
 sg13g2_fill_2 FILLER_56_1139 ();
 sg13g2_fill_2 FILLER_56_1176 ();
 sg13g2_fill_1 FILLER_56_1226 ();
 sg13g2_fill_2 FILLER_56_1259 ();
 sg13g2_fill_1 FILLER_56_1261 ();
 sg13g2_fill_2 FILLER_56_1294 ();
 sg13g2_fill_2 FILLER_56_1373 ();
 sg13g2_fill_1 FILLER_56_1375 ();
 sg13g2_fill_2 FILLER_56_1380 ();
 sg13g2_fill_1 FILLER_56_1409 ();
 sg13g2_fill_1 FILLER_56_1451 ();
 sg13g2_fill_2 FILLER_56_1466 ();
 sg13g2_fill_1 FILLER_56_1468 ();
 sg13g2_fill_2 FILLER_56_1480 ();
 sg13g2_fill_1 FILLER_56_1487 ();
 sg13g2_fill_2 FILLER_56_1493 ();
 sg13g2_fill_2 FILLER_56_1500 ();
 sg13g2_fill_2 FILLER_56_1529 ();
 sg13g2_fill_1 FILLER_56_1531 ();
 sg13g2_fill_1 FILLER_56_1563 ();
 sg13g2_decap_8 FILLER_56_1645 ();
 sg13g2_fill_1 FILLER_56_1652 ();
 sg13g2_fill_2 FILLER_56_1694 ();
 sg13g2_fill_1 FILLER_56_1732 ();
 sg13g2_fill_2 FILLER_56_1776 ();
 sg13g2_fill_2 FILLER_56_1803 ();
 sg13g2_fill_1 FILLER_56_1805 ();
 sg13g2_fill_1 FILLER_56_1896 ();
 sg13g2_decap_8 FILLER_56_1983 ();
 sg13g2_fill_1 FILLER_56_1990 ();
 sg13g2_fill_2 FILLER_56_2012 ();
 sg13g2_fill_1 FILLER_56_2014 ();
 sg13g2_fill_1 FILLER_56_2056 ();
 sg13g2_fill_2 FILLER_56_2094 ();
 sg13g2_fill_1 FILLER_56_2096 ();
 sg13g2_decap_8 FILLER_56_2125 ();
 sg13g2_decap_4 FILLER_56_2132 ();
 sg13g2_fill_1 FILLER_56_2145 ();
 sg13g2_fill_1 FILLER_56_2151 ();
 sg13g2_fill_2 FILLER_56_2179 ();
 sg13g2_fill_1 FILLER_56_2181 ();
 sg13g2_fill_2 FILLER_56_2200 ();
 sg13g2_fill_2 FILLER_56_2238 ();
 sg13g2_fill_1 FILLER_56_2240 ();
 sg13g2_decap_8 FILLER_56_2312 ();
 sg13g2_fill_2 FILLER_56_2319 ();
 sg13g2_fill_1 FILLER_56_2321 ();
 sg13g2_fill_1 FILLER_56_2326 ();
 sg13g2_fill_1 FILLER_56_2341 ();
 sg13g2_fill_1 FILLER_56_2351 ();
 sg13g2_fill_1 FILLER_56_2404 ();
 sg13g2_decap_8 FILLER_56_2422 ();
 sg13g2_decap_8 FILLER_56_2429 ();
 sg13g2_decap_8 FILLER_56_2436 ();
 sg13g2_decap_8 FILLER_56_2443 ();
 sg13g2_decap_8 FILLER_56_2450 ();
 sg13g2_decap_8 FILLER_56_2457 ();
 sg13g2_decap_8 FILLER_56_2464 ();
 sg13g2_decap_8 FILLER_56_2471 ();
 sg13g2_decap_8 FILLER_56_2478 ();
 sg13g2_decap_8 FILLER_56_2485 ();
 sg13g2_decap_8 FILLER_56_2492 ();
 sg13g2_decap_8 FILLER_56_2499 ();
 sg13g2_decap_8 FILLER_56_2506 ();
 sg13g2_decap_8 FILLER_56_2513 ();
 sg13g2_decap_8 FILLER_56_2520 ();
 sg13g2_decap_8 FILLER_56_2527 ();
 sg13g2_decap_8 FILLER_56_2534 ();
 sg13g2_decap_8 FILLER_56_2541 ();
 sg13g2_decap_8 FILLER_56_2548 ();
 sg13g2_decap_8 FILLER_56_2555 ();
 sg13g2_decap_8 FILLER_56_2562 ();
 sg13g2_decap_8 FILLER_56_2569 ();
 sg13g2_decap_8 FILLER_56_2576 ();
 sg13g2_decap_8 FILLER_56_2583 ();
 sg13g2_decap_8 FILLER_56_2590 ();
 sg13g2_decap_8 FILLER_56_2597 ();
 sg13g2_decap_8 FILLER_56_2604 ();
 sg13g2_decap_8 FILLER_56_2611 ();
 sg13g2_decap_8 FILLER_56_2618 ();
 sg13g2_decap_8 FILLER_56_2625 ();
 sg13g2_decap_8 FILLER_56_2632 ();
 sg13g2_decap_8 FILLER_56_2639 ();
 sg13g2_decap_8 FILLER_56_2646 ();
 sg13g2_decap_8 FILLER_56_2653 ();
 sg13g2_decap_8 FILLER_56_2660 ();
 sg13g2_decap_8 FILLER_56_2667 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_9 ();
 sg13g2_fill_2 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_120 ();
 sg13g2_fill_1 FILLER_57_199 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_decap_4 FILLER_57_229 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_fill_2 FILLER_57_286 ();
 sg13g2_fill_1 FILLER_57_288 ();
 sg13g2_decap_4 FILLER_57_329 ();
 sg13g2_fill_1 FILLER_57_333 ();
 sg13g2_fill_1 FILLER_57_343 ();
 sg13g2_fill_2 FILLER_57_385 ();
 sg13g2_fill_2 FILLER_57_396 ();
 sg13g2_fill_2 FILLER_57_411 ();
 sg13g2_decap_4 FILLER_57_435 ();
 sg13g2_fill_1 FILLER_57_439 ();
 sg13g2_fill_1 FILLER_57_459 ();
 sg13g2_fill_2 FILLER_57_505 ();
 sg13g2_fill_1 FILLER_57_507 ();
 sg13g2_fill_2 FILLER_57_543 ();
 sg13g2_fill_1 FILLER_57_623 ();
 sg13g2_fill_1 FILLER_57_661 ();
 sg13g2_fill_2 FILLER_57_719 ();
 sg13g2_fill_1 FILLER_57_721 ();
 sg13g2_fill_1 FILLER_57_731 ();
 sg13g2_fill_1 FILLER_57_842 ();
 sg13g2_fill_2 FILLER_57_861 ();
 sg13g2_fill_1 FILLER_57_863 ();
 sg13g2_fill_1 FILLER_57_891 ();
 sg13g2_fill_1 FILLER_57_943 ();
 sg13g2_decap_8 FILLER_57_1007 ();
 sg13g2_fill_1 FILLER_57_1014 ();
 sg13g2_decap_4 FILLER_57_1046 ();
 sg13g2_fill_2 FILLER_57_1070 ();
 sg13g2_fill_1 FILLER_57_1072 ();
 sg13g2_fill_2 FILLER_57_1082 ();
 sg13g2_decap_8 FILLER_57_1093 ();
 sg13g2_fill_2 FILLER_57_1100 ();
 sg13g2_fill_1 FILLER_57_1102 ();
 sg13g2_fill_1 FILLER_57_1131 ();
 sg13g2_fill_2 FILLER_57_1150 ();
 sg13g2_fill_2 FILLER_57_1218 ();
 sg13g2_fill_1 FILLER_57_1220 ();
 sg13g2_fill_2 FILLER_57_1251 ();
 sg13g2_fill_1 FILLER_57_1253 ();
 sg13g2_decap_4 FILLER_57_1264 ();
 sg13g2_fill_2 FILLER_57_1268 ();
 sg13g2_decap_8 FILLER_57_1361 ();
 sg13g2_fill_2 FILLER_57_1368 ();
 sg13g2_decap_4 FILLER_57_1375 ();
 sg13g2_fill_2 FILLER_57_1384 ();
 sg13g2_fill_1 FILLER_57_1395 ();
 sg13g2_decap_4 FILLER_57_1439 ();
 sg13g2_fill_2 FILLER_57_1487 ();
 sg13g2_fill_2 FILLER_57_1498 ();
 sg13g2_fill_2 FILLER_57_1519 ();
 sg13g2_fill_1 FILLER_57_1521 ();
 sg13g2_decap_8 FILLER_57_1531 ();
 sg13g2_decap_8 FILLER_57_1538 ();
 sg13g2_fill_2 FILLER_57_1545 ();
 sg13g2_fill_1 FILLER_57_1575 ();
 sg13g2_fill_1 FILLER_57_1589 ();
 sg13g2_fill_1 FILLER_57_1613 ();
 sg13g2_fill_2 FILLER_57_1713 ();
 sg13g2_decap_4 FILLER_57_1778 ();
 sg13g2_fill_1 FILLER_57_1782 ();
 sg13g2_fill_2 FILLER_57_1812 ();
 sg13g2_fill_1 FILLER_57_1843 ();
 sg13g2_fill_1 FILLER_57_1848 ();
 sg13g2_fill_2 FILLER_57_1888 ();
 sg13g2_fill_1 FILLER_57_1943 ();
 sg13g2_fill_1 FILLER_57_1962 ();
 sg13g2_decap_4 FILLER_57_1985 ();
 sg13g2_fill_2 FILLER_57_1989 ();
 sg13g2_fill_2 FILLER_57_2006 ();
 sg13g2_fill_1 FILLER_57_2032 ();
 sg13g2_decap_8 FILLER_57_2048 ();
 sg13g2_fill_2 FILLER_57_2055 ();
 sg13g2_fill_1 FILLER_57_2067 ();
 sg13g2_decap_8 FILLER_57_2084 ();
 sg13g2_decap_4 FILLER_57_2091 ();
 sg13g2_fill_2 FILLER_57_2095 ();
 sg13g2_fill_1 FILLER_57_2115 ();
 sg13g2_fill_1 FILLER_57_2134 ();
 sg13g2_fill_2 FILLER_57_2148 ();
 sg13g2_decap_4 FILLER_57_2163 ();
 sg13g2_fill_1 FILLER_57_2167 ();
 sg13g2_fill_2 FILLER_57_2238 ();
 sg13g2_decap_8 FILLER_57_2327 ();
 sg13g2_fill_2 FILLER_57_2334 ();
 sg13g2_fill_1 FILLER_57_2336 ();
 sg13g2_fill_1 FILLER_57_2363 ();
 sg13g2_fill_1 FILLER_57_2374 ();
 sg13g2_decap_8 FILLER_57_2426 ();
 sg13g2_decap_8 FILLER_57_2433 ();
 sg13g2_decap_8 FILLER_57_2440 ();
 sg13g2_decap_8 FILLER_57_2447 ();
 sg13g2_decap_8 FILLER_57_2454 ();
 sg13g2_decap_8 FILLER_57_2461 ();
 sg13g2_decap_8 FILLER_57_2468 ();
 sg13g2_decap_8 FILLER_57_2475 ();
 sg13g2_decap_8 FILLER_57_2482 ();
 sg13g2_decap_8 FILLER_57_2489 ();
 sg13g2_decap_8 FILLER_57_2496 ();
 sg13g2_decap_8 FILLER_57_2503 ();
 sg13g2_decap_8 FILLER_57_2510 ();
 sg13g2_decap_8 FILLER_57_2517 ();
 sg13g2_decap_8 FILLER_57_2524 ();
 sg13g2_decap_8 FILLER_57_2531 ();
 sg13g2_decap_8 FILLER_57_2538 ();
 sg13g2_decap_8 FILLER_57_2545 ();
 sg13g2_decap_8 FILLER_57_2552 ();
 sg13g2_decap_8 FILLER_57_2559 ();
 sg13g2_decap_8 FILLER_57_2566 ();
 sg13g2_decap_8 FILLER_57_2573 ();
 sg13g2_decap_8 FILLER_57_2580 ();
 sg13g2_decap_8 FILLER_57_2587 ();
 sg13g2_decap_8 FILLER_57_2594 ();
 sg13g2_decap_8 FILLER_57_2601 ();
 sg13g2_decap_8 FILLER_57_2608 ();
 sg13g2_decap_8 FILLER_57_2615 ();
 sg13g2_decap_8 FILLER_57_2622 ();
 sg13g2_decap_8 FILLER_57_2629 ();
 sg13g2_decap_8 FILLER_57_2636 ();
 sg13g2_decap_8 FILLER_57_2643 ();
 sg13g2_decap_8 FILLER_57_2650 ();
 sg13g2_decap_8 FILLER_57_2657 ();
 sg13g2_decap_8 FILLER_57_2664 ();
 sg13g2_fill_2 FILLER_57_2671 ();
 sg13g2_fill_1 FILLER_57_2673 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_105 ();
 sg13g2_fill_2 FILLER_58_109 ();
 sg13g2_decap_8 FILLER_58_124 ();
 sg13g2_fill_2 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_193 ();
 sg13g2_fill_2 FILLER_58_238 ();
 sg13g2_fill_2 FILLER_58_245 ();
 sg13g2_fill_1 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_395 ();
 sg13g2_fill_2 FILLER_58_460 ();
 sg13g2_fill_1 FILLER_58_462 ();
 sg13g2_decap_8 FILLER_58_495 ();
 sg13g2_decap_8 FILLER_58_502 ();
 sg13g2_decap_4 FILLER_58_509 ();
 sg13g2_fill_2 FILLER_58_513 ();
 sg13g2_decap_4 FILLER_58_520 ();
 sg13g2_fill_2 FILLER_58_524 ();
 sg13g2_fill_2 FILLER_58_539 ();
 sg13g2_fill_1 FILLER_58_541 ();
 sg13g2_fill_1 FILLER_58_545 ();
 sg13g2_fill_2 FILLER_58_598 ();
 sg13g2_fill_1 FILLER_58_600 ();
 sg13g2_fill_2 FILLER_58_652 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_fill_2 FILLER_58_750 ();
 sg13g2_fill_1 FILLER_58_806 ();
 sg13g2_fill_1 FILLER_58_857 ();
 sg13g2_fill_1 FILLER_58_876 ();
 sg13g2_fill_2 FILLER_58_886 ();
 sg13g2_fill_1 FILLER_58_904 ();
 sg13g2_fill_2 FILLER_58_923 ();
 sg13g2_decap_8 FILLER_58_931 ();
 sg13g2_decap_4 FILLER_58_938 ();
 sg13g2_fill_1 FILLER_58_942 ();
 sg13g2_decap_8 FILLER_58_946 ();
 sg13g2_fill_2 FILLER_58_953 ();
 sg13g2_fill_1 FILLER_58_955 ();
 sg13g2_decap_8 FILLER_58_969 ();
 sg13g2_fill_2 FILLER_58_989 ();
 sg13g2_decap_8 FILLER_58_997 ();
 sg13g2_decap_8 FILLER_58_1004 ();
 sg13g2_fill_2 FILLER_58_1011 ();
 sg13g2_decap_4 FILLER_58_1019 ();
 sg13g2_fill_2 FILLER_58_1023 ();
 sg13g2_fill_2 FILLER_58_1048 ();
 sg13g2_decap_4 FILLER_58_1087 ();
 sg13g2_fill_1 FILLER_58_1091 ();
 sg13g2_decap_8 FILLER_58_1105 ();
 sg13g2_decap_4 FILLER_58_1112 ();
 sg13g2_fill_1 FILLER_58_1198 ();
 sg13g2_fill_1 FILLER_58_1235 ();
 sg13g2_fill_2 FILLER_58_1277 ();
 sg13g2_fill_2 FILLER_58_1296 ();
 sg13g2_fill_1 FILLER_58_1308 ();
 sg13g2_fill_2 FILLER_58_1368 ();
 sg13g2_decap_4 FILLER_58_1375 ();
 sg13g2_fill_2 FILLER_58_1410 ();
 sg13g2_fill_1 FILLER_58_1412 ();
 sg13g2_fill_1 FILLER_58_1424 ();
 sg13g2_fill_2 FILLER_58_1467 ();
 sg13g2_fill_1 FILLER_58_1469 ();
 sg13g2_fill_2 FILLER_58_1488 ();
 sg13g2_fill_1 FILLER_58_1505 ();
 sg13g2_decap_8 FILLER_58_1531 ();
 sg13g2_decap_8 FILLER_58_1538 ();
 sg13g2_decap_8 FILLER_58_1545 ();
 sg13g2_fill_1 FILLER_58_1552 ();
 sg13g2_fill_2 FILLER_58_1558 ();
 sg13g2_fill_1 FILLER_58_1560 ();
 sg13g2_fill_1 FILLER_58_1574 ();
 sg13g2_decap_4 FILLER_58_1585 ();
 sg13g2_fill_2 FILLER_58_1597 ();
 sg13g2_fill_1 FILLER_58_1599 ();
 sg13g2_decap_8 FILLER_58_1645 ();
 sg13g2_fill_1 FILLER_58_1652 ();
 sg13g2_fill_2 FILLER_58_1730 ();
 sg13g2_fill_2 FILLER_58_1741 ();
 sg13g2_fill_2 FILLER_58_1781 ();
 sg13g2_fill_1 FILLER_58_1783 ();
 sg13g2_fill_1 FILLER_58_1797 ();
 sg13g2_fill_2 FILLER_58_1813 ();
 sg13g2_fill_2 FILLER_58_1839 ();
 sg13g2_fill_1 FILLER_58_1841 ();
 sg13g2_fill_1 FILLER_58_1923 ();
 sg13g2_fill_2 FILLER_58_1998 ();
 sg13g2_fill_2 FILLER_58_2008 ();
 sg13g2_fill_1 FILLER_58_2010 ();
 sg13g2_fill_1 FILLER_58_2037 ();
 sg13g2_fill_1 FILLER_58_2057 ();
 sg13g2_fill_2 FILLER_58_2071 ();
 sg13g2_fill_2 FILLER_58_2085 ();
 sg13g2_decap_8 FILLER_58_2166 ();
 sg13g2_decap_8 FILLER_58_2173 ();
 sg13g2_decap_4 FILLER_58_2180 ();
 sg13g2_fill_1 FILLER_58_2184 ();
 sg13g2_fill_2 FILLER_58_2198 ();
 sg13g2_fill_2 FILLER_58_2254 ();
 sg13g2_fill_2 FILLER_58_2340 ();
 sg13g2_fill_2 FILLER_58_2355 ();
 sg13g2_fill_1 FILLER_58_2370 ();
 sg13g2_decap_8 FILLER_58_2417 ();
 sg13g2_decap_8 FILLER_58_2424 ();
 sg13g2_decap_8 FILLER_58_2431 ();
 sg13g2_decap_8 FILLER_58_2438 ();
 sg13g2_decap_8 FILLER_58_2445 ();
 sg13g2_decap_8 FILLER_58_2452 ();
 sg13g2_decap_8 FILLER_58_2459 ();
 sg13g2_decap_8 FILLER_58_2466 ();
 sg13g2_decap_8 FILLER_58_2473 ();
 sg13g2_decap_8 FILLER_58_2480 ();
 sg13g2_decap_8 FILLER_58_2487 ();
 sg13g2_decap_8 FILLER_58_2494 ();
 sg13g2_decap_8 FILLER_58_2501 ();
 sg13g2_decap_8 FILLER_58_2508 ();
 sg13g2_decap_8 FILLER_58_2515 ();
 sg13g2_decap_8 FILLER_58_2522 ();
 sg13g2_decap_8 FILLER_58_2529 ();
 sg13g2_decap_8 FILLER_58_2536 ();
 sg13g2_decap_8 FILLER_58_2543 ();
 sg13g2_decap_8 FILLER_58_2550 ();
 sg13g2_decap_8 FILLER_58_2557 ();
 sg13g2_decap_8 FILLER_58_2564 ();
 sg13g2_decap_8 FILLER_58_2571 ();
 sg13g2_decap_8 FILLER_58_2578 ();
 sg13g2_decap_8 FILLER_58_2585 ();
 sg13g2_decap_8 FILLER_58_2592 ();
 sg13g2_decap_8 FILLER_58_2599 ();
 sg13g2_decap_8 FILLER_58_2606 ();
 sg13g2_decap_8 FILLER_58_2613 ();
 sg13g2_decap_8 FILLER_58_2620 ();
 sg13g2_decap_8 FILLER_58_2627 ();
 sg13g2_decap_8 FILLER_58_2634 ();
 sg13g2_decap_8 FILLER_58_2641 ();
 sg13g2_decap_8 FILLER_58_2648 ();
 sg13g2_decap_8 FILLER_58_2655 ();
 sg13g2_decap_8 FILLER_58_2662 ();
 sg13g2_decap_4 FILLER_58_2669 ();
 sg13g2_fill_1 FILLER_58_2673 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_43 ();
 sg13g2_fill_2 FILLER_59_58 ();
 sg13g2_fill_1 FILLER_59_60 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_1 FILLER_59_90 ();
 sg13g2_decap_8 FILLER_59_104 ();
 sg13g2_decap_8 FILLER_59_111 ();
 sg13g2_decap_4 FILLER_59_118 ();
 sg13g2_fill_1 FILLER_59_122 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_190 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_2 FILLER_59_274 ();
 sg13g2_fill_1 FILLER_59_276 ();
 sg13g2_fill_2 FILLER_59_290 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_fill_2 FILLER_59_362 ();
 sg13g2_fill_1 FILLER_59_387 ();
 sg13g2_fill_1 FILLER_59_459 ();
 sg13g2_fill_1 FILLER_59_474 ();
 sg13g2_decap_4 FILLER_59_501 ();
 sg13g2_decap_4 FILLER_59_532 ();
 sg13g2_fill_2 FILLER_59_561 ();
 sg13g2_fill_2 FILLER_59_596 ();
 sg13g2_fill_1 FILLER_59_598 ();
 sg13g2_fill_2 FILLER_59_632 ();
 sg13g2_fill_1 FILLER_59_742 ();
 sg13g2_fill_2 FILLER_59_820 ();
 sg13g2_fill_1 FILLER_59_822 ();
 sg13g2_fill_1 FILLER_59_837 ();
 sg13g2_fill_1 FILLER_59_882 ();
 sg13g2_decap_4 FILLER_59_897 ();
 sg13g2_decap_8 FILLER_59_910 ();
 sg13g2_decap_8 FILLER_59_920 ();
 sg13g2_decap_8 FILLER_59_927 ();
 sg13g2_decap_8 FILLER_59_934 ();
 sg13g2_decap_8 FILLER_59_941 ();
 sg13g2_decap_8 FILLER_59_948 ();
 sg13g2_decap_8 FILLER_59_955 ();
 sg13g2_decap_8 FILLER_59_962 ();
 sg13g2_decap_8 FILLER_59_969 ();
 sg13g2_decap_8 FILLER_59_993 ();
 sg13g2_decap_8 FILLER_59_1000 ();
 sg13g2_decap_4 FILLER_59_1007 ();
 sg13g2_fill_2 FILLER_59_1011 ();
 sg13g2_decap_4 FILLER_59_1026 ();
 sg13g2_fill_2 FILLER_59_1076 ();
 sg13g2_fill_2 FILLER_59_1106 ();
 sg13g2_fill_1 FILLER_59_1108 ();
 sg13g2_fill_1 FILLER_59_1179 ();
 sg13g2_fill_2 FILLER_59_1217 ();
 sg13g2_fill_1 FILLER_59_1251 ();
 sg13g2_fill_2 FILLER_59_1289 ();
 sg13g2_fill_1 FILLER_59_1331 ();
 sg13g2_fill_2 FILLER_59_1370 ();
 sg13g2_fill_1 FILLER_59_1372 ();
 sg13g2_decap_8 FILLER_59_1378 ();
 sg13g2_fill_2 FILLER_59_1385 ();
 sg13g2_fill_2 FILLER_59_1404 ();
 sg13g2_fill_1 FILLER_59_1406 ();
 sg13g2_fill_1 FILLER_59_1469 ();
 sg13g2_fill_1 FILLER_59_1535 ();
 sg13g2_fill_2 FILLER_59_1546 ();
 sg13g2_fill_1 FILLER_59_1554 ();
 sg13g2_fill_2 FILLER_59_1559 ();
 sg13g2_fill_1 FILLER_59_1561 ();
 sg13g2_decap_8 FILLER_59_1579 ();
 sg13g2_fill_1 FILLER_59_1586 ();
 sg13g2_fill_1 FILLER_59_1595 ();
 sg13g2_decap_8 FILLER_59_1627 ();
 sg13g2_fill_2 FILLER_59_1638 ();
 sg13g2_fill_1 FILLER_59_1640 ();
 sg13g2_fill_2 FILLER_59_1645 ();
 sg13g2_fill_1 FILLER_59_1647 ();
 sg13g2_decap_4 FILLER_59_1659 ();
 sg13g2_fill_1 FILLER_59_1680 ();
 sg13g2_fill_2 FILLER_59_1720 ();
 sg13g2_fill_1 FILLER_59_1759 ();
 sg13g2_fill_1 FILLER_59_1788 ();
 sg13g2_fill_2 FILLER_59_1802 ();
 sg13g2_fill_2 FILLER_59_1819 ();
 sg13g2_fill_1 FILLER_59_1895 ();
 sg13g2_fill_1 FILLER_59_1900 ();
 sg13g2_fill_2 FILLER_59_1912 ();
 sg13g2_fill_2 FILLER_59_1928 ();
 sg13g2_fill_1 FILLER_59_1996 ();
 sg13g2_fill_2 FILLER_59_2042 ();
 sg13g2_fill_1 FILLER_59_2044 ();
 sg13g2_decap_4 FILLER_59_2058 ();
 sg13g2_fill_1 FILLER_59_2072 ();
 sg13g2_fill_2 FILLER_59_2083 ();
 sg13g2_fill_2 FILLER_59_2113 ();
 sg13g2_fill_1 FILLER_59_2115 ();
 sg13g2_decap_4 FILLER_59_2149 ();
 sg13g2_fill_2 FILLER_59_2163 ();
 sg13g2_fill_2 FILLER_59_2187 ();
 sg13g2_fill_1 FILLER_59_2189 ();
 sg13g2_fill_2 FILLER_59_2208 ();
 sg13g2_fill_1 FILLER_59_2232 ();
 sg13g2_fill_2 FILLER_59_2242 ();
 sg13g2_fill_1 FILLER_59_2244 ();
 sg13g2_fill_2 FILLER_59_2288 ();
 sg13g2_decap_4 FILLER_59_2336 ();
 sg13g2_fill_2 FILLER_59_2340 ();
 sg13g2_fill_1 FILLER_59_2375 ();
 sg13g2_decap_8 FILLER_59_2416 ();
 sg13g2_decap_8 FILLER_59_2423 ();
 sg13g2_decap_8 FILLER_59_2430 ();
 sg13g2_decap_8 FILLER_59_2437 ();
 sg13g2_decap_8 FILLER_59_2444 ();
 sg13g2_decap_8 FILLER_59_2451 ();
 sg13g2_decap_8 FILLER_59_2458 ();
 sg13g2_decap_8 FILLER_59_2465 ();
 sg13g2_decap_8 FILLER_59_2472 ();
 sg13g2_decap_8 FILLER_59_2479 ();
 sg13g2_decap_8 FILLER_59_2486 ();
 sg13g2_decap_8 FILLER_59_2493 ();
 sg13g2_decap_8 FILLER_59_2500 ();
 sg13g2_decap_8 FILLER_59_2507 ();
 sg13g2_decap_8 FILLER_59_2514 ();
 sg13g2_decap_8 FILLER_59_2521 ();
 sg13g2_decap_8 FILLER_59_2528 ();
 sg13g2_decap_8 FILLER_59_2535 ();
 sg13g2_decap_8 FILLER_59_2542 ();
 sg13g2_decap_8 FILLER_59_2549 ();
 sg13g2_decap_8 FILLER_59_2556 ();
 sg13g2_decap_8 FILLER_59_2563 ();
 sg13g2_decap_8 FILLER_59_2570 ();
 sg13g2_decap_8 FILLER_59_2577 ();
 sg13g2_decap_8 FILLER_59_2584 ();
 sg13g2_decap_8 FILLER_59_2591 ();
 sg13g2_decap_8 FILLER_59_2598 ();
 sg13g2_decap_8 FILLER_59_2605 ();
 sg13g2_decap_8 FILLER_59_2612 ();
 sg13g2_decap_8 FILLER_59_2619 ();
 sg13g2_decap_8 FILLER_59_2626 ();
 sg13g2_decap_8 FILLER_59_2633 ();
 sg13g2_decap_8 FILLER_59_2640 ();
 sg13g2_decap_8 FILLER_59_2647 ();
 sg13g2_decap_8 FILLER_59_2654 ();
 sg13g2_decap_8 FILLER_59_2661 ();
 sg13g2_decap_4 FILLER_59_2668 ();
 sg13g2_fill_2 FILLER_59_2672 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_118 ();
 sg13g2_fill_2 FILLER_60_161 ();
 sg13g2_fill_1 FILLER_60_163 ();
 sg13g2_fill_2 FILLER_60_179 ();
 sg13g2_fill_1 FILLER_60_226 ();
 sg13g2_fill_1 FILLER_60_245 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_fill_2 FILLER_60_301 ();
 sg13g2_fill_2 FILLER_60_321 ();
 sg13g2_fill_1 FILLER_60_323 ();
 sg13g2_fill_2 FILLER_60_343 ();
 sg13g2_fill_1 FILLER_60_345 ();
 sg13g2_fill_2 FILLER_60_355 ();
 sg13g2_fill_1 FILLER_60_420 ();
 sg13g2_fill_1 FILLER_60_439 ();
 sg13g2_fill_1 FILLER_60_499 ();
 sg13g2_fill_2 FILLER_60_537 ();
 sg13g2_fill_1 FILLER_60_539 ();
 sg13g2_fill_2 FILLER_60_617 ();
 sg13g2_fill_1 FILLER_60_669 ();
 sg13g2_fill_2 FILLER_60_743 ();
 sg13g2_fill_1 FILLER_60_745 ();
 sg13g2_fill_2 FILLER_60_783 ();
 sg13g2_fill_2 FILLER_60_803 ();
 sg13g2_fill_2 FILLER_60_900 ();
 sg13g2_fill_1 FILLER_60_902 ();
 sg13g2_decap_8 FILLER_60_921 ();
 sg13g2_fill_2 FILLER_60_928 ();
 sg13g2_decap_4 FILLER_60_944 ();
 sg13g2_decap_8 FILLER_60_956 ();
 sg13g2_decap_4 FILLER_60_963 ();
 sg13g2_fill_1 FILLER_60_967 ();
 sg13g2_fill_2 FILLER_60_986 ();
 sg13g2_fill_1 FILLER_60_988 ();
 sg13g2_fill_2 FILLER_60_994 ();
 sg13g2_fill_2 FILLER_60_1007 ();
 sg13g2_fill_1 FILLER_60_1031 ();
 sg13g2_fill_2 FILLER_60_1037 ();
 sg13g2_fill_1 FILLER_60_1039 ();
 sg13g2_fill_2 FILLER_60_1059 ();
 sg13g2_fill_1 FILLER_60_1061 ();
 sg13g2_decap_4 FILLER_60_1090 ();
 sg13g2_fill_1 FILLER_60_1172 ();
 sg13g2_fill_1 FILLER_60_1216 ();
 sg13g2_fill_2 FILLER_60_1258 ();
 sg13g2_fill_1 FILLER_60_1260 ();
 sg13g2_fill_2 FILLER_60_1325 ();
 sg13g2_fill_1 FILLER_60_1327 ();
 sg13g2_fill_2 FILLER_60_1361 ();
 sg13g2_fill_1 FILLER_60_1363 ();
 sg13g2_fill_2 FILLER_60_1376 ();
 sg13g2_decap_4 FILLER_60_1403 ();
 sg13g2_fill_2 FILLER_60_1407 ();
 sg13g2_fill_2 FILLER_60_1445 ();
 sg13g2_decap_4 FILLER_60_1462 ();
 sg13g2_fill_2 FILLER_60_1484 ();
 sg13g2_fill_1 FILLER_60_1486 ();
 sg13g2_decap_8 FILLER_60_1584 ();
 sg13g2_decap_8 FILLER_60_1591 ();
 sg13g2_decap_8 FILLER_60_1622 ();
 sg13g2_fill_1 FILLER_60_1635 ();
 sg13g2_fill_1 FILLER_60_1706 ();
 sg13g2_fill_2 FILLER_60_1748 ();
 sg13g2_fill_1 FILLER_60_1750 ();
 sg13g2_fill_2 FILLER_60_1788 ();
 sg13g2_fill_1 FILLER_60_1790 ();
 sg13g2_fill_2 FILLER_60_1851 ();
 sg13g2_fill_1 FILLER_60_1870 ();
 sg13g2_fill_1 FILLER_60_1911 ();
 sg13g2_fill_2 FILLER_60_1928 ();
 sg13g2_fill_1 FILLER_60_1967 ();
 sg13g2_decap_4 FILLER_60_1995 ();
 sg13g2_fill_2 FILLER_60_1999 ();
 sg13g2_fill_2 FILLER_60_2051 ();
 sg13g2_fill_2 FILLER_60_2072 ();
 sg13g2_fill_1 FILLER_60_2082 ();
 sg13g2_fill_2 FILLER_60_2104 ();
 sg13g2_fill_2 FILLER_60_2155 ();
 sg13g2_fill_1 FILLER_60_2157 ();
 sg13g2_fill_2 FILLER_60_2186 ();
 sg13g2_fill_1 FILLER_60_2197 ();
 sg13g2_fill_1 FILLER_60_2203 ();
 sg13g2_fill_1 FILLER_60_2222 ();
 sg13g2_fill_2 FILLER_60_2251 ();
 sg13g2_fill_2 FILLER_60_2266 ();
 sg13g2_fill_1 FILLER_60_2268 ();
 sg13g2_fill_1 FILLER_60_2346 ();
 sg13g2_fill_2 FILLER_60_2351 ();
 sg13g2_fill_1 FILLER_60_2353 ();
 sg13g2_fill_1 FILLER_60_2387 ();
 sg13g2_decap_8 FILLER_60_2410 ();
 sg13g2_decap_8 FILLER_60_2417 ();
 sg13g2_decap_8 FILLER_60_2424 ();
 sg13g2_decap_8 FILLER_60_2431 ();
 sg13g2_decap_8 FILLER_60_2438 ();
 sg13g2_decap_8 FILLER_60_2445 ();
 sg13g2_decap_8 FILLER_60_2452 ();
 sg13g2_decap_8 FILLER_60_2459 ();
 sg13g2_decap_8 FILLER_60_2466 ();
 sg13g2_decap_8 FILLER_60_2473 ();
 sg13g2_decap_8 FILLER_60_2480 ();
 sg13g2_decap_8 FILLER_60_2487 ();
 sg13g2_decap_8 FILLER_60_2494 ();
 sg13g2_decap_8 FILLER_60_2501 ();
 sg13g2_decap_8 FILLER_60_2508 ();
 sg13g2_decap_8 FILLER_60_2515 ();
 sg13g2_decap_8 FILLER_60_2522 ();
 sg13g2_decap_8 FILLER_60_2529 ();
 sg13g2_decap_8 FILLER_60_2536 ();
 sg13g2_decap_8 FILLER_60_2543 ();
 sg13g2_decap_8 FILLER_60_2550 ();
 sg13g2_decap_8 FILLER_60_2557 ();
 sg13g2_decap_8 FILLER_60_2564 ();
 sg13g2_decap_8 FILLER_60_2571 ();
 sg13g2_decap_8 FILLER_60_2578 ();
 sg13g2_decap_8 FILLER_60_2585 ();
 sg13g2_decap_8 FILLER_60_2592 ();
 sg13g2_decap_8 FILLER_60_2599 ();
 sg13g2_decap_8 FILLER_60_2606 ();
 sg13g2_decap_8 FILLER_60_2613 ();
 sg13g2_decap_8 FILLER_60_2620 ();
 sg13g2_decap_8 FILLER_60_2627 ();
 sg13g2_decap_8 FILLER_60_2634 ();
 sg13g2_decap_8 FILLER_60_2641 ();
 sg13g2_decap_8 FILLER_60_2648 ();
 sg13g2_decap_8 FILLER_60_2655 ();
 sg13g2_decap_8 FILLER_60_2662 ();
 sg13g2_decap_4 FILLER_60_2669 ();
 sg13g2_fill_1 FILLER_60_2673 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_2 FILLER_61_43 ();
 sg13g2_fill_2 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_87 ();
 sg13g2_fill_2 FILLER_61_127 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_fill_2 FILLER_61_214 ();
 sg13g2_fill_1 FILLER_61_216 ();
 sg13g2_fill_2 FILLER_61_225 ();
 sg13g2_fill_1 FILLER_61_227 ();
 sg13g2_decap_8 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_241 ();
 sg13g2_fill_1 FILLER_61_273 ();
 sg13g2_fill_2 FILLER_61_283 ();
 sg13g2_fill_1 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_339 ();
 sg13g2_fill_2 FILLER_61_400 ();
 sg13g2_fill_2 FILLER_61_455 ();
 sg13g2_fill_1 FILLER_61_457 ();
 sg13g2_fill_2 FILLER_61_475 ();
 sg13g2_fill_1 FILLER_61_477 ();
 sg13g2_fill_2 FILLER_61_544 ();
 sg13g2_fill_1 FILLER_61_549 ();
 sg13g2_fill_2 FILLER_61_627 ();
 sg13g2_fill_1 FILLER_61_697 ();
 sg13g2_fill_2 FILLER_61_746 ();
 sg13g2_fill_1 FILLER_61_817 ();
 sg13g2_decap_8 FILLER_61_878 ();
 sg13g2_fill_1 FILLER_61_885 ();
 sg13g2_fill_2 FILLER_61_890 ();
 sg13g2_fill_1 FILLER_61_897 ();
 sg13g2_fill_1 FILLER_61_903 ();
 sg13g2_decap_8 FILLER_61_922 ();
 sg13g2_fill_2 FILLER_61_929 ();
 sg13g2_decap_4 FILLER_61_962 ();
 sg13g2_fill_1 FILLER_61_966 ();
 sg13g2_fill_2 FILLER_61_974 ();
 sg13g2_fill_2 FILLER_61_981 ();
 sg13g2_fill_2 FILLER_61_1043 ();
 sg13g2_fill_2 FILLER_61_1058 ();
 sg13g2_fill_1 FILLER_61_1060 ();
 sg13g2_fill_1 FILLER_61_1247 ();
 sg13g2_decap_4 FILLER_61_1330 ();
 sg13g2_decap_4 FILLER_61_1372 ();
 sg13g2_fill_2 FILLER_61_1380 ();
 sg13g2_fill_1 FILLER_61_1478 ();
 sg13g2_fill_2 FILLER_61_1525 ();
 sg13g2_fill_1 FILLER_61_1527 ();
 sg13g2_fill_2 FILLER_61_1537 ();
 sg13g2_fill_1 FILLER_61_1539 ();
 sg13g2_fill_1 FILLER_61_1554 ();
 sg13g2_decap_4 FILLER_61_1568 ();
 sg13g2_fill_2 FILLER_61_1572 ();
 sg13g2_decap_4 FILLER_61_1595 ();
 sg13g2_fill_1 FILLER_61_1599 ();
 sg13g2_fill_1 FILLER_61_1623 ();
 sg13g2_fill_1 FILLER_61_1670 ();
 sg13g2_decap_8 FILLER_61_1689 ();
 sg13g2_fill_1 FILLER_61_1696 ();
 sg13g2_fill_1 FILLER_61_1750 ();
 sg13g2_fill_2 FILLER_61_1836 ();
 sg13g2_fill_1 FILLER_61_1838 ();
 sg13g2_fill_1 FILLER_61_1861 ();
 sg13g2_fill_1 FILLER_61_1890 ();
 sg13g2_fill_2 FILLER_61_1896 ();
 sg13g2_fill_1 FILLER_61_1912 ();
 sg13g2_fill_1 FILLER_61_1921 ();
 sg13g2_fill_2 FILLER_61_1949 ();
 sg13g2_decap_8 FILLER_61_1999 ();
 sg13g2_decap_8 FILLER_61_2006 ();
 sg13g2_decap_4 FILLER_61_2017 ();
 sg13g2_decap_4 FILLER_61_2053 ();
 sg13g2_fill_1 FILLER_61_2057 ();
 sg13g2_fill_1 FILLER_61_2074 ();
 sg13g2_fill_1 FILLER_61_2109 ();
 sg13g2_fill_2 FILLER_61_2123 ();
 sg13g2_fill_1 FILLER_61_2182 ();
 sg13g2_fill_1 FILLER_61_2194 ();
 sg13g2_fill_1 FILLER_61_2209 ();
 sg13g2_fill_1 FILLER_61_2252 ();
 sg13g2_fill_1 FILLER_61_2282 ();
 sg13g2_fill_1 FILLER_61_2307 ();
 sg13g2_decap_4 FILLER_61_2349 ();
 sg13g2_fill_1 FILLER_61_2353 ();
 sg13g2_fill_2 FILLER_61_2362 ();
 sg13g2_fill_1 FILLER_61_2364 ();
 sg13g2_decap_8 FILLER_61_2401 ();
 sg13g2_decap_8 FILLER_61_2408 ();
 sg13g2_decap_8 FILLER_61_2415 ();
 sg13g2_decap_8 FILLER_61_2422 ();
 sg13g2_decap_8 FILLER_61_2429 ();
 sg13g2_decap_8 FILLER_61_2436 ();
 sg13g2_decap_8 FILLER_61_2443 ();
 sg13g2_decap_8 FILLER_61_2450 ();
 sg13g2_decap_8 FILLER_61_2457 ();
 sg13g2_decap_8 FILLER_61_2464 ();
 sg13g2_decap_8 FILLER_61_2471 ();
 sg13g2_decap_8 FILLER_61_2478 ();
 sg13g2_decap_8 FILLER_61_2485 ();
 sg13g2_decap_8 FILLER_61_2492 ();
 sg13g2_decap_8 FILLER_61_2499 ();
 sg13g2_decap_8 FILLER_61_2506 ();
 sg13g2_decap_8 FILLER_61_2513 ();
 sg13g2_decap_8 FILLER_61_2520 ();
 sg13g2_decap_8 FILLER_61_2527 ();
 sg13g2_decap_8 FILLER_61_2534 ();
 sg13g2_decap_8 FILLER_61_2541 ();
 sg13g2_decap_8 FILLER_61_2548 ();
 sg13g2_decap_8 FILLER_61_2555 ();
 sg13g2_decap_8 FILLER_61_2562 ();
 sg13g2_decap_8 FILLER_61_2569 ();
 sg13g2_decap_8 FILLER_61_2576 ();
 sg13g2_decap_8 FILLER_61_2583 ();
 sg13g2_decap_8 FILLER_61_2590 ();
 sg13g2_decap_8 FILLER_61_2597 ();
 sg13g2_decap_8 FILLER_61_2604 ();
 sg13g2_decap_8 FILLER_61_2611 ();
 sg13g2_decap_8 FILLER_61_2618 ();
 sg13g2_decap_8 FILLER_61_2625 ();
 sg13g2_decap_8 FILLER_61_2632 ();
 sg13g2_decap_8 FILLER_61_2639 ();
 sg13g2_decap_8 FILLER_61_2646 ();
 sg13g2_decap_8 FILLER_61_2653 ();
 sg13g2_decap_8 FILLER_61_2660 ();
 sg13g2_decap_8 FILLER_61_2667 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_fill_2 FILLER_62_39 ();
 sg13g2_fill_1 FILLER_62_50 ();
 sg13g2_decap_4 FILLER_62_81 ();
 sg13g2_fill_2 FILLER_62_121 ();
 sg13g2_fill_1 FILLER_62_123 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_decap_8 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_fill_2 FILLER_62_231 ();
 sg13g2_fill_1 FILLER_62_233 ();
 sg13g2_fill_2 FILLER_62_263 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_fill_2 FILLER_62_324 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_decap_8 FILLER_62_398 ();
 sg13g2_fill_1 FILLER_62_436 ();
 sg13g2_decap_4 FILLER_62_481 ();
 sg13g2_fill_2 FILLER_62_485 ();
 sg13g2_decap_8 FILLER_62_500 ();
 sg13g2_decap_4 FILLER_62_542 ();
 sg13g2_decap_4 FILLER_62_559 ();
 sg13g2_fill_2 FILLER_62_572 ();
 sg13g2_fill_1 FILLER_62_592 ();
 sg13g2_fill_1 FILLER_62_630 ();
 sg13g2_fill_1 FILLER_62_704 ();
 sg13g2_fill_1 FILLER_62_720 ();
 sg13g2_fill_2 FILLER_62_735 ();
 sg13g2_fill_2 FILLER_62_828 ();
 sg13g2_fill_1 FILLER_62_830 ();
 sg13g2_decap_8 FILLER_62_881 ();
 sg13g2_decap_8 FILLER_62_888 ();
 sg13g2_fill_2 FILLER_62_899 ();
 sg13g2_fill_1 FILLER_62_901 ();
 sg13g2_decap_8 FILLER_62_909 ();
 sg13g2_decap_8 FILLER_62_916 ();
 sg13g2_decap_8 FILLER_62_923 ();
 sg13g2_decap_4 FILLER_62_930 ();
 sg13g2_decap_8 FILLER_62_944 ();
 sg13g2_decap_4 FILLER_62_955 ();
 sg13g2_fill_1 FILLER_62_959 ();
 sg13g2_fill_2 FILLER_62_965 ();
 sg13g2_fill_1 FILLER_62_975 ();
 sg13g2_decap_8 FILLER_62_991 ();
 sg13g2_decap_8 FILLER_62_998 ();
 sg13g2_fill_1 FILLER_62_1005 ();
 sg13g2_decap_4 FILLER_62_1019 ();
 sg13g2_fill_1 FILLER_62_1023 ();
 sg13g2_decap_8 FILLER_62_1044 ();
 sg13g2_decap_8 FILLER_62_1051 ();
 sg13g2_decap_4 FILLER_62_1058 ();
 sg13g2_fill_2 FILLER_62_1062 ();
 sg13g2_fill_2 FILLER_62_1069 ();
 sg13g2_fill_1 FILLER_62_1071 ();
 sg13g2_fill_1 FILLER_62_1219 ();
 sg13g2_fill_2 FILLER_62_1262 ();
 sg13g2_fill_2 FILLER_62_1282 ();
 sg13g2_decap_8 FILLER_62_1377 ();
 sg13g2_decap_4 FILLER_62_1384 ();
 sg13g2_fill_1 FILLER_62_1388 ();
 sg13g2_decap_8 FILLER_62_1564 ();
 sg13g2_fill_1 FILLER_62_1571 ();
 sg13g2_fill_2 FILLER_62_1576 ();
 sg13g2_fill_1 FILLER_62_1578 ();
 sg13g2_fill_2 FILLER_62_1645 ();
 sg13g2_fill_2 FILLER_62_1662 ();
 sg13g2_fill_1 FILLER_62_1664 ();
 sg13g2_fill_2 FILLER_62_1706 ();
 sg13g2_fill_1 FILLER_62_1746 ();
 sg13g2_fill_1 FILLER_62_1798 ();
 sg13g2_fill_2 FILLER_62_1877 ();
 sg13g2_fill_2 FILLER_62_1911 ();
 sg13g2_fill_1 FILLER_62_1925 ();
 sg13g2_fill_2 FILLER_62_1984 ();
 sg13g2_fill_2 FILLER_62_2015 ();
 sg13g2_fill_2 FILLER_62_2038 ();
 sg13g2_fill_2 FILLER_62_2057 ();
 sg13g2_fill_2 FILLER_62_2073 ();
 sg13g2_fill_1 FILLER_62_2102 ();
 sg13g2_fill_1 FILLER_62_2120 ();
 sg13g2_fill_1 FILLER_62_2145 ();
 sg13g2_fill_1 FILLER_62_2159 ();
 sg13g2_fill_2 FILLER_62_2200 ();
 sg13g2_fill_1 FILLER_62_2217 ();
 sg13g2_fill_2 FILLER_62_2264 ();
 sg13g2_fill_1 FILLER_62_2279 ();
 sg13g2_fill_1 FILLER_62_2314 ();
 sg13g2_decap_4 FILLER_62_2337 ();
 sg13g2_fill_2 FILLER_62_2373 ();
 sg13g2_fill_2 FILLER_62_2379 ();
 sg13g2_fill_1 FILLER_62_2381 ();
 sg13g2_fill_1 FILLER_62_2395 ();
 sg13g2_decap_8 FILLER_62_2405 ();
 sg13g2_decap_8 FILLER_62_2412 ();
 sg13g2_decap_8 FILLER_62_2419 ();
 sg13g2_decap_8 FILLER_62_2426 ();
 sg13g2_decap_8 FILLER_62_2433 ();
 sg13g2_decap_8 FILLER_62_2440 ();
 sg13g2_decap_8 FILLER_62_2447 ();
 sg13g2_decap_8 FILLER_62_2454 ();
 sg13g2_decap_8 FILLER_62_2461 ();
 sg13g2_decap_8 FILLER_62_2468 ();
 sg13g2_decap_8 FILLER_62_2475 ();
 sg13g2_decap_8 FILLER_62_2482 ();
 sg13g2_decap_8 FILLER_62_2489 ();
 sg13g2_decap_8 FILLER_62_2496 ();
 sg13g2_decap_8 FILLER_62_2503 ();
 sg13g2_decap_8 FILLER_62_2510 ();
 sg13g2_decap_8 FILLER_62_2517 ();
 sg13g2_decap_8 FILLER_62_2524 ();
 sg13g2_decap_8 FILLER_62_2531 ();
 sg13g2_decap_8 FILLER_62_2538 ();
 sg13g2_decap_8 FILLER_62_2545 ();
 sg13g2_decap_8 FILLER_62_2552 ();
 sg13g2_decap_8 FILLER_62_2559 ();
 sg13g2_decap_8 FILLER_62_2566 ();
 sg13g2_decap_8 FILLER_62_2573 ();
 sg13g2_decap_8 FILLER_62_2580 ();
 sg13g2_decap_8 FILLER_62_2587 ();
 sg13g2_decap_8 FILLER_62_2594 ();
 sg13g2_decap_8 FILLER_62_2601 ();
 sg13g2_decap_8 FILLER_62_2608 ();
 sg13g2_decap_8 FILLER_62_2615 ();
 sg13g2_decap_8 FILLER_62_2622 ();
 sg13g2_decap_8 FILLER_62_2629 ();
 sg13g2_decap_8 FILLER_62_2636 ();
 sg13g2_decap_8 FILLER_62_2643 ();
 sg13g2_decap_8 FILLER_62_2650 ();
 sg13g2_decap_8 FILLER_62_2657 ();
 sg13g2_decap_8 FILLER_62_2664 ();
 sg13g2_fill_2 FILLER_62_2671 ();
 sg13g2_fill_1 FILLER_62_2673 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_123 ();
 sg13g2_fill_2 FILLER_63_128 ();
 sg13g2_fill_1 FILLER_63_130 ();
 sg13g2_fill_2 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_fill_2 FILLER_63_269 ();
 sg13g2_decap_4 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_2 FILLER_63_325 ();
 sg13g2_fill_1 FILLER_63_363 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_decap_8 FILLER_63_403 ();
 sg13g2_fill_1 FILLER_63_419 ();
 sg13g2_fill_2 FILLER_63_452 ();
 sg13g2_fill_1 FILLER_63_454 ();
 sg13g2_fill_2 FILLER_63_464 ();
 sg13g2_fill_2 FILLER_63_475 ();
 sg13g2_fill_1 FILLER_63_477 ();
 sg13g2_decap_8 FILLER_63_491 ();
 sg13g2_decap_8 FILLER_63_498 ();
 sg13g2_decap_4 FILLER_63_505 ();
 sg13g2_fill_2 FILLER_63_509 ();
 sg13g2_fill_2 FILLER_63_549 ();
 sg13g2_decap_4 FILLER_63_582 ();
 sg13g2_fill_2 FILLER_63_604 ();
 sg13g2_fill_2 FILLER_63_619 ();
 sg13g2_fill_2 FILLER_63_770 ();
 sg13g2_fill_1 FILLER_63_772 ();
 sg13g2_fill_2 FILLER_63_822 ();
 sg13g2_decap_8 FILLER_63_877 ();
 sg13g2_decap_8 FILLER_63_884 ();
 sg13g2_decap_8 FILLER_63_905 ();
 sg13g2_decap_8 FILLER_63_912 ();
 sg13g2_decap_8 FILLER_63_919 ();
 sg13g2_decap_8 FILLER_63_926 ();
 sg13g2_decap_8 FILLER_63_933 ();
 sg13g2_decap_8 FILLER_63_940 ();
 sg13g2_decap_8 FILLER_63_947 ();
 sg13g2_decap_8 FILLER_63_954 ();
 sg13g2_decap_8 FILLER_63_961 ();
 sg13g2_decap_8 FILLER_63_968 ();
 sg13g2_decap_8 FILLER_63_975 ();
 sg13g2_decap_4 FILLER_63_990 ();
 sg13g2_fill_1 FILLER_63_994 ();
 sg13g2_decap_4 FILLER_63_1001 ();
 sg13g2_decap_4 FILLER_63_1029 ();
 sg13g2_decap_8 FILLER_63_1037 ();
 sg13g2_decap_8 FILLER_63_1044 ();
 sg13g2_decap_8 FILLER_63_1051 ();
 sg13g2_fill_1 FILLER_63_1058 ();
 sg13g2_decap_8 FILLER_63_1073 ();
 sg13g2_decap_8 FILLER_63_1080 ();
 sg13g2_decap_4 FILLER_63_1087 ();
 sg13g2_fill_2 FILLER_63_1091 ();
 sg13g2_fill_2 FILLER_63_1098 ();
 sg13g2_fill_1 FILLER_63_1100 ();
 sg13g2_fill_1 FILLER_63_1117 ();
 sg13g2_fill_2 FILLER_63_1140 ();
 sg13g2_fill_2 FILLER_63_1169 ();
 sg13g2_fill_1 FILLER_63_1171 ();
 sg13g2_decap_4 FILLER_63_1213 ();
 sg13g2_fill_2 FILLER_63_1226 ();
 sg13g2_fill_1 FILLER_63_1228 ();
 sg13g2_fill_2 FILLER_63_1242 ();
 sg13g2_fill_1 FILLER_63_1286 ();
 sg13g2_decap_4 FILLER_63_1331 ();
 sg13g2_fill_1 FILLER_63_1386 ();
 sg13g2_fill_2 FILLER_63_1413 ();
 sg13g2_fill_1 FILLER_63_1462 ();
 sg13g2_fill_2 FILLER_63_1495 ();
 sg13g2_fill_2 FILLER_63_1501 ();
 sg13g2_decap_4 FILLER_63_1537 ();
 sg13g2_fill_1 FILLER_63_1557 ();
 sg13g2_decap_4 FILLER_63_1588 ();
 sg13g2_fill_2 FILLER_63_1613 ();
 sg13g2_fill_2 FILLER_63_1656 ();
 sg13g2_decap_4 FILLER_63_1714 ();
 sg13g2_fill_2 FILLER_63_1718 ();
 sg13g2_fill_2 FILLER_63_1765 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_fill_1 FILLER_63_1849 ();
 sg13g2_fill_1 FILLER_63_1876 ();
 sg13g2_fill_2 FILLER_63_1921 ();
 sg13g2_fill_2 FILLER_63_1955 ();
 sg13g2_fill_1 FILLER_63_1985 ();
 sg13g2_fill_2 FILLER_63_2008 ();
 sg13g2_fill_1 FILLER_63_2024 ();
 sg13g2_fill_2 FILLER_63_2095 ();
 sg13g2_fill_1 FILLER_63_2097 ();
 sg13g2_fill_2 FILLER_63_2112 ();
 sg13g2_fill_1 FILLER_63_2114 ();
 sg13g2_fill_2 FILLER_63_2155 ();
 sg13g2_decap_4 FILLER_63_2170 ();
 sg13g2_fill_2 FILLER_63_2219 ();
 sg13g2_fill_2 FILLER_63_2230 ();
 sg13g2_fill_2 FILLER_63_2279 ();
 sg13g2_fill_1 FILLER_63_2281 ();
 sg13g2_decap_8 FILLER_63_2336 ();
 sg13g2_decap_4 FILLER_63_2343 ();
 sg13g2_decap_8 FILLER_63_2424 ();
 sg13g2_decap_8 FILLER_63_2431 ();
 sg13g2_decap_8 FILLER_63_2438 ();
 sg13g2_decap_8 FILLER_63_2445 ();
 sg13g2_decap_8 FILLER_63_2452 ();
 sg13g2_decap_8 FILLER_63_2459 ();
 sg13g2_decap_8 FILLER_63_2466 ();
 sg13g2_decap_8 FILLER_63_2473 ();
 sg13g2_decap_8 FILLER_63_2480 ();
 sg13g2_decap_8 FILLER_63_2487 ();
 sg13g2_decap_8 FILLER_63_2494 ();
 sg13g2_decap_8 FILLER_63_2501 ();
 sg13g2_decap_8 FILLER_63_2508 ();
 sg13g2_decap_8 FILLER_63_2515 ();
 sg13g2_decap_8 FILLER_63_2522 ();
 sg13g2_decap_8 FILLER_63_2529 ();
 sg13g2_decap_8 FILLER_63_2536 ();
 sg13g2_decap_8 FILLER_63_2543 ();
 sg13g2_decap_8 FILLER_63_2550 ();
 sg13g2_decap_8 FILLER_63_2557 ();
 sg13g2_decap_8 FILLER_63_2564 ();
 sg13g2_decap_8 FILLER_63_2571 ();
 sg13g2_decap_8 FILLER_63_2578 ();
 sg13g2_decap_8 FILLER_63_2585 ();
 sg13g2_decap_8 FILLER_63_2592 ();
 sg13g2_decap_8 FILLER_63_2599 ();
 sg13g2_decap_8 FILLER_63_2606 ();
 sg13g2_decap_8 FILLER_63_2613 ();
 sg13g2_decap_8 FILLER_63_2620 ();
 sg13g2_decap_8 FILLER_63_2627 ();
 sg13g2_decap_8 FILLER_63_2634 ();
 sg13g2_decap_8 FILLER_63_2641 ();
 sg13g2_decap_8 FILLER_63_2648 ();
 sg13g2_decap_8 FILLER_63_2655 ();
 sg13g2_decap_8 FILLER_63_2662 ();
 sg13g2_decap_4 FILLER_63_2669 ();
 sg13g2_fill_1 FILLER_63_2673 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_2 FILLER_64_62 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_fill_1 FILLER_64_93 ();
 sg13g2_decap_4 FILLER_64_103 ();
 sg13g2_fill_2 FILLER_64_107 ();
 sg13g2_decap_8 FILLER_64_113 ();
 sg13g2_decap_8 FILLER_64_120 ();
 sg13g2_decap_8 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_171 ();
 sg13g2_decap_4 FILLER_64_204 ();
 sg13g2_fill_2 FILLER_64_208 ();
 sg13g2_decap_8 FILLER_64_286 ();
 sg13g2_fill_2 FILLER_64_293 ();
 sg13g2_fill_1 FILLER_64_328 ();
 sg13g2_fill_2 FILLER_64_361 ();
 sg13g2_fill_1 FILLER_64_377 ();
 sg13g2_decap_8 FILLER_64_387 ();
 sg13g2_decap_8 FILLER_64_394 ();
 sg13g2_decap_8 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_4 FILLER_64_419 ();
 sg13g2_fill_2 FILLER_64_525 ();
 sg13g2_fill_1 FILLER_64_537 ();
 sg13g2_decap_8 FILLER_64_576 ();
 sg13g2_decap_8 FILLER_64_583 ();
 sg13g2_decap_8 FILLER_64_590 ();
 sg13g2_fill_1 FILLER_64_597 ();
 sg13g2_fill_2 FILLER_64_699 ();
 sg13g2_fill_2 FILLER_64_777 ();
 sg13g2_fill_1 FILLER_64_818 ();
 sg13g2_fill_2 FILLER_64_828 ();
 sg13g2_decap_8 FILLER_64_866 ();
 sg13g2_decap_8 FILLER_64_873 ();
 sg13g2_decap_8 FILLER_64_880 ();
 sg13g2_decap_8 FILLER_64_887 ();
 sg13g2_fill_2 FILLER_64_894 ();
 sg13g2_fill_1 FILLER_64_896 ();
 sg13g2_fill_2 FILLER_64_902 ();
 sg13g2_fill_1 FILLER_64_904 ();
 sg13g2_fill_1 FILLER_64_914 ();
 sg13g2_decap_8 FILLER_64_920 ();
 sg13g2_fill_2 FILLER_64_932 ();
 sg13g2_decap_8 FILLER_64_940 ();
 sg13g2_decap_8 FILLER_64_952 ();
 sg13g2_fill_2 FILLER_64_959 ();
 sg13g2_fill_2 FILLER_64_966 ();
 sg13g2_fill_2 FILLER_64_994 ();
 sg13g2_fill_1 FILLER_64_996 ();
 sg13g2_decap_4 FILLER_64_1002 ();
 sg13g2_fill_2 FILLER_64_1006 ();
 sg13g2_fill_1 FILLER_64_1017 ();
 sg13g2_decap_4 FILLER_64_1025 ();
 sg13g2_decap_8 FILLER_64_1035 ();
 sg13g2_decap_8 FILLER_64_1042 ();
 sg13g2_decap_8 FILLER_64_1049 ();
 sg13g2_decap_4 FILLER_64_1056 ();
 sg13g2_decap_8 FILLER_64_1064 ();
 sg13g2_decap_8 FILLER_64_1071 ();
 sg13g2_decap_8 FILLER_64_1078 ();
 sg13g2_decap_8 FILLER_64_1085 ();
 sg13g2_fill_2 FILLER_64_1092 ();
 sg13g2_fill_1 FILLER_64_1094 ();
 sg13g2_fill_1 FILLER_64_1149 ();
 sg13g2_fill_1 FILLER_64_1163 ();
 sg13g2_fill_2 FILLER_64_1209 ();
 sg13g2_fill_1 FILLER_64_1264 ();
 sg13g2_fill_2 FILLER_64_1283 ();
 sg13g2_fill_1 FILLER_64_1285 ();
 sg13g2_fill_2 FILLER_64_1341 ();
 sg13g2_fill_1 FILLER_64_1343 ();
 sg13g2_fill_1 FILLER_64_1350 ();
 sg13g2_fill_1 FILLER_64_1407 ();
 sg13g2_fill_2 FILLER_64_1414 ();
 sg13g2_fill_1 FILLER_64_1452 ();
 sg13g2_decap_8 FILLER_64_1501 ();
 sg13g2_fill_2 FILLER_64_1508 ();
 sg13g2_fill_1 FILLER_64_1518 ();
 sg13g2_fill_1 FILLER_64_1544 ();
 sg13g2_fill_1 FILLER_64_1553 ();
 sg13g2_decap_4 FILLER_64_1565 ();
 sg13g2_fill_1 FILLER_64_1576 ();
 sg13g2_fill_2 FILLER_64_1609 ();
 sg13g2_fill_1 FILLER_64_1611 ();
 sg13g2_fill_2 FILLER_64_1638 ();
 sg13g2_fill_1 FILLER_64_1640 ();
 sg13g2_decap_4 FILLER_64_1706 ();
 sg13g2_fill_2 FILLER_64_1818 ();
 sg13g2_fill_2 FILLER_64_1847 ();
 sg13g2_fill_1 FILLER_64_1849 ();
 sg13g2_fill_2 FILLER_64_1876 ();
 sg13g2_fill_2 FILLER_64_1891 ();
 sg13g2_fill_1 FILLER_64_1958 ();
 sg13g2_fill_1 FILLER_64_2045 ();
 sg13g2_fill_1 FILLER_64_2161 ();
 sg13g2_decap_8 FILLER_64_2172 ();
 sg13g2_decap_4 FILLER_64_2179 ();
 sg13g2_fill_1 FILLER_64_2240 ();
 sg13g2_fill_2 FILLER_64_2250 ();
 sg13g2_fill_1 FILLER_64_2270 ();
 sg13g2_fill_2 FILLER_64_2324 ();
 sg13g2_fill_1 FILLER_64_2326 ();
 sg13g2_decap_4 FILLER_64_2341 ();
 sg13g2_fill_1 FILLER_64_2345 ();
 sg13g2_fill_2 FILLER_64_2350 ();
 sg13g2_fill_1 FILLER_64_2352 ();
 sg13g2_fill_2 FILLER_64_2379 ();
 sg13g2_fill_2 FILLER_64_2391 ();
 sg13g2_decap_8 FILLER_64_2430 ();
 sg13g2_decap_8 FILLER_64_2437 ();
 sg13g2_decap_8 FILLER_64_2444 ();
 sg13g2_decap_8 FILLER_64_2451 ();
 sg13g2_decap_8 FILLER_64_2458 ();
 sg13g2_decap_8 FILLER_64_2465 ();
 sg13g2_decap_8 FILLER_64_2472 ();
 sg13g2_decap_8 FILLER_64_2479 ();
 sg13g2_decap_8 FILLER_64_2486 ();
 sg13g2_decap_8 FILLER_64_2493 ();
 sg13g2_decap_8 FILLER_64_2500 ();
 sg13g2_decap_8 FILLER_64_2507 ();
 sg13g2_decap_8 FILLER_64_2514 ();
 sg13g2_decap_8 FILLER_64_2521 ();
 sg13g2_decap_8 FILLER_64_2528 ();
 sg13g2_decap_8 FILLER_64_2535 ();
 sg13g2_decap_8 FILLER_64_2542 ();
 sg13g2_decap_8 FILLER_64_2549 ();
 sg13g2_decap_8 FILLER_64_2556 ();
 sg13g2_decap_8 FILLER_64_2563 ();
 sg13g2_decap_8 FILLER_64_2570 ();
 sg13g2_decap_8 FILLER_64_2577 ();
 sg13g2_decap_8 FILLER_64_2584 ();
 sg13g2_decap_8 FILLER_64_2591 ();
 sg13g2_decap_8 FILLER_64_2598 ();
 sg13g2_decap_8 FILLER_64_2605 ();
 sg13g2_decap_8 FILLER_64_2612 ();
 sg13g2_decap_8 FILLER_64_2619 ();
 sg13g2_decap_8 FILLER_64_2626 ();
 sg13g2_decap_8 FILLER_64_2633 ();
 sg13g2_decap_8 FILLER_64_2640 ();
 sg13g2_decap_8 FILLER_64_2647 ();
 sg13g2_decap_8 FILLER_64_2654 ();
 sg13g2_decap_8 FILLER_64_2661 ();
 sg13g2_decap_4 FILLER_64_2668 ();
 sg13g2_fill_2 FILLER_64_2672 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_2 ();
 sg13g2_fill_1 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_97 ();
 sg13g2_fill_2 FILLER_65_104 ();
 sg13g2_fill_1 FILLER_65_106 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_fill_2 FILLER_65_229 ();
 sg13g2_decap_8 FILLER_65_253 ();
 sg13g2_decap_8 FILLER_65_260 ();
 sg13g2_decap_4 FILLER_65_267 ();
 sg13g2_decap_8 FILLER_65_284 ();
 sg13g2_decap_8 FILLER_65_291 ();
 sg13g2_decap_4 FILLER_65_298 ();
 sg13g2_fill_2 FILLER_65_302 ();
 sg13g2_fill_2 FILLER_65_322 ();
 sg13g2_fill_1 FILLER_65_324 ();
 sg13g2_decap_4 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_333 ();
 sg13g2_fill_2 FILLER_65_339 ();
 sg13g2_fill_2 FILLER_65_350 ();
 sg13g2_fill_1 FILLER_65_352 ();
 sg13g2_fill_2 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_367 ();
 sg13g2_decap_8 FILLER_65_374 ();
 sg13g2_decap_8 FILLER_65_381 ();
 sg13g2_decap_4 FILLER_65_388 ();
 sg13g2_fill_1 FILLER_65_392 ();
 sg13g2_decap_4 FILLER_65_397 ();
 sg13g2_fill_1 FILLER_65_401 ();
 sg13g2_fill_2 FILLER_65_420 ();
 sg13g2_fill_1 FILLER_65_430 ();
 sg13g2_fill_2 FILLER_65_448 ();
 sg13g2_decap_8 FILLER_65_453 ();
 sg13g2_fill_1 FILLER_65_460 ();
 sg13g2_decap_8 FILLER_65_465 ();
 sg13g2_decap_8 FILLER_65_472 ();
 sg13g2_decap_8 FILLER_65_479 ();
 sg13g2_fill_1 FILLER_65_532 ();
 sg13g2_fill_2 FILLER_65_586 ();
 sg13g2_fill_1 FILLER_65_588 ();
 sg13g2_fill_1 FILLER_65_597 ();
 sg13g2_decap_4 FILLER_65_602 ();
 sg13g2_fill_2 FILLER_65_673 ();
 sg13g2_fill_2 FILLER_65_713 ();
 sg13g2_fill_1 FILLER_65_765 ();
 sg13g2_fill_1 FILLER_65_794 ();
 sg13g2_fill_2 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_65_872 ();
 sg13g2_decap_8 FILLER_65_879 ();
 sg13g2_fill_2 FILLER_65_922 ();
 sg13g2_fill_1 FILLER_65_924 ();
 sg13g2_fill_1 FILLER_65_938 ();
 sg13g2_decap_4 FILLER_65_970 ();
 sg13g2_fill_2 FILLER_65_1017 ();
 sg13g2_fill_1 FILLER_65_1019 ();
 sg13g2_fill_2 FILLER_65_1033 ();
 sg13g2_fill_1 FILLER_65_1035 ();
 sg13g2_decap_8 FILLER_65_1041 ();
 sg13g2_decap_4 FILLER_65_1048 ();
 sg13g2_fill_1 FILLER_65_1052 ();
 sg13g2_fill_2 FILLER_65_1071 ();
 sg13g2_decap_8 FILLER_65_1081 ();
 sg13g2_fill_2 FILLER_65_1088 ();
 sg13g2_fill_1 FILLER_65_1090 ();
 sg13g2_fill_2 FILLER_65_1138 ();
 sg13g2_fill_2 FILLER_65_1207 ();
 sg13g2_fill_1 FILLER_65_1209 ();
 sg13g2_decap_8 FILLER_65_1307 ();
 sg13g2_decap_8 FILLER_65_1318 ();
 sg13g2_decap_8 FILLER_65_1325 ();
 sg13g2_decap_4 FILLER_65_1332 ();
 sg13g2_fill_2 FILLER_65_1336 ();
 sg13g2_decap_8 FILLER_65_1343 ();
 sg13g2_decap_8 FILLER_65_1350 ();
 sg13g2_fill_2 FILLER_65_1357 ();
 sg13g2_fill_1 FILLER_65_1377 ();
 sg13g2_fill_2 FILLER_65_1452 ();
 sg13g2_fill_2 FILLER_65_1473 ();
 sg13g2_fill_2 FILLER_65_1499 ();
 sg13g2_fill_1 FILLER_65_1501 ();
 sg13g2_fill_1 FILLER_65_1525 ();
 sg13g2_fill_2 FILLER_65_1534 ();
 sg13g2_fill_1 FILLER_65_1536 ();
 sg13g2_fill_1 FILLER_65_1559 ();
 sg13g2_fill_2 FILLER_65_1594 ();
 sg13g2_fill_1 FILLER_65_1596 ();
 sg13g2_fill_2 FILLER_65_1648 ();
 sg13g2_fill_1 FILLER_65_1650 ();
 sg13g2_fill_1 FILLER_65_1669 ();
 sg13g2_fill_2 FILLER_65_1679 ();
 sg13g2_fill_1 FILLER_65_1681 ();
 sg13g2_fill_2 FILLER_65_1691 ();
 sg13g2_fill_1 FILLER_65_1693 ();
 sg13g2_fill_2 FILLER_65_1699 ();
 sg13g2_fill_1 FILLER_65_1701 ();
 sg13g2_fill_1 FILLER_65_1707 ();
 sg13g2_fill_2 FILLER_65_1739 ();
 sg13g2_fill_2 FILLER_65_1786 ();
 sg13g2_fill_2 FILLER_65_1847 ();
 sg13g2_fill_1 FILLER_65_1908 ();
 sg13g2_fill_2 FILLER_65_1986 ();
 sg13g2_fill_1 FILLER_65_2020 ();
 sg13g2_decap_8 FILLER_65_2032 ();
 sg13g2_fill_2 FILLER_65_2039 ();
 sg13g2_fill_1 FILLER_65_2041 ();
 sg13g2_fill_2 FILLER_65_2092 ();
 sg13g2_fill_1 FILLER_65_2094 ();
 sg13g2_fill_2 FILLER_65_2150 ();
 sg13g2_fill_1 FILLER_65_2179 ();
 sg13g2_fill_2 FILLER_65_2187 ();
 sg13g2_fill_1 FILLER_65_2189 ();
 sg13g2_fill_1 FILLER_65_2226 ();
 sg13g2_fill_1 FILLER_65_2258 ();
 sg13g2_fill_2 FILLER_65_2296 ();
 sg13g2_fill_1 FILLER_65_2308 ();
 sg13g2_fill_1 FILLER_65_2354 ();
 sg13g2_decap_8 FILLER_65_2438 ();
 sg13g2_decap_8 FILLER_65_2445 ();
 sg13g2_decap_8 FILLER_65_2452 ();
 sg13g2_decap_8 FILLER_65_2459 ();
 sg13g2_decap_8 FILLER_65_2466 ();
 sg13g2_decap_8 FILLER_65_2473 ();
 sg13g2_decap_8 FILLER_65_2480 ();
 sg13g2_decap_8 FILLER_65_2487 ();
 sg13g2_decap_8 FILLER_65_2494 ();
 sg13g2_decap_8 FILLER_65_2501 ();
 sg13g2_decap_8 FILLER_65_2508 ();
 sg13g2_decap_8 FILLER_65_2515 ();
 sg13g2_decap_8 FILLER_65_2522 ();
 sg13g2_decap_8 FILLER_65_2529 ();
 sg13g2_decap_8 FILLER_65_2536 ();
 sg13g2_decap_8 FILLER_65_2543 ();
 sg13g2_decap_8 FILLER_65_2550 ();
 sg13g2_decap_8 FILLER_65_2557 ();
 sg13g2_decap_8 FILLER_65_2564 ();
 sg13g2_decap_8 FILLER_65_2571 ();
 sg13g2_decap_8 FILLER_65_2578 ();
 sg13g2_decap_8 FILLER_65_2585 ();
 sg13g2_decap_8 FILLER_65_2592 ();
 sg13g2_decap_8 FILLER_65_2599 ();
 sg13g2_decap_8 FILLER_65_2606 ();
 sg13g2_decap_8 FILLER_65_2613 ();
 sg13g2_decap_8 FILLER_65_2620 ();
 sg13g2_decap_8 FILLER_65_2627 ();
 sg13g2_decap_8 FILLER_65_2634 ();
 sg13g2_decap_8 FILLER_65_2641 ();
 sg13g2_decap_8 FILLER_65_2648 ();
 sg13g2_decap_8 FILLER_65_2655 ();
 sg13g2_decap_8 FILLER_65_2662 ();
 sg13g2_decap_4 FILLER_65_2669 ();
 sg13g2_fill_1 FILLER_65_2673 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_fill_1 FILLER_66_46 ();
 sg13g2_decap_8 FILLER_66_90 ();
 sg13g2_decap_8 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_2 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_219 ();
 sg13g2_decap_4 FILLER_66_226 ();
 sg13g2_fill_1 FILLER_66_230 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_4 FILLER_66_266 ();
 sg13g2_fill_1 FILLER_66_270 ();
 sg13g2_fill_2 FILLER_66_288 ();
 sg13g2_fill_2 FILLER_66_296 ();
 sg13g2_decap_8 FILLER_66_304 ();
 sg13g2_decap_8 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_323 ();
 sg13g2_fill_2 FILLER_66_328 ();
 sg13g2_fill_2 FILLER_66_343 ();
 sg13g2_fill_1 FILLER_66_345 ();
 sg13g2_fill_1 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_376 ();
 sg13g2_fill_1 FILLER_66_383 ();
 sg13g2_fill_1 FILLER_66_416 ();
 sg13g2_decap_4 FILLER_66_449 ();
 sg13g2_fill_1 FILLER_66_453 ();
 sg13g2_decap_8 FILLER_66_482 ();
 sg13g2_fill_1 FILLER_66_493 ();
 sg13g2_fill_2 FILLER_66_543 ();
 sg13g2_fill_1 FILLER_66_545 ();
 sg13g2_fill_2 FILLER_66_555 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_fill_2 FILLER_66_696 ();
 sg13g2_fill_1 FILLER_66_760 ();
 sg13g2_fill_2 FILLER_66_765 ();
 sg13g2_fill_1 FILLER_66_767 ();
 sg13g2_fill_1 FILLER_66_794 ();
 sg13g2_fill_2 FILLER_66_856 ();
 sg13g2_fill_1 FILLER_66_884 ();
 sg13g2_fill_2 FILLER_66_904 ();
 sg13g2_fill_2 FILLER_66_931 ();
 sg13g2_decap_8 FILLER_66_987 ();
 sg13g2_fill_1 FILLER_66_994 ();
 sg13g2_fill_2 FILLER_66_1010 ();
 sg13g2_fill_2 FILLER_66_1017 ();
 sg13g2_fill_1 FILLER_66_1019 ();
 sg13g2_fill_1 FILLER_66_1026 ();
 sg13g2_fill_2 FILLER_66_1043 ();
 sg13g2_fill_1 FILLER_66_1045 ();
 sg13g2_decap_8 FILLER_66_1051 ();
 sg13g2_decap_8 FILLER_66_1058 ();
 sg13g2_fill_2 FILLER_66_1065 ();
 sg13g2_fill_1 FILLER_66_1080 ();
 sg13g2_fill_2 FILLER_66_1141 ();
 sg13g2_fill_1 FILLER_66_1143 ();
 sg13g2_fill_2 FILLER_66_1202 ();
 sg13g2_fill_1 FILLER_66_1204 ();
 sg13g2_fill_1 FILLER_66_1237 ();
 sg13g2_fill_1 FILLER_66_1260 ();
 sg13g2_decap_8 FILLER_66_1298 ();
 sg13g2_fill_1 FILLER_66_1305 ();
 sg13g2_decap_8 FILLER_66_1326 ();
 sg13g2_decap_8 FILLER_66_1333 ();
 sg13g2_decap_4 FILLER_66_1340 ();
 sg13g2_fill_2 FILLER_66_1352 ();
 sg13g2_fill_2 FILLER_66_1391 ();
 sg13g2_fill_1 FILLER_66_1406 ();
 sg13g2_fill_2 FILLER_66_1466 ();
 sg13g2_fill_1 FILLER_66_1468 ();
 sg13g2_fill_2 FILLER_66_1495 ();
 sg13g2_fill_2 FILLER_66_1539 ();
 sg13g2_fill_1 FILLER_66_1541 ();
 sg13g2_fill_1 FILLER_66_1566 ();
 sg13g2_fill_2 FILLER_66_1622 ();
 sg13g2_fill_1 FILLER_66_1624 ();
 sg13g2_fill_2 FILLER_66_1739 ();
 sg13g2_fill_2 FILLER_66_1799 ();
 sg13g2_fill_1 FILLER_66_1801 ();
 sg13g2_fill_2 FILLER_66_1847 ();
 sg13g2_fill_2 FILLER_66_1876 ();
 sg13g2_fill_1 FILLER_66_1940 ();
 sg13g2_fill_1 FILLER_66_1949 ();
 sg13g2_fill_2 FILLER_66_1964 ();
 sg13g2_fill_2 FILLER_66_1994 ();
 sg13g2_fill_2 FILLER_66_2005 ();
 sg13g2_fill_1 FILLER_66_2007 ();
 sg13g2_decap_8 FILLER_66_2028 ();
 sg13g2_decap_4 FILLER_66_2035 ();
 sg13g2_fill_1 FILLER_66_2058 ();
 sg13g2_fill_1 FILLER_66_2123 ();
 sg13g2_fill_2 FILLER_66_2151 ();
 sg13g2_fill_2 FILLER_66_2180 ();
 sg13g2_decap_4 FILLER_66_2298 ();
 sg13g2_fill_2 FILLER_66_2302 ();
 sg13g2_fill_2 FILLER_66_2313 ();
 sg13g2_fill_1 FILLER_66_2315 ();
 sg13g2_fill_2 FILLER_66_2351 ();
 sg13g2_fill_1 FILLER_66_2353 ();
 sg13g2_fill_2 FILLER_66_2368 ();
 sg13g2_decap_8 FILLER_66_2431 ();
 sg13g2_decap_8 FILLER_66_2438 ();
 sg13g2_decap_8 FILLER_66_2445 ();
 sg13g2_decap_8 FILLER_66_2452 ();
 sg13g2_decap_8 FILLER_66_2459 ();
 sg13g2_decap_8 FILLER_66_2466 ();
 sg13g2_decap_8 FILLER_66_2473 ();
 sg13g2_decap_8 FILLER_66_2480 ();
 sg13g2_decap_8 FILLER_66_2487 ();
 sg13g2_decap_8 FILLER_66_2494 ();
 sg13g2_decap_8 FILLER_66_2501 ();
 sg13g2_decap_8 FILLER_66_2508 ();
 sg13g2_decap_8 FILLER_66_2515 ();
 sg13g2_decap_8 FILLER_66_2522 ();
 sg13g2_decap_8 FILLER_66_2529 ();
 sg13g2_decap_8 FILLER_66_2536 ();
 sg13g2_decap_8 FILLER_66_2543 ();
 sg13g2_decap_8 FILLER_66_2550 ();
 sg13g2_decap_8 FILLER_66_2557 ();
 sg13g2_decap_8 FILLER_66_2564 ();
 sg13g2_decap_8 FILLER_66_2571 ();
 sg13g2_decap_8 FILLER_66_2578 ();
 sg13g2_decap_8 FILLER_66_2585 ();
 sg13g2_decap_8 FILLER_66_2592 ();
 sg13g2_decap_8 FILLER_66_2599 ();
 sg13g2_decap_8 FILLER_66_2606 ();
 sg13g2_decap_8 FILLER_66_2613 ();
 sg13g2_decap_8 FILLER_66_2620 ();
 sg13g2_decap_8 FILLER_66_2627 ();
 sg13g2_decap_8 FILLER_66_2634 ();
 sg13g2_decap_8 FILLER_66_2641 ();
 sg13g2_decap_8 FILLER_66_2648 ();
 sg13g2_decap_8 FILLER_66_2655 ();
 sg13g2_decap_8 FILLER_66_2662 ();
 sg13g2_decap_4 FILLER_66_2669 ();
 sg13g2_fill_1 FILLER_66_2673 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_1 FILLER_67_79 ();
 sg13g2_decap_4 FILLER_67_90 ();
 sg13g2_fill_1 FILLER_67_99 ();
 sg13g2_fill_2 FILLER_67_152 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_fill_1 FILLER_67_174 ();
 sg13g2_fill_2 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_349 ();
 sg13g2_fill_2 FILLER_67_404 ();
 sg13g2_decap_8 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_446 ();
 sg13g2_fill_2 FILLER_67_453 ();
 sg13g2_fill_1 FILLER_67_526 ();
 sg13g2_fill_1 FILLER_67_536 ();
 sg13g2_fill_2 FILLER_67_569 ();
 sg13g2_fill_2 FILLER_67_598 ();
 sg13g2_fill_1 FILLER_67_600 ();
 sg13g2_fill_1 FILLER_67_647 ();
 sg13g2_fill_2 FILLER_67_744 ();
 sg13g2_decap_8 FILLER_67_860 ();
 sg13g2_decap_8 FILLER_67_867 ();
 sg13g2_decap_4 FILLER_67_874 ();
 sg13g2_fill_2 FILLER_67_878 ();
 sg13g2_decap_8 FILLER_67_895 ();
 sg13g2_decap_4 FILLER_67_902 ();
 sg13g2_fill_1 FILLER_67_906 ();
 sg13g2_fill_1 FILLER_67_911 ();
 sg13g2_fill_2 FILLER_67_926 ();
 sg13g2_decap_8 FILLER_67_933 ();
 sg13g2_decap_4 FILLER_67_940 ();
 sg13g2_fill_2 FILLER_67_944 ();
 sg13g2_fill_2 FILLER_67_951 ();
 sg13g2_fill_1 FILLER_67_953 ();
 sg13g2_fill_2 FILLER_67_959 ();
 sg13g2_fill_1 FILLER_67_961 ();
 sg13g2_decap_8 FILLER_67_966 ();
 sg13g2_fill_2 FILLER_67_973 ();
 sg13g2_fill_1 FILLER_67_975 ();
 sg13g2_decap_4 FILLER_67_981 ();
 sg13g2_fill_2 FILLER_67_985 ();
 sg13g2_decap_8 FILLER_67_993 ();
 sg13g2_fill_2 FILLER_67_1000 ();
 sg13g2_decap_8 FILLER_67_1017 ();
 sg13g2_fill_2 FILLER_67_1024 ();
 sg13g2_fill_2 FILLER_67_1030 ();
 sg13g2_fill_1 FILLER_67_1050 ();
 sg13g2_decap_8 FILLER_67_1059 ();
 sg13g2_decap_8 FILLER_67_1066 ();
 sg13g2_fill_2 FILLER_67_1073 ();
 sg13g2_decap_8 FILLER_67_1084 ();
 sg13g2_decap_4 FILLER_67_1091 ();
 sg13g2_decap_4 FILLER_67_1108 ();
 sg13g2_decap_8 FILLER_67_1291 ();
 sg13g2_fill_2 FILLER_67_1298 ();
 sg13g2_fill_2 FILLER_67_1341 ();
 sg13g2_fill_1 FILLER_67_1343 ();
 sg13g2_fill_2 FILLER_67_1423 ();
 sg13g2_fill_1 FILLER_67_1502 ();
 sg13g2_fill_2 FILLER_67_1511 ();
 sg13g2_fill_1 FILLER_67_1513 ();
 sg13g2_fill_1 FILLER_67_1520 ();
 sg13g2_fill_1 FILLER_67_1565 ();
 sg13g2_decap_4 FILLER_67_1588 ();
 sg13g2_fill_1 FILLER_67_1592 ();
 sg13g2_decap_4 FILLER_67_1597 ();
 sg13g2_fill_1 FILLER_67_1651 ();
 sg13g2_fill_2 FILLER_67_1697 ();
 sg13g2_fill_1 FILLER_67_1744 ();
 sg13g2_fill_2 FILLER_67_1816 ();
 sg13g2_fill_2 FILLER_67_1930 ();
 sg13g2_fill_1 FILLER_67_1963 ();
 sg13g2_fill_1 FILLER_67_1978 ();
 sg13g2_fill_2 FILLER_67_2032 ();
 sg13g2_fill_2 FILLER_67_2038 ();
 sg13g2_fill_2 FILLER_67_2061 ();
 sg13g2_fill_1 FILLER_67_2072 ();
 sg13g2_fill_1 FILLER_67_2109 ();
 sg13g2_decap_8 FILLER_67_2146 ();
 sg13g2_decap_4 FILLER_67_2153 ();
 sg13g2_fill_1 FILLER_67_2157 ();
 sg13g2_decap_4 FILLER_67_2309 ();
 sg13g2_fill_2 FILLER_67_2313 ();
 sg13g2_fill_2 FILLER_67_2402 ();
 sg13g2_decap_8 FILLER_67_2422 ();
 sg13g2_decap_8 FILLER_67_2429 ();
 sg13g2_decap_8 FILLER_67_2436 ();
 sg13g2_decap_8 FILLER_67_2443 ();
 sg13g2_decap_8 FILLER_67_2450 ();
 sg13g2_decap_8 FILLER_67_2457 ();
 sg13g2_decap_8 FILLER_67_2464 ();
 sg13g2_decap_8 FILLER_67_2471 ();
 sg13g2_decap_8 FILLER_67_2478 ();
 sg13g2_decap_8 FILLER_67_2485 ();
 sg13g2_decap_8 FILLER_67_2492 ();
 sg13g2_decap_8 FILLER_67_2499 ();
 sg13g2_decap_8 FILLER_67_2506 ();
 sg13g2_decap_8 FILLER_67_2513 ();
 sg13g2_decap_8 FILLER_67_2520 ();
 sg13g2_decap_8 FILLER_67_2527 ();
 sg13g2_decap_8 FILLER_67_2534 ();
 sg13g2_decap_8 FILLER_67_2541 ();
 sg13g2_decap_8 FILLER_67_2548 ();
 sg13g2_decap_8 FILLER_67_2555 ();
 sg13g2_decap_8 FILLER_67_2562 ();
 sg13g2_decap_8 FILLER_67_2569 ();
 sg13g2_decap_8 FILLER_67_2576 ();
 sg13g2_decap_8 FILLER_67_2583 ();
 sg13g2_decap_8 FILLER_67_2590 ();
 sg13g2_decap_8 FILLER_67_2597 ();
 sg13g2_decap_8 FILLER_67_2604 ();
 sg13g2_decap_8 FILLER_67_2611 ();
 sg13g2_decap_8 FILLER_67_2618 ();
 sg13g2_decap_8 FILLER_67_2625 ();
 sg13g2_decap_8 FILLER_67_2632 ();
 sg13g2_decap_8 FILLER_67_2639 ();
 sg13g2_decap_8 FILLER_67_2646 ();
 sg13g2_decap_8 FILLER_67_2653 ();
 sg13g2_decap_8 FILLER_67_2660 ();
 sg13g2_decap_8 FILLER_67_2667 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_1 FILLER_68_52 ();
 sg13g2_decap_4 FILLER_68_78 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_305 ();
 sg13g2_fill_1 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_decap_4 FILLER_68_407 ();
 sg13g2_fill_1 FILLER_68_411 ();
 sg13g2_decap_8 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_4 FILLER_68_453 ();
 sg13g2_fill_1 FILLER_68_457 ();
 sg13g2_fill_1 FILLER_68_574 ();
 sg13g2_fill_1 FILLER_68_588 ();
 sg13g2_fill_2 FILLER_68_603 ();
 sg13g2_fill_1 FILLER_68_605 ();
 sg13g2_fill_2 FILLER_68_634 ();
 sg13g2_fill_1 FILLER_68_636 ();
 sg13g2_decap_8 FILLER_68_641 ();
 sg13g2_fill_1 FILLER_68_653 ();
 sg13g2_fill_2 FILLER_68_722 ();
 sg13g2_fill_1 FILLER_68_746 ();
 sg13g2_fill_1 FILLER_68_775 ();
 sg13g2_fill_1 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_878 ();
 sg13g2_decap_8 FILLER_68_885 ();
 sg13g2_decap_8 FILLER_68_892 ();
 sg13g2_decap_8 FILLER_68_899 ();
 sg13g2_decap_8 FILLER_68_906 ();
 sg13g2_decap_8 FILLER_68_913 ();
 sg13g2_decap_4 FILLER_68_920 ();
 sg13g2_fill_1 FILLER_68_924 ();
 sg13g2_decap_8 FILLER_68_941 ();
 sg13g2_decap_8 FILLER_68_948 ();
 sg13g2_fill_1 FILLER_68_955 ();
 sg13g2_decap_8 FILLER_68_962 ();
 sg13g2_decap_8 FILLER_68_969 ();
 sg13g2_decap_8 FILLER_68_976 ();
 sg13g2_decap_8 FILLER_68_983 ();
 sg13g2_decap_8 FILLER_68_990 ();
 sg13g2_decap_8 FILLER_68_997 ();
 sg13g2_decap_8 FILLER_68_1004 ();
 sg13g2_decap_8 FILLER_68_1011 ();
 sg13g2_decap_8 FILLER_68_1018 ();
 sg13g2_decap_8 FILLER_68_1025 ();
 sg13g2_decap_8 FILLER_68_1032 ();
 sg13g2_decap_8 FILLER_68_1039 ();
 sg13g2_decap_8 FILLER_68_1046 ();
 sg13g2_decap_4 FILLER_68_1053 ();
 sg13g2_fill_2 FILLER_68_1057 ();
 sg13g2_decap_4 FILLER_68_1076 ();
 sg13g2_fill_2 FILLER_68_1080 ();
 sg13g2_decap_8 FILLER_68_1095 ();
 sg13g2_decap_8 FILLER_68_1115 ();
 sg13g2_fill_1 FILLER_68_1122 ();
 sg13g2_fill_2 FILLER_68_1132 ();
 sg13g2_fill_1 FILLER_68_1175 ();
 sg13g2_fill_2 FILLER_68_1185 ();
 sg13g2_fill_1 FILLER_68_1205 ();
 sg13g2_fill_1 FILLER_68_1225 ();
 sg13g2_fill_2 FILLER_68_1293 ();
 sg13g2_fill_2 FILLER_68_1317 ();
 sg13g2_fill_1 FILLER_68_1368 ();
 sg13g2_decap_4 FILLER_68_1402 ();
 sg13g2_fill_2 FILLER_68_1436 ();
 sg13g2_fill_2 FILLER_68_1495 ();
 sg13g2_fill_1 FILLER_68_1497 ();
 sg13g2_fill_2 FILLER_68_1503 ();
 sg13g2_decap_8 FILLER_68_1514 ();
 sg13g2_decap_8 FILLER_68_1521 ();
 sg13g2_decap_8 FILLER_68_1528 ();
 sg13g2_fill_1 FILLER_68_1535 ();
 sg13g2_decap_8 FILLER_68_1562 ();
 sg13g2_fill_2 FILLER_68_1569 ();
 sg13g2_decap_8 FILLER_68_1599 ();
 sg13g2_fill_1 FILLER_68_1606 ();
 sg13g2_fill_2 FILLER_68_1677 ();
 sg13g2_fill_1 FILLER_68_1743 ();
 sg13g2_fill_2 FILLER_68_1939 ();
 sg13g2_fill_1 FILLER_68_1954 ();
 sg13g2_fill_2 FILLER_68_2000 ();
 sg13g2_fill_2 FILLER_68_2039 ();
 sg13g2_fill_2 FILLER_68_2119 ();
 sg13g2_decap_8 FILLER_68_2140 ();
 sg13g2_decap_8 FILLER_68_2147 ();
 sg13g2_decap_8 FILLER_68_2154 ();
 sg13g2_fill_2 FILLER_68_2161 ();
 sg13g2_fill_1 FILLER_68_2163 ();
 sg13g2_fill_2 FILLER_68_2218 ();
 sg13g2_decap_8 FILLER_68_2260 ();
 sg13g2_decap_8 FILLER_68_2272 ();
 sg13g2_decap_8 FILLER_68_2279 ();
 sg13g2_fill_2 FILLER_68_2286 ();
 sg13g2_fill_1 FILLER_68_2288 ();
 sg13g2_fill_1 FILLER_68_2299 ();
 sg13g2_fill_1 FILLER_68_2354 ();
 sg13g2_fill_2 FILLER_68_2360 ();
 sg13g2_fill_1 FILLER_68_2362 ();
 sg13g2_fill_1 FILLER_68_2368 ();
 sg13g2_fill_2 FILLER_68_2388 ();
 sg13g2_decap_8 FILLER_68_2416 ();
 sg13g2_decap_8 FILLER_68_2423 ();
 sg13g2_decap_8 FILLER_68_2430 ();
 sg13g2_decap_8 FILLER_68_2437 ();
 sg13g2_decap_8 FILLER_68_2444 ();
 sg13g2_decap_8 FILLER_68_2451 ();
 sg13g2_decap_8 FILLER_68_2458 ();
 sg13g2_decap_8 FILLER_68_2465 ();
 sg13g2_decap_8 FILLER_68_2472 ();
 sg13g2_decap_8 FILLER_68_2479 ();
 sg13g2_decap_8 FILLER_68_2486 ();
 sg13g2_decap_8 FILLER_68_2493 ();
 sg13g2_decap_8 FILLER_68_2500 ();
 sg13g2_decap_8 FILLER_68_2507 ();
 sg13g2_decap_8 FILLER_68_2514 ();
 sg13g2_decap_8 FILLER_68_2521 ();
 sg13g2_decap_8 FILLER_68_2528 ();
 sg13g2_decap_8 FILLER_68_2535 ();
 sg13g2_decap_8 FILLER_68_2542 ();
 sg13g2_decap_8 FILLER_68_2549 ();
 sg13g2_decap_8 FILLER_68_2556 ();
 sg13g2_decap_8 FILLER_68_2563 ();
 sg13g2_decap_8 FILLER_68_2570 ();
 sg13g2_decap_8 FILLER_68_2577 ();
 sg13g2_decap_8 FILLER_68_2584 ();
 sg13g2_decap_8 FILLER_68_2591 ();
 sg13g2_decap_8 FILLER_68_2598 ();
 sg13g2_decap_8 FILLER_68_2605 ();
 sg13g2_decap_8 FILLER_68_2612 ();
 sg13g2_decap_8 FILLER_68_2619 ();
 sg13g2_decap_8 FILLER_68_2626 ();
 sg13g2_decap_8 FILLER_68_2633 ();
 sg13g2_decap_8 FILLER_68_2640 ();
 sg13g2_decap_8 FILLER_68_2647 ();
 sg13g2_decap_8 FILLER_68_2654 ();
 sg13g2_decap_8 FILLER_68_2661 ();
 sg13g2_decap_4 FILLER_68_2668 ();
 sg13g2_fill_2 FILLER_68_2672 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_50 ();
 sg13g2_fill_1 FILLER_69_52 ();
 sg13g2_decap_8 FILLER_69_87 ();
 sg13g2_fill_2 FILLER_69_94 ();
 sg13g2_fill_2 FILLER_69_115 ();
 sg13g2_decap_4 FILLER_69_128 ();
 sg13g2_fill_2 FILLER_69_168 ();
 sg13g2_fill_1 FILLER_69_170 ();
 sg13g2_decap_8 FILLER_69_232 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_fill_1 FILLER_69_283 ();
 sg13g2_decap_8 FILLER_69_313 ();
 sg13g2_fill_1 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_352 ();
 sg13g2_decap_4 FILLER_69_384 ();
 sg13g2_fill_2 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_438 ();
 sg13g2_fill_2 FILLER_69_445 ();
 sg13g2_fill_1 FILLER_69_488 ();
 sg13g2_fill_1 FILLER_69_566 ();
 sg13g2_fill_2 FILLER_69_612 ();
 sg13g2_fill_2 FILLER_69_632 ();
 sg13g2_fill_2 FILLER_69_647 ();
 sg13g2_fill_2 FILLER_69_708 ();
 sg13g2_fill_2 FILLER_69_725 ();
 sg13g2_fill_1 FILLER_69_727 ();
 sg13g2_fill_2 FILLER_69_743 ();
 sg13g2_fill_1 FILLER_69_745 ();
 sg13g2_fill_1 FILLER_69_764 ();
 sg13g2_fill_2 FILLER_69_784 ();
 sg13g2_fill_1 FILLER_69_786 ();
 sg13g2_fill_2 FILLER_69_817 ();
 sg13g2_decap_4 FILLER_69_854 ();
 sg13g2_fill_2 FILLER_69_858 ();
 sg13g2_decap_4 FILLER_69_865 ();
 sg13g2_fill_1 FILLER_69_869 ();
 sg13g2_fill_2 FILLER_69_879 ();
 sg13g2_decap_8 FILLER_69_890 ();
 sg13g2_fill_2 FILLER_69_897 ();
 sg13g2_fill_1 FILLER_69_899 ();
 sg13g2_decap_8 FILLER_69_905 ();
 sg13g2_decap_8 FILLER_69_924 ();
 sg13g2_decap_8 FILLER_69_931 ();
 sg13g2_decap_8 FILLER_69_938 ();
 sg13g2_decap_8 FILLER_69_945 ();
 sg13g2_fill_2 FILLER_69_952 ();
 sg13g2_fill_1 FILLER_69_954 ();
 sg13g2_decap_8 FILLER_69_959 ();
 sg13g2_decap_4 FILLER_69_966 ();
 sg13g2_fill_1 FILLER_69_970 ();
 sg13g2_decap_8 FILLER_69_978 ();
 sg13g2_fill_2 FILLER_69_985 ();
 sg13g2_decap_8 FILLER_69_1018 ();
 sg13g2_decap_4 FILLER_69_1025 ();
 sg13g2_fill_1 FILLER_69_1029 ();
 sg13g2_decap_8 FILLER_69_1035 ();
 sg13g2_decap_8 FILLER_69_1042 ();
 sg13g2_decap_8 FILLER_69_1049 ();
 sg13g2_decap_8 FILLER_69_1056 ();
 sg13g2_decap_4 FILLER_69_1063 ();
 sg13g2_fill_2 FILLER_69_1067 ();
 sg13g2_decap_8 FILLER_69_1076 ();
 sg13g2_fill_2 FILLER_69_1083 ();
 sg13g2_fill_1 FILLER_69_1085 ();
 sg13g2_fill_1 FILLER_69_1134 ();
 sg13g2_fill_2 FILLER_69_1175 ();
 sg13g2_fill_2 FILLER_69_1191 ();
 sg13g2_fill_2 FILLER_69_1225 ();
 sg13g2_fill_2 FILLER_69_1299 ();
 sg13g2_fill_1 FILLER_69_1310 ();
 sg13g2_fill_2 FILLER_69_1330 ();
 sg13g2_fill_2 FILLER_69_1357 ();
 sg13g2_decap_8 FILLER_69_1390 ();
 sg13g2_decap_4 FILLER_69_1397 ();
 sg13g2_fill_2 FILLER_69_1401 ();
 sg13g2_fill_2 FILLER_69_1413 ();
 sg13g2_fill_1 FILLER_69_1443 ();
 sg13g2_fill_2 FILLER_69_1467 ();
 sg13g2_fill_1 FILLER_69_1469 ();
 sg13g2_fill_2 FILLER_69_1491 ();
 sg13g2_fill_2 FILLER_69_1497 ();
 sg13g2_fill_1 FILLER_69_1499 ();
 sg13g2_fill_2 FILLER_69_1510 ();
 sg13g2_decap_8 FILLER_69_1521 ();
 sg13g2_decap_8 FILLER_69_1528 ();
 sg13g2_decap_4 FILLER_69_1535 ();
 sg13g2_decap_8 FILLER_69_1568 ();
 sg13g2_fill_1 FILLER_69_1575 ();
 sg13g2_decap_4 FILLER_69_1580 ();
 sg13g2_fill_2 FILLER_69_1584 ();
 sg13g2_decap_8 FILLER_69_1599 ();
 sg13g2_fill_2 FILLER_69_1606 ();
 sg13g2_fill_2 FILLER_69_1658 ();
 sg13g2_fill_2 FILLER_69_1674 ();
 sg13g2_fill_2 FILLER_69_1737 ();
 sg13g2_fill_1 FILLER_69_1752 ();
 sg13g2_fill_2 FILLER_69_1763 ();
 sg13g2_fill_1 FILLER_69_1765 ();
 sg13g2_fill_2 FILLER_69_1775 ();
 sg13g2_fill_1 FILLER_69_1786 ();
 sg13g2_fill_2 FILLER_69_1818 ();
 sg13g2_fill_2 FILLER_69_1895 ();
 sg13g2_fill_1 FILLER_69_1964 ();
 sg13g2_fill_1 FILLER_69_2128 ();
 sg13g2_decap_4 FILLER_69_2146 ();
 sg13g2_fill_2 FILLER_69_2150 ();
 sg13g2_decap_4 FILLER_69_2179 ();
 sg13g2_fill_1 FILLER_69_2197 ();
 sg13g2_fill_2 FILLER_69_2238 ();
 sg13g2_fill_1 FILLER_69_2240 ();
 sg13g2_decap_8 FILLER_69_2263 ();
 sg13g2_decap_8 FILLER_69_2270 ();
 sg13g2_decap_8 FILLER_69_2277 ();
 sg13g2_fill_2 FILLER_69_2321 ();
 sg13g2_decap_8 FILLER_69_2401 ();
 sg13g2_decap_8 FILLER_69_2408 ();
 sg13g2_decap_8 FILLER_69_2415 ();
 sg13g2_decap_8 FILLER_69_2422 ();
 sg13g2_decap_8 FILLER_69_2429 ();
 sg13g2_decap_8 FILLER_69_2436 ();
 sg13g2_decap_8 FILLER_69_2443 ();
 sg13g2_decap_8 FILLER_69_2450 ();
 sg13g2_decap_8 FILLER_69_2457 ();
 sg13g2_decap_8 FILLER_69_2464 ();
 sg13g2_decap_8 FILLER_69_2471 ();
 sg13g2_decap_8 FILLER_69_2478 ();
 sg13g2_decap_8 FILLER_69_2485 ();
 sg13g2_decap_8 FILLER_69_2492 ();
 sg13g2_decap_8 FILLER_69_2499 ();
 sg13g2_decap_8 FILLER_69_2506 ();
 sg13g2_decap_8 FILLER_69_2513 ();
 sg13g2_decap_8 FILLER_69_2520 ();
 sg13g2_decap_8 FILLER_69_2527 ();
 sg13g2_decap_8 FILLER_69_2534 ();
 sg13g2_decap_8 FILLER_69_2541 ();
 sg13g2_decap_8 FILLER_69_2548 ();
 sg13g2_decap_8 FILLER_69_2555 ();
 sg13g2_decap_8 FILLER_69_2562 ();
 sg13g2_decap_8 FILLER_69_2569 ();
 sg13g2_decap_8 FILLER_69_2576 ();
 sg13g2_decap_8 FILLER_69_2583 ();
 sg13g2_decap_8 FILLER_69_2590 ();
 sg13g2_decap_8 FILLER_69_2597 ();
 sg13g2_decap_8 FILLER_69_2604 ();
 sg13g2_decap_8 FILLER_69_2611 ();
 sg13g2_decap_8 FILLER_69_2618 ();
 sg13g2_decap_8 FILLER_69_2625 ();
 sg13g2_decap_8 FILLER_69_2632 ();
 sg13g2_decap_8 FILLER_69_2639 ();
 sg13g2_decap_8 FILLER_69_2646 ();
 sg13g2_decap_8 FILLER_69_2653 ();
 sg13g2_decap_8 FILLER_69_2660 ();
 sg13g2_decap_8 FILLER_69_2667 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_85 ();
 sg13g2_decap_8 FILLER_70_92 ();
 sg13g2_decap_8 FILLER_70_99 ();
 sg13g2_decap_4 FILLER_70_106 ();
 sg13g2_fill_1 FILLER_70_110 ();
 sg13g2_decap_4 FILLER_70_122 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_224 ();
 sg13g2_decap_4 FILLER_70_234 ();
 sg13g2_fill_2 FILLER_70_238 ();
 sg13g2_fill_2 FILLER_70_249 ();
 sg13g2_fill_2 FILLER_70_291 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_decap_4 FILLER_70_309 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_2 FILLER_70_414 ();
 sg13g2_fill_1 FILLER_70_422 ();
 sg13g2_decap_4 FILLER_70_441 ();
 sg13g2_fill_1 FILLER_70_445 ();
 sg13g2_fill_1 FILLER_70_459 ();
 sg13g2_fill_2 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_519 ();
 sg13g2_fill_2 FILLER_70_526 ();
 sg13g2_fill_2 FILLER_70_589 ();
 sg13g2_fill_1 FILLER_70_591 ();
 sg13g2_fill_2 FILLER_70_598 ();
 sg13g2_fill_2 FILLER_70_628 ();
 sg13g2_fill_1 FILLER_70_630 ();
 sg13g2_fill_1 FILLER_70_660 ();
 sg13g2_fill_1 FILLER_70_683 ();
 sg13g2_fill_2 FILLER_70_761 ();
 sg13g2_fill_1 FILLER_70_763 ();
 sg13g2_fill_2 FILLER_70_768 ();
 sg13g2_fill_1 FILLER_70_786 ();
 sg13g2_fill_1 FILLER_70_882 ();
 sg13g2_fill_1 FILLER_70_896 ();
 sg13g2_decap_4 FILLER_70_936 ();
 sg13g2_fill_2 FILLER_70_940 ();
 sg13g2_fill_2 FILLER_70_945 ();
 sg13g2_fill_1 FILLER_70_947 ();
 sg13g2_decap_8 FILLER_70_966 ();
 sg13g2_decap_4 FILLER_70_973 ();
 sg13g2_fill_1 FILLER_70_983 ();
 sg13g2_fill_2 FILLER_70_997 ();
 sg13g2_fill_1 FILLER_70_999 ();
 sg13g2_decap_8 FILLER_70_1023 ();
 sg13g2_decap_4 FILLER_70_1030 ();
 sg13g2_decap_8 FILLER_70_1045 ();
 sg13g2_decap_8 FILLER_70_1052 ();
 sg13g2_fill_1 FILLER_70_1059 ();
 sg13g2_decap_8 FILLER_70_1065 ();
 sg13g2_decap_8 FILLER_70_1072 ();
 sg13g2_decap_8 FILLER_70_1079 ();
 sg13g2_decap_4 FILLER_70_1086 ();
 sg13g2_fill_1 FILLER_70_1095 ();
 sg13g2_fill_2 FILLER_70_1146 ();
 sg13g2_fill_1 FILLER_70_1148 ();
 sg13g2_fill_1 FILLER_70_1235 ();
 sg13g2_fill_2 FILLER_70_1245 ();
 sg13g2_fill_2 FILLER_70_1257 ();
 sg13g2_fill_1 FILLER_70_1259 ();
 sg13g2_fill_2 FILLER_70_1275 ();
 sg13g2_fill_1 FILLER_70_1277 ();
 sg13g2_fill_2 FILLER_70_1287 ();
 sg13g2_fill_1 FILLER_70_1298 ();
 sg13g2_fill_2 FILLER_70_1320 ();
 sg13g2_fill_1 FILLER_70_1322 ();
 sg13g2_fill_2 FILLER_70_1342 ();
 sg13g2_fill_1 FILLER_70_1344 ();
 sg13g2_fill_1 FILLER_70_1350 ();
 sg13g2_decap_8 FILLER_70_1394 ();
 sg13g2_decap_4 FILLER_70_1401 ();
 sg13g2_fill_2 FILLER_70_1418 ();
 sg13g2_fill_2 FILLER_70_1433 ();
 sg13g2_fill_2 FILLER_70_1478 ();
 sg13g2_fill_2 FILLER_70_1500 ();
 sg13g2_fill_1 FILLER_70_1502 ();
 sg13g2_fill_1 FILLER_70_1538 ();
 sg13g2_fill_1 FILLER_70_1590 ();
 sg13g2_fill_1 FILLER_70_1607 ();
 sg13g2_fill_1 FILLER_70_1659 ();
 sg13g2_fill_2 FILLER_70_1684 ();
 sg13g2_fill_1 FILLER_70_1700 ();
 sg13g2_fill_2 FILLER_70_1767 ();
 sg13g2_fill_1 FILLER_70_1769 ();
 sg13g2_fill_2 FILLER_70_1894 ();
 sg13g2_fill_2 FILLER_70_1935 ();
 sg13g2_fill_1 FILLER_70_1955 ();
 sg13g2_fill_1 FILLER_70_1991 ();
 sg13g2_fill_1 FILLER_70_2001 ();
 sg13g2_fill_2 FILLER_70_2061 ();
 sg13g2_fill_2 FILLER_70_2128 ();
 sg13g2_fill_1 FILLER_70_2165 ();
 sg13g2_fill_2 FILLER_70_2190 ();
 sg13g2_fill_1 FILLER_70_2192 ();
 sg13g2_fill_1 FILLER_70_2213 ();
 sg13g2_fill_1 FILLER_70_2219 ();
 sg13g2_fill_2 FILLER_70_2230 ();
 sg13g2_fill_2 FILLER_70_2265 ();
 sg13g2_fill_1 FILLER_70_2267 ();
 sg13g2_decap_4 FILLER_70_2291 ();
 sg13g2_fill_2 FILLER_70_2340 ();
 sg13g2_fill_1 FILLER_70_2342 ();
 sg13g2_fill_1 FILLER_70_2348 ();
 sg13g2_decap_8 FILLER_70_2390 ();
 sg13g2_decap_8 FILLER_70_2397 ();
 sg13g2_decap_8 FILLER_70_2404 ();
 sg13g2_decap_8 FILLER_70_2411 ();
 sg13g2_decap_8 FILLER_70_2418 ();
 sg13g2_decap_8 FILLER_70_2425 ();
 sg13g2_decap_8 FILLER_70_2432 ();
 sg13g2_decap_8 FILLER_70_2439 ();
 sg13g2_decap_8 FILLER_70_2446 ();
 sg13g2_decap_8 FILLER_70_2453 ();
 sg13g2_decap_8 FILLER_70_2460 ();
 sg13g2_decap_8 FILLER_70_2467 ();
 sg13g2_decap_8 FILLER_70_2474 ();
 sg13g2_decap_8 FILLER_70_2481 ();
 sg13g2_decap_8 FILLER_70_2488 ();
 sg13g2_decap_8 FILLER_70_2495 ();
 sg13g2_decap_8 FILLER_70_2502 ();
 sg13g2_decap_8 FILLER_70_2509 ();
 sg13g2_decap_8 FILLER_70_2516 ();
 sg13g2_decap_8 FILLER_70_2523 ();
 sg13g2_decap_8 FILLER_70_2530 ();
 sg13g2_decap_8 FILLER_70_2537 ();
 sg13g2_decap_8 FILLER_70_2544 ();
 sg13g2_decap_8 FILLER_70_2551 ();
 sg13g2_decap_8 FILLER_70_2558 ();
 sg13g2_decap_8 FILLER_70_2565 ();
 sg13g2_decap_8 FILLER_70_2572 ();
 sg13g2_decap_8 FILLER_70_2579 ();
 sg13g2_decap_8 FILLER_70_2586 ();
 sg13g2_decap_8 FILLER_70_2593 ();
 sg13g2_decap_8 FILLER_70_2600 ();
 sg13g2_decap_8 FILLER_70_2607 ();
 sg13g2_decap_8 FILLER_70_2614 ();
 sg13g2_decap_8 FILLER_70_2621 ();
 sg13g2_decap_8 FILLER_70_2628 ();
 sg13g2_decap_8 FILLER_70_2635 ();
 sg13g2_decap_8 FILLER_70_2642 ();
 sg13g2_decap_8 FILLER_70_2649 ();
 sg13g2_decap_8 FILLER_70_2656 ();
 sg13g2_decap_8 FILLER_70_2663 ();
 sg13g2_decap_4 FILLER_70_2670 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_4 ();
 sg13g2_fill_2 FILLER_71_45 ();
 sg13g2_fill_1 FILLER_71_66 ();
 sg13g2_decap_4 FILLER_71_90 ();
 sg13g2_fill_1 FILLER_71_103 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_129 ();
 sg13g2_fill_2 FILLER_71_139 ();
 sg13g2_fill_1 FILLER_71_141 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_fill_2 FILLER_71_204 ();
 sg13g2_fill_1 FILLER_71_206 ();
 sg13g2_fill_2 FILLER_71_274 ();
 sg13g2_fill_1 FILLER_71_276 ();
 sg13g2_fill_1 FILLER_71_494 ();
 sg13g2_fill_2 FILLER_71_535 ();
 sg13g2_fill_2 FILLER_71_596 ();
 sg13g2_fill_1 FILLER_71_598 ();
 sg13g2_fill_1 FILLER_71_688 ();
 sg13g2_fill_2 FILLER_71_700 ();
 sg13g2_fill_1 FILLER_71_725 ();
 sg13g2_fill_1 FILLER_71_736 ();
 sg13g2_fill_2 FILLER_71_747 ();
 sg13g2_fill_2 FILLER_71_776 ();
 sg13g2_fill_1 FILLER_71_778 ();
 sg13g2_fill_2 FILLER_71_838 ();
 sg13g2_fill_1 FILLER_71_840 ();
 sg13g2_fill_2 FILLER_71_851 ();
 sg13g2_fill_1 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_881 ();
 sg13g2_fill_1 FILLER_71_883 ();
 sg13g2_decap_4 FILLER_71_907 ();
 sg13g2_decap_4 FILLER_71_924 ();
 sg13g2_fill_1 FILLER_71_928 ();
 sg13g2_decap_8 FILLER_71_933 ();
 sg13g2_fill_1 FILLER_71_940 ();
 sg13g2_fill_1 FILLER_71_947 ();
 sg13g2_fill_1 FILLER_71_953 ();
 sg13g2_fill_2 FILLER_71_964 ();
 sg13g2_fill_1 FILLER_71_966 ();
 sg13g2_decap_8 FILLER_71_975 ();
 sg13g2_decap_4 FILLER_71_982 ();
 sg13g2_fill_1 FILLER_71_986 ();
 sg13g2_decap_4 FILLER_71_1015 ();
 sg13g2_fill_2 FILLER_71_1019 ();
 sg13g2_fill_1 FILLER_71_1030 ();
 sg13g2_decap_8 FILLER_71_1044 ();
 sg13g2_fill_2 FILLER_71_1051 ();
 sg13g2_fill_1 FILLER_71_1053 ();
 sg13g2_decap_8 FILLER_71_1073 ();
 sg13g2_decap_8 FILLER_71_1080 ();
 sg13g2_decap_8 FILLER_71_1087 ();
 sg13g2_decap_4 FILLER_71_1094 ();
 sg13g2_fill_2 FILLER_71_1098 ();
 sg13g2_fill_2 FILLER_71_1113 ();
 sg13g2_fill_2 FILLER_71_1133 ();
 sg13g2_fill_1 FILLER_71_1148 ();
 sg13g2_fill_2 FILLER_71_1201 ();
 sg13g2_fill_2 FILLER_71_1282 ();
 sg13g2_fill_2 FILLER_71_1301 ();
 sg13g2_fill_2 FILLER_71_1307 ();
 sg13g2_fill_1 FILLER_71_1309 ();
 sg13g2_fill_2 FILLER_71_1335 ();
 sg13g2_fill_1 FILLER_71_1337 ();
 sg13g2_fill_2 FILLER_71_1381 ();
 sg13g2_fill_1 FILLER_71_1383 ();
 sg13g2_decap_8 FILLER_71_1389 ();
 sg13g2_fill_2 FILLER_71_1396 ();
 sg13g2_fill_1 FILLER_71_1398 ();
 sg13g2_fill_2 FILLER_71_1550 ();
 sg13g2_fill_2 FILLER_71_1592 ();
 sg13g2_fill_2 FILLER_71_1603 ();
 sg13g2_fill_2 FILLER_71_1757 ();
 sg13g2_fill_2 FILLER_71_1772 ();
 sg13g2_fill_1 FILLER_71_1774 ();
 sg13g2_fill_2 FILLER_71_1789 ();
 sg13g2_fill_1 FILLER_71_1791 ();
 sg13g2_fill_2 FILLER_71_1836 ();
 sg13g2_fill_1 FILLER_71_1865 ();
 sg13g2_fill_1 FILLER_71_1932 ();
 sg13g2_fill_2 FILLER_71_1938 ();
 sg13g2_fill_1 FILLER_71_1940 ();
 sg13g2_fill_2 FILLER_71_1954 ();
 sg13g2_fill_1 FILLER_71_1956 ();
 sg13g2_fill_2 FILLER_71_1980 ();
 sg13g2_fill_2 FILLER_71_1987 ();
 sg13g2_fill_2 FILLER_71_2019 ();
 sg13g2_fill_2 FILLER_71_2035 ();
 sg13g2_fill_1 FILLER_71_2037 ();
 sg13g2_fill_2 FILLER_71_2219 ();
 sg13g2_fill_1 FILLER_71_2221 ();
 sg13g2_fill_2 FILLER_71_2240 ();
 sg13g2_fill_2 FILLER_71_2296 ();
 sg13g2_fill_1 FILLER_71_2298 ();
 sg13g2_decap_8 FILLER_71_2382 ();
 sg13g2_decap_8 FILLER_71_2389 ();
 sg13g2_decap_8 FILLER_71_2396 ();
 sg13g2_decap_8 FILLER_71_2403 ();
 sg13g2_decap_8 FILLER_71_2410 ();
 sg13g2_decap_8 FILLER_71_2417 ();
 sg13g2_decap_8 FILLER_71_2424 ();
 sg13g2_decap_8 FILLER_71_2431 ();
 sg13g2_decap_8 FILLER_71_2438 ();
 sg13g2_decap_8 FILLER_71_2445 ();
 sg13g2_decap_8 FILLER_71_2452 ();
 sg13g2_decap_8 FILLER_71_2459 ();
 sg13g2_decap_8 FILLER_71_2466 ();
 sg13g2_decap_8 FILLER_71_2473 ();
 sg13g2_decap_8 FILLER_71_2480 ();
 sg13g2_decap_8 FILLER_71_2487 ();
 sg13g2_decap_8 FILLER_71_2494 ();
 sg13g2_decap_8 FILLER_71_2501 ();
 sg13g2_decap_8 FILLER_71_2508 ();
 sg13g2_decap_8 FILLER_71_2515 ();
 sg13g2_decap_8 FILLER_71_2522 ();
 sg13g2_decap_8 FILLER_71_2529 ();
 sg13g2_decap_8 FILLER_71_2536 ();
 sg13g2_decap_8 FILLER_71_2543 ();
 sg13g2_decap_8 FILLER_71_2550 ();
 sg13g2_decap_8 FILLER_71_2557 ();
 sg13g2_decap_8 FILLER_71_2564 ();
 sg13g2_decap_8 FILLER_71_2571 ();
 sg13g2_decap_8 FILLER_71_2578 ();
 sg13g2_decap_8 FILLER_71_2585 ();
 sg13g2_decap_8 FILLER_71_2592 ();
 sg13g2_decap_8 FILLER_71_2599 ();
 sg13g2_decap_8 FILLER_71_2606 ();
 sg13g2_decap_8 FILLER_71_2613 ();
 sg13g2_decap_8 FILLER_71_2620 ();
 sg13g2_decap_8 FILLER_71_2627 ();
 sg13g2_decap_8 FILLER_71_2634 ();
 sg13g2_decap_8 FILLER_71_2641 ();
 sg13g2_decap_8 FILLER_71_2648 ();
 sg13g2_decap_8 FILLER_71_2655 ();
 sg13g2_decap_8 FILLER_71_2662 ();
 sg13g2_decap_4 FILLER_71_2669 ();
 sg13g2_fill_1 FILLER_71_2673 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_41 ();
 sg13g2_fill_2 FILLER_72_55 ();
 sg13g2_fill_1 FILLER_72_151 ();
 sg13g2_fill_2 FILLER_72_188 ();
 sg13g2_fill_1 FILLER_72_190 ();
 sg13g2_fill_1 FILLER_72_232 ();
 sg13g2_fill_2 FILLER_72_355 ();
 sg13g2_fill_1 FILLER_72_357 ();
 sg13g2_fill_2 FILLER_72_408 ();
 sg13g2_decap_4 FILLER_72_442 ();
 sg13g2_fill_1 FILLER_72_446 ();
 sg13g2_fill_1 FILLER_72_501 ();
 sg13g2_fill_2 FILLER_72_518 ();
 sg13g2_fill_2 FILLER_72_526 ();
 sg13g2_fill_1 FILLER_72_528 ();
 sg13g2_fill_2 FILLER_72_556 ();
 sg13g2_fill_2 FILLER_72_589 ();
 sg13g2_fill_1 FILLER_72_591 ();
 sg13g2_fill_1 FILLER_72_623 ();
 sg13g2_fill_2 FILLER_72_654 ();
 sg13g2_fill_1 FILLER_72_709 ();
 sg13g2_fill_2 FILLER_72_809 ();
 sg13g2_fill_1 FILLER_72_829 ();
 sg13g2_fill_2 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_884 ();
 sg13g2_decap_4 FILLER_72_891 ();
 sg13g2_fill_2 FILLER_72_895 ();
 sg13g2_decap_8 FILLER_72_917 ();
 sg13g2_decap_8 FILLER_72_924 ();
 sg13g2_decap_8 FILLER_72_931 ();
 sg13g2_decap_8 FILLER_72_972 ();
 sg13g2_decap_8 FILLER_72_979 ();
 sg13g2_fill_1 FILLER_72_986 ();
 sg13g2_decap_8 FILLER_72_997 ();
 sg13g2_decap_8 FILLER_72_1004 ();
 sg13g2_fill_2 FILLER_72_1011 ();
 sg13g2_fill_1 FILLER_72_1013 ();
 sg13g2_decap_4 FILLER_72_1019 ();
 sg13g2_fill_2 FILLER_72_1042 ();
 sg13g2_fill_1 FILLER_72_1044 ();
 sg13g2_decap_8 FILLER_72_1050 ();
 sg13g2_decap_8 FILLER_72_1057 ();
 sg13g2_decap_4 FILLER_72_1064 ();
 sg13g2_decap_4 FILLER_72_1073 ();
 sg13g2_decap_4 FILLER_72_1085 ();
 sg13g2_fill_1 FILLER_72_1089 ();
 sg13g2_decap_4 FILLER_72_1220 ();
 sg13g2_fill_1 FILLER_72_1246 ();
 sg13g2_decap_8 FILLER_72_1269 ();
 sg13g2_fill_1 FILLER_72_1276 ();
 sg13g2_fill_2 FILLER_72_1317 ();
 sg13g2_fill_1 FILLER_72_1319 ();
 sg13g2_decap_4 FILLER_72_1346 ();
 sg13g2_fill_1 FILLER_72_1350 ();
 sg13g2_fill_1 FILLER_72_1405 ();
 sg13g2_fill_1 FILLER_72_1444 ();
 sg13g2_fill_1 FILLER_72_1598 ();
 sg13g2_fill_2 FILLER_72_1646 ();
 sg13g2_fill_2 FILLER_72_1666 ();
 sg13g2_fill_2 FILLER_72_1681 ();
 sg13g2_fill_1 FILLER_72_1683 ();
 sg13g2_fill_1 FILLER_72_1691 ();
 sg13g2_fill_1 FILLER_72_1786 ();
 sg13g2_fill_1 FILLER_72_1811 ();
 sg13g2_fill_1 FILLER_72_1857 ();
 sg13g2_fill_2 FILLER_72_1867 ();
 sg13g2_fill_2 FILLER_72_1883 ();
 sg13g2_fill_1 FILLER_72_1916 ();
 sg13g2_fill_2 FILLER_72_1966 ();
 sg13g2_fill_2 FILLER_72_1995 ();
 sg13g2_fill_1 FILLER_72_1997 ();
 sg13g2_fill_1 FILLER_72_2020 ();
 sg13g2_fill_1 FILLER_72_2048 ();
 sg13g2_fill_2 FILLER_72_2071 ();
 sg13g2_fill_2 FILLER_72_2114 ();
 sg13g2_decap_8 FILLER_72_2167 ();
 sg13g2_fill_2 FILLER_72_2174 ();
 sg13g2_fill_1 FILLER_72_2176 ();
 sg13g2_fill_2 FILLER_72_2192 ();
 sg13g2_fill_1 FILLER_72_2227 ();
 sg13g2_fill_1 FILLER_72_2233 ();
 sg13g2_decap_4 FILLER_72_2290 ();
 sg13g2_fill_2 FILLER_72_2294 ();
 sg13g2_fill_2 FILLER_72_2338 ();
 sg13g2_decap_8 FILLER_72_2376 ();
 sg13g2_decap_8 FILLER_72_2383 ();
 sg13g2_decap_8 FILLER_72_2390 ();
 sg13g2_decap_8 FILLER_72_2397 ();
 sg13g2_decap_8 FILLER_72_2404 ();
 sg13g2_decap_8 FILLER_72_2411 ();
 sg13g2_decap_8 FILLER_72_2418 ();
 sg13g2_decap_8 FILLER_72_2425 ();
 sg13g2_decap_8 FILLER_72_2432 ();
 sg13g2_decap_8 FILLER_72_2439 ();
 sg13g2_decap_8 FILLER_72_2446 ();
 sg13g2_decap_8 FILLER_72_2453 ();
 sg13g2_decap_8 FILLER_72_2460 ();
 sg13g2_decap_8 FILLER_72_2467 ();
 sg13g2_decap_8 FILLER_72_2474 ();
 sg13g2_decap_8 FILLER_72_2481 ();
 sg13g2_decap_8 FILLER_72_2488 ();
 sg13g2_decap_8 FILLER_72_2495 ();
 sg13g2_decap_8 FILLER_72_2502 ();
 sg13g2_decap_8 FILLER_72_2509 ();
 sg13g2_decap_8 FILLER_72_2516 ();
 sg13g2_decap_8 FILLER_72_2523 ();
 sg13g2_decap_8 FILLER_72_2530 ();
 sg13g2_decap_8 FILLER_72_2537 ();
 sg13g2_decap_8 FILLER_72_2544 ();
 sg13g2_decap_8 FILLER_72_2551 ();
 sg13g2_decap_8 FILLER_72_2558 ();
 sg13g2_decap_8 FILLER_72_2565 ();
 sg13g2_decap_8 FILLER_72_2572 ();
 sg13g2_decap_8 FILLER_72_2579 ();
 sg13g2_decap_8 FILLER_72_2586 ();
 sg13g2_decap_8 FILLER_72_2593 ();
 sg13g2_decap_8 FILLER_72_2600 ();
 sg13g2_decap_8 FILLER_72_2607 ();
 sg13g2_decap_8 FILLER_72_2614 ();
 sg13g2_decap_8 FILLER_72_2621 ();
 sg13g2_decap_8 FILLER_72_2628 ();
 sg13g2_decap_8 FILLER_72_2635 ();
 sg13g2_decap_8 FILLER_72_2642 ();
 sg13g2_decap_8 FILLER_72_2649 ();
 sg13g2_decap_8 FILLER_72_2656 ();
 sg13g2_decap_8 FILLER_72_2663 ();
 sg13g2_decap_4 FILLER_72_2670 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_1 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_134 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_265 ();
 sg13g2_decap_4 FILLER_73_275 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_fill_2 FILLER_73_323 ();
 sg13g2_fill_2 FILLER_73_396 ();
 sg13g2_decap_4 FILLER_73_439 ();
 sg13g2_fill_1 FILLER_73_443 ();
 sg13g2_fill_1 FILLER_73_457 ();
 sg13g2_fill_1 FILLER_73_480 ();
 sg13g2_fill_2 FILLER_73_518 ();
 sg13g2_fill_1 FILLER_73_520 ();
 sg13g2_fill_1 FILLER_73_529 ();
 sg13g2_decap_8 FILLER_73_624 ();
 sg13g2_fill_1 FILLER_73_653 ();
 sg13g2_fill_1 FILLER_73_687 ();
 sg13g2_fill_2 FILLER_73_756 ();
 sg13g2_fill_1 FILLER_73_758 ();
 sg13g2_fill_2 FILLER_73_810 ();
 sg13g2_fill_1 FILLER_73_812 ();
 sg13g2_fill_1 FILLER_73_832 ();
 sg13g2_fill_2 FILLER_73_846 ();
 sg13g2_decap_8 FILLER_73_865 ();
 sg13g2_fill_2 FILLER_73_872 ();
 sg13g2_fill_1 FILLER_73_874 ();
 sg13g2_decap_8 FILLER_73_889 ();
 sg13g2_decap_4 FILLER_73_896 ();
 sg13g2_decap_8 FILLER_73_905 ();
 sg13g2_decap_8 FILLER_73_912 ();
 sg13g2_decap_8 FILLER_73_919 ();
 sg13g2_decap_8 FILLER_73_926 ();
 sg13g2_decap_8 FILLER_73_933 ();
 sg13g2_decap_4 FILLER_73_940 ();
 sg13g2_fill_2 FILLER_73_944 ();
 sg13g2_fill_1 FILLER_73_966 ();
 sg13g2_fill_1 FILLER_73_977 ();
 sg13g2_decap_8 FILLER_73_984 ();
 sg13g2_decap_8 FILLER_73_991 ();
 sg13g2_fill_2 FILLER_73_998 ();
 sg13g2_decap_8 FILLER_73_1006 ();
 sg13g2_decap_8 FILLER_73_1013 ();
 sg13g2_decap_4 FILLER_73_1020 ();
 sg13g2_fill_1 FILLER_73_1024 ();
 sg13g2_decap_8 FILLER_73_1031 ();
 sg13g2_decap_4 FILLER_73_1038 ();
 sg13g2_fill_2 FILLER_73_1042 ();
 sg13g2_fill_2 FILLER_73_1058 ();
 sg13g2_fill_1 FILLER_73_1060 ();
 sg13g2_fill_1 FILLER_73_1077 ();
 sg13g2_fill_2 FILLER_73_1127 ();
 sg13g2_fill_1 FILLER_73_1129 ();
 sg13g2_fill_2 FILLER_73_1162 ();
 sg13g2_fill_1 FILLER_73_1164 ();
 sg13g2_fill_2 FILLER_73_1218 ();
 sg13g2_decap_4 FILLER_73_1230 ();
 sg13g2_fill_1 FILLER_73_1234 ();
 sg13g2_decap_4 FILLER_73_1262 ();
 sg13g2_fill_2 FILLER_73_1266 ();
 sg13g2_fill_2 FILLER_73_1296 ();
 sg13g2_decap_4 FILLER_73_1352 ();
 sg13g2_fill_1 FILLER_73_1361 ();
 sg13g2_decap_4 FILLER_73_1379 ();
 sg13g2_fill_1 FILLER_73_1383 ();
 sg13g2_fill_1 FILLER_73_1397 ();
 sg13g2_fill_2 FILLER_73_1426 ();
 sg13g2_fill_1 FILLER_73_1428 ();
 sg13g2_fill_2 FILLER_73_1536 ();
 sg13g2_fill_1 FILLER_73_1551 ();
 sg13g2_fill_1 FILLER_73_1591 ();
 sg13g2_fill_1 FILLER_73_1658 ();
 sg13g2_fill_2 FILLER_73_1685 ();
 sg13g2_fill_1 FILLER_73_1715 ();
 sg13g2_fill_2 FILLER_73_1743 ();
 sg13g2_fill_1 FILLER_73_1771 ();
 sg13g2_fill_1 FILLER_73_1847 ();
 sg13g2_fill_1 FILLER_73_1897 ();
 sg13g2_fill_1 FILLER_73_2118 ();
 sg13g2_fill_1 FILLER_73_2159 ();
 sg13g2_fill_1 FILLER_73_2194 ();
 sg13g2_fill_2 FILLER_73_2202 ();
 sg13g2_fill_1 FILLER_73_2204 ();
 sg13g2_fill_2 FILLER_73_2211 ();
 sg13g2_fill_1 FILLER_73_2213 ();
 sg13g2_fill_2 FILLER_73_2228 ();
 sg13g2_fill_1 FILLER_73_2230 ();
 sg13g2_decap_8 FILLER_73_2266 ();
 sg13g2_fill_1 FILLER_73_2273 ();
 sg13g2_fill_2 FILLER_73_2298 ();
 sg13g2_decap_8 FILLER_73_2381 ();
 sg13g2_decap_8 FILLER_73_2388 ();
 sg13g2_decap_8 FILLER_73_2395 ();
 sg13g2_decap_8 FILLER_73_2402 ();
 sg13g2_decap_8 FILLER_73_2409 ();
 sg13g2_decap_8 FILLER_73_2416 ();
 sg13g2_decap_8 FILLER_73_2423 ();
 sg13g2_decap_8 FILLER_73_2430 ();
 sg13g2_decap_8 FILLER_73_2437 ();
 sg13g2_decap_8 FILLER_73_2444 ();
 sg13g2_decap_8 FILLER_73_2451 ();
 sg13g2_decap_8 FILLER_73_2458 ();
 sg13g2_decap_8 FILLER_73_2465 ();
 sg13g2_decap_8 FILLER_73_2472 ();
 sg13g2_decap_8 FILLER_73_2479 ();
 sg13g2_decap_8 FILLER_73_2486 ();
 sg13g2_decap_8 FILLER_73_2493 ();
 sg13g2_decap_8 FILLER_73_2500 ();
 sg13g2_decap_8 FILLER_73_2507 ();
 sg13g2_decap_8 FILLER_73_2514 ();
 sg13g2_decap_8 FILLER_73_2521 ();
 sg13g2_decap_8 FILLER_73_2528 ();
 sg13g2_decap_8 FILLER_73_2535 ();
 sg13g2_decap_8 FILLER_73_2542 ();
 sg13g2_decap_8 FILLER_73_2549 ();
 sg13g2_decap_8 FILLER_73_2556 ();
 sg13g2_decap_8 FILLER_73_2563 ();
 sg13g2_decap_8 FILLER_73_2570 ();
 sg13g2_decap_8 FILLER_73_2577 ();
 sg13g2_decap_8 FILLER_73_2584 ();
 sg13g2_decap_8 FILLER_73_2591 ();
 sg13g2_decap_8 FILLER_73_2598 ();
 sg13g2_decap_8 FILLER_73_2605 ();
 sg13g2_decap_8 FILLER_73_2612 ();
 sg13g2_decap_8 FILLER_73_2619 ();
 sg13g2_decap_8 FILLER_73_2626 ();
 sg13g2_decap_8 FILLER_73_2633 ();
 sg13g2_decap_8 FILLER_73_2640 ();
 sg13g2_decap_8 FILLER_73_2647 ();
 sg13g2_decap_8 FILLER_73_2654 ();
 sg13g2_decap_8 FILLER_73_2661 ();
 sg13g2_decap_4 FILLER_73_2668 ();
 sg13g2_fill_2 FILLER_73_2672 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_131 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_2 FILLER_74_228 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_decap_4 FILLER_74_310 ();
 sg13g2_fill_2 FILLER_74_373 ();
 sg13g2_fill_2 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_403 ();
 sg13g2_decap_8 FILLER_74_432 ();
 sg13g2_fill_2 FILLER_74_460 ();
 sg13g2_fill_1 FILLER_74_471 ();
 sg13g2_fill_1 FILLER_74_522 ();
 sg13g2_fill_1 FILLER_74_577 ();
 sg13g2_decap_8 FILLER_74_614 ();
 sg13g2_fill_2 FILLER_74_621 ();
 sg13g2_fill_1 FILLER_74_623 ();
 sg13g2_fill_1 FILLER_74_640 ();
 sg13g2_fill_2 FILLER_74_656 ();
 sg13g2_fill_2 FILLER_74_714 ();
 sg13g2_fill_1 FILLER_74_722 ();
 sg13g2_fill_2 FILLER_74_729 ();
 sg13g2_fill_1 FILLER_74_754 ();
 sg13g2_fill_1 FILLER_74_835 ();
 sg13g2_fill_2 FILLER_74_863 ();
 sg13g2_fill_1 FILLER_74_865 ();
 sg13g2_decap_8 FILLER_74_871 ();
 sg13g2_decap_4 FILLER_74_878 ();
 sg13g2_decap_8 FILLER_74_901 ();
 sg13g2_decap_8 FILLER_74_908 ();
 sg13g2_fill_2 FILLER_74_915 ();
 sg13g2_fill_1 FILLER_74_917 ();
 sg13g2_fill_1 FILLER_74_926 ();
 sg13g2_decap_8 FILLER_74_936 ();
 sg13g2_decap_8 FILLER_74_943 ();
 sg13g2_decap_8 FILLER_74_950 ();
 sg13g2_decap_8 FILLER_74_957 ();
 sg13g2_decap_8 FILLER_74_964 ();
 sg13g2_decap_4 FILLER_74_971 ();
 sg13g2_fill_2 FILLER_74_975 ();
 sg13g2_decap_8 FILLER_74_987 ();
 sg13g2_decap_8 FILLER_74_994 ();
 sg13g2_decap_8 FILLER_74_1001 ();
 sg13g2_fill_2 FILLER_74_1008 ();
 sg13g2_fill_1 FILLER_74_1014 ();
 sg13g2_decap_8 FILLER_74_1021 ();
 sg13g2_decap_8 FILLER_74_1028 ();
 sg13g2_decap_8 FILLER_74_1035 ();
 sg13g2_decap_8 FILLER_74_1042 ();
 sg13g2_decap_8 FILLER_74_1049 ();
 sg13g2_fill_2 FILLER_74_1056 ();
 sg13g2_fill_1 FILLER_74_1058 ();
 sg13g2_fill_2 FILLER_74_1090 ();
 sg13g2_fill_1 FILLER_74_1113 ();
 sg13g2_fill_1 FILLER_74_1185 ();
 sg13g2_fill_2 FILLER_74_1226 ();
 sg13g2_fill_1 FILLER_74_1228 ();
 sg13g2_fill_1 FILLER_74_1266 ();
 sg13g2_fill_1 FILLER_74_1326 ();
 sg13g2_decap_8 FILLER_74_1342 ();
 sg13g2_decap_4 FILLER_74_1363 ();
 sg13g2_decap_8 FILLER_74_1380 ();
 sg13g2_fill_2 FILLER_74_1387 ();
 sg13g2_fill_1 FILLER_74_1389 ();
 sg13g2_fill_1 FILLER_74_1407 ();
 sg13g2_fill_1 FILLER_74_1413 ();
 sg13g2_fill_1 FILLER_74_1499 ();
 sg13g2_fill_1 FILLER_74_1512 ();
 sg13g2_fill_1 FILLER_74_1540 ();
 sg13g2_fill_2 FILLER_74_1554 ();
 sg13g2_fill_1 FILLER_74_1640 ();
 sg13g2_fill_2 FILLER_74_1704 ();
 sg13g2_fill_1 FILLER_74_1706 ();
 sg13g2_fill_2 FILLER_74_1734 ();
 sg13g2_fill_2 FILLER_74_1847 ();
 sg13g2_fill_1 FILLER_74_1886 ();
 sg13g2_fill_2 FILLER_74_1910 ();
 sg13g2_fill_2 FILLER_74_1980 ();
 sg13g2_fill_2 FILLER_74_2009 ();
 sg13g2_fill_1 FILLER_74_2011 ();
 sg13g2_fill_1 FILLER_74_2033 ();
 sg13g2_fill_1 FILLER_74_2053 ();
 sg13g2_fill_2 FILLER_74_2060 ();
 sg13g2_fill_1 FILLER_74_2202 ();
 sg13g2_fill_1 FILLER_74_2227 ();
 sg13g2_fill_2 FILLER_74_2233 ();
 sg13g2_fill_1 FILLER_74_2235 ();
 sg13g2_fill_2 FILLER_74_2271 ();
 sg13g2_decap_8 FILLER_74_2373 ();
 sg13g2_decap_8 FILLER_74_2380 ();
 sg13g2_decap_8 FILLER_74_2387 ();
 sg13g2_decap_8 FILLER_74_2394 ();
 sg13g2_decap_8 FILLER_74_2401 ();
 sg13g2_decap_8 FILLER_74_2408 ();
 sg13g2_decap_8 FILLER_74_2415 ();
 sg13g2_decap_8 FILLER_74_2422 ();
 sg13g2_decap_8 FILLER_74_2429 ();
 sg13g2_decap_8 FILLER_74_2436 ();
 sg13g2_decap_8 FILLER_74_2443 ();
 sg13g2_decap_8 FILLER_74_2450 ();
 sg13g2_decap_8 FILLER_74_2457 ();
 sg13g2_decap_8 FILLER_74_2464 ();
 sg13g2_decap_8 FILLER_74_2471 ();
 sg13g2_decap_8 FILLER_74_2478 ();
 sg13g2_decap_8 FILLER_74_2485 ();
 sg13g2_decap_8 FILLER_74_2492 ();
 sg13g2_decap_8 FILLER_74_2499 ();
 sg13g2_decap_8 FILLER_74_2506 ();
 sg13g2_decap_8 FILLER_74_2513 ();
 sg13g2_decap_8 FILLER_74_2520 ();
 sg13g2_decap_8 FILLER_74_2527 ();
 sg13g2_decap_8 FILLER_74_2534 ();
 sg13g2_decap_8 FILLER_74_2541 ();
 sg13g2_decap_8 FILLER_74_2548 ();
 sg13g2_decap_8 FILLER_74_2555 ();
 sg13g2_decap_8 FILLER_74_2562 ();
 sg13g2_decap_8 FILLER_74_2569 ();
 sg13g2_decap_8 FILLER_74_2576 ();
 sg13g2_decap_8 FILLER_74_2583 ();
 sg13g2_decap_8 FILLER_74_2590 ();
 sg13g2_decap_8 FILLER_74_2597 ();
 sg13g2_decap_8 FILLER_74_2604 ();
 sg13g2_decap_8 FILLER_74_2611 ();
 sg13g2_decap_8 FILLER_74_2618 ();
 sg13g2_decap_8 FILLER_74_2625 ();
 sg13g2_decap_8 FILLER_74_2632 ();
 sg13g2_decap_8 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2646 ();
 sg13g2_decap_8 FILLER_74_2653 ();
 sg13g2_decap_8 FILLER_74_2660 ();
 sg13g2_decap_8 FILLER_74_2667 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_41 ();
 sg13g2_fill_1 FILLER_75_43 ();
 sg13g2_fill_2 FILLER_75_67 ();
 sg13g2_fill_2 FILLER_75_125 ();
 sg13g2_fill_2 FILLER_75_136 ();
 sg13g2_fill_2 FILLER_75_174 ();
 sg13g2_fill_2 FILLER_75_198 ();
 sg13g2_fill_2 FILLER_75_247 ();
 sg13g2_fill_2 FILLER_75_303 ();
 sg13g2_fill_2 FILLER_75_313 ();
 sg13g2_fill_1 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_366 ();
 sg13g2_fill_1 FILLER_75_368 ();
 sg13g2_fill_1 FILLER_75_426 ();
 sg13g2_decap_4 FILLER_75_433 ();
 sg13g2_fill_1 FILLER_75_451 ();
 sg13g2_fill_2 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_500 ();
 sg13g2_fill_2 FILLER_75_525 ();
 sg13g2_fill_2 FILLER_75_558 ();
 sg13g2_fill_1 FILLER_75_560 ();
 sg13g2_fill_2 FILLER_75_568 ();
 sg13g2_fill_2 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_619 ();
 sg13g2_fill_1 FILLER_75_844 ();
 sg13g2_fill_1 FILLER_75_917 ();
 sg13g2_decap_8 FILLER_75_943 ();
 sg13g2_decap_8 FILLER_75_950 ();
 sg13g2_fill_1 FILLER_75_957 ();
 sg13g2_decap_4 FILLER_75_962 ();
 sg13g2_decap_8 FILLER_75_970 ();
 sg13g2_decap_8 FILLER_75_977 ();
 sg13g2_decap_8 FILLER_75_984 ();
 sg13g2_decap_8 FILLER_75_991 ();
 sg13g2_fill_2 FILLER_75_998 ();
 sg13g2_fill_1 FILLER_75_1000 ();
 sg13g2_decap_8 FILLER_75_1024 ();
 sg13g2_decap_4 FILLER_75_1031 ();
 sg13g2_fill_2 FILLER_75_1035 ();
 sg13g2_decap_8 FILLER_75_1042 ();
 sg13g2_fill_2 FILLER_75_1049 ();
 sg13g2_fill_1 FILLER_75_1074 ();
 sg13g2_fill_1 FILLER_75_1125 ();
 sg13g2_decap_4 FILLER_75_1234 ();
 sg13g2_fill_2 FILLER_75_1315 ();
 sg13g2_fill_1 FILLER_75_1324 ();
 sg13g2_fill_2 FILLER_75_1340 ();
 sg13g2_fill_1 FILLER_75_1342 ();
 sg13g2_decap_4 FILLER_75_1352 ();
 sg13g2_fill_1 FILLER_75_1356 ();
 sg13g2_fill_2 FILLER_75_1385 ();
 sg13g2_fill_1 FILLER_75_1433 ();
 sg13g2_fill_1 FILLER_75_1481 ();
 sg13g2_fill_2 FILLER_75_1495 ();
 sg13g2_fill_1 FILLER_75_1537 ();
 sg13g2_fill_2 FILLER_75_1584 ();
 sg13g2_fill_1 FILLER_75_1595 ();
 sg13g2_fill_1 FILLER_75_1605 ();
 sg13g2_fill_1 FILLER_75_1620 ();
 sg13g2_fill_2 FILLER_75_1634 ();
 sg13g2_fill_1 FILLER_75_1684 ();
 sg13g2_fill_2 FILLER_75_1730 ();
 sg13g2_fill_2 FILLER_75_1768 ();
 sg13g2_fill_1 FILLER_75_1770 ();
 sg13g2_fill_1 FILLER_75_1785 ();
 sg13g2_fill_2 FILLER_75_1822 ();
 sg13g2_fill_1 FILLER_75_1824 ();
 sg13g2_fill_1 FILLER_75_1838 ();
 sg13g2_fill_1 FILLER_75_1935 ();
 sg13g2_fill_1 FILLER_75_1974 ();
 sg13g2_fill_2 FILLER_75_1984 ();
 sg13g2_fill_1 FILLER_75_1986 ();
 sg13g2_fill_2 FILLER_75_2021 ();
 sg13g2_fill_1 FILLER_75_2023 ();
 sg13g2_fill_1 FILLER_75_2073 ();
 sg13g2_fill_1 FILLER_75_2104 ();
 sg13g2_fill_1 FILLER_75_2138 ();
 sg13g2_decap_8 FILLER_75_2148 ();
 sg13g2_decap_4 FILLER_75_2155 ();
 sg13g2_fill_1 FILLER_75_2159 ();
 sg13g2_fill_1 FILLER_75_2174 ();
 sg13g2_fill_1 FILLER_75_2203 ();
 sg13g2_fill_1 FILLER_75_2227 ();
 sg13g2_fill_1 FILLER_75_2245 ();
 sg13g2_fill_2 FILLER_75_2313 ();
 sg13g2_fill_1 FILLER_75_2315 ();
 sg13g2_fill_1 FILLER_75_2352 ();
 sg13g2_decap_8 FILLER_75_2375 ();
 sg13g2_decap_8 FILLER_75_2382 ();
 sg13g2_decap_8 FILLER_75_2389 ();
 sg13g2_decap_8 FILLER_75_2396 ();
 sg13g2_decap_8 FILLER_75_2403 ();
 sg13g2_decap_8 FILLER_75_2410 ();
 sg13g2_decap_8 FILLER_75_2417 ();
 sg13g2_decap_8 FILLER_75_2424 ();
 sg13g2_decap_8 FILLER_75_2431 ();
 sg13g2_decap_8 FILLER_75_2438 ();
 sg13g2_decap_8 FILLER_75_2445 ();
 sg13g2_decap_8 FILLER_75_2452 ();
 sg13g2_decap_8 FILLER_75_2459 ();
 sg13g2_decap_8 FILLER_75_2466 ();
 sg13g2_decap_8 FILLER_75_2473 ();
 sg13g2_decap_8 FILLER_75_2480 ();
 sg13g2_decap_8 FILLER_75_2487 ();
 sg13g2_decap_8 FILLER_75_2494 ();
 sg13g2_decap_8 FILLER_75_2501 ();
 sg13g2_decap_8 FILLER_75_2508 ();
 sg13g2_decap_8 FILLER_75_2515 ();
 sg13g2_decap_8 FILLER_75_2522 ();
 sg13g2_decap_8 FILLER_75_2529 ();
 sg13g2_decap_8 FILLER_75_2536 ();
 sg13g2_decap_8 FILLER_75_2543 ();
 sg13g2_decap_8 FILLER_75_2550 ();
 sg13g2_decap_8 FILLER_75_2557 ();
 sg13g2_decap_8 FILLER_75_2564 ();
 sg13g2_decap_8 FILLER_75_2571 ();
 sg13g2_decap_8 FILLER_75_2578 ();
 sg13g2_decap_8 FILLER_75_2585 ();
 sg13g2_decap_8 FILLER_75_2592 ();
 sg13g2_decap_8 FILLER_75_2599 ();
 sg13g2_decap_8 FILLER_75_2606 ();
 sg13g2_decap_8 FILLER_75_2613 ();
 sg13g2_decap_8 FILLER_75_2620 ();
 sg13g2_decap_8 FILLER_75_2627 ();
 sg13g2_decap_8 FILLER_75_2634 ();
 sg13g2_decap_8 FILLER_75_2641 ();
 sg13g2_decap_8 FILLER_75_2648 ();
 sg13g2_decap_8 FILLER_75_2655 ();
 sg13g2_decap_8 FILLER_75_2662 ();
 sg13g2_decap_4 FILLER_75_2669 ();
 sg13g2_fill_1 FILLER_75_2673 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_69 ();
 sg13g2_fill_1 FILLER_76_83 ();
 sg13g2_fill_1 FILLER_76_144 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_fill_1 FILLER_76_200 ();
 sg13g2_fill_1 FILLER_76_205 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_4 FILLER_76_273 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_fill_1 FILLER_76_320 ();
 sg13g2_fill_2 FILLER_76_398 ();
 sg13g2_fill_1 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_432 ();
 sg13g2_fill_1 FILLER_76_495 ();
 sg13g2_fill_2 FILLER_76_506 ();
 sg13g2_fill_1 FILLER_76_508 ();
 sg13g2_fill_1 FILLER_76_519 ();
 sg13g2_fill_2 FILLER_76_588 ();
 sg13g2_fill_1 FILLER_76_621 ();
 sg13g2_fill_2 FILLER_76_790 ();
 sg13g2_fill_1 FILLER_76_871 ();
 sg13g2_fill_2 FILLER_76_885 ();
 sg13g2_decap_4 FILLER_76_900 ();
 sg13g2_fill_2 FILLER_76_917 ();
 sg13g2_fill_1 FILLER_76_942 ();
 sg13g2_decap_8 FILLER_76_947 ();
 sg13g2_decap_4 FILLER_76_954 ();
 sg13g2_decap_8 FILLER_76_982 ();
 sg13g2_fill_2 FILLER_76_989 ();
 sg13g2_decap_4 FILLER_76_1039 ();
 sg13g2_fill_2 FILLER_76_1043 ();
 sg13g2_decap_4 FILLER_76_1053 ();
 sg13g2_fill_1 FILLER_76_1057 ();
 sg13g2_decap_8 FILLER_76_1069 ();
 sg13g2_fill_2 FILLER_76_1076 ();
 sg13g2_fill_1 FILLER_76_1100 ();
 sg13g2_fill_2 FILLER_76_1115 ();
 sg13g2_fill_2 FILLER_76_1218 ();
 sg13g2_fill_1 FILLER_76_1220 ();
 sg13g2_decap_4 FILLER_76_1239 ();
 sg13g2_fill_2 FILLER_76_1252 ();
 sg13g2_decap_8 FILLER_76_1267 ();
 sg13g2_fill_1 FILLER_76_1274 ();
 sg13g2_fill_1 FILLER_76_1288 ();
 sg13g2_fill_2 FILLER_76_1341 ();
 sg13g2_fill_1 FILLER_76_1343 ();
 sg13g2_fill_2 FILLER_76_1372 ();
 sg13g2_fill_1 FILLER_76_1374 ();
 sg13g2_fill_2 FILLER_76_1428 ();
 sg13g2_fill_1 FILLER_76_1430 ();
 sg13g2_fill_2 FILLER_76_1488 ();
 sg13g2_fill_2 FILLER_76_1540 ();
 sg13g2_fill_2 FILLER_76_1582 ();
 sg13g2_fill_1 FILLER_76_1611 ();
 sg13g2_fill_2 FILLER_76_1708 ();
 sg13g2_fill_2 FILLER_76_1766 ();
 sg13g2_fill_2 FILLER_76_1777 ();
 sg13g2_fill_1 FILLER_76_1801 ();
 sg13g2_fill_2 FILLER_76_1846 ();
 sg13g2_fill_1 FILLER_76_1887 ();
 sg13g2_fill_2 FILLER_76_1942 ();
 sg13g2_decap_8 FILLER_76_2023 ();
 sg13g2_decap_8 FILLER_76_2137 ();
 sg13g2_decap_8 FILLER_76_2144 ();
 sg13g2_decap_8 FILLER_76_2151 ();
 sg13g2_decap_8 FILLER_76_2158 ();
 sg13g2_decap_8 FILLER_76_2165 ();
 sg13g2_fill_2 FILLER_76_2172 ();
 sg13g2_fill_2 FILLER_76_2235 ();
 sg13g2_fill_1 FILLER_76_2237 ();
 sg13g2_decap_4 FILLER_76_2289 ();
 sg13g2_fill_2 FILLER_76_2302 ();
 sg13g2_fill_1 FILLER_76_2340 ();
 sg13g2_decap_8 FILLER_76_2364 ();
 sg13g2_decap_8 FILLER_76_2371 ();
 sg13g2_decap_8 FILLER_76_2378 ();
 sg13g2_decap_8 FILLER_76_2385 ();
 sg13g2_decap_8 FILLER_76_2392 ();
 sg13g2_decap_8 FILLER_76_2399 ();
 sg13g2_decap_8 FILLER_76_2406 ();
 sg13g2_decap_8 FILLER_76_2413 ();
 sg13g2_decap_8 FILLER_76_2420 ();
 sg13g2_decap_8 FILLER_76_2427 ();
 sg13g2_decap_8 FILLER_76_2434 ();
 sg13g2_decap_8 FILLER_76_2441 ();
 sg13g2_decap_8 FILLER_76_2448 ();
 sg13g2_decap_8 FILLER_76_2455 ();
 sg13g2_decap_8 FILLER_76_2462 ();
 sg13g2_decap_8 FILLER_76_2469 ();
 sg13g2_decap_8 FILLER_76_2476 ();
 sg13g2_decap_8 FILLER_76_2483 ();
 sg13g2_decap_8 FILLER_76_2490 ();
 sg13g2_decap_8 FILLER_76_2497 ();
 sg13g2_decap_8 FILLER_76_2504 ();
 sg13g2_decap_8 FILLER_76_2511 ();
 sg13g2_decap_8 FILLER_76_2518 ();
 sg13g2_decap_8 FILLER_76_2525 ();
 sg13g2_decap_8 FILLER_76_2532 ();
 sg13g2_decap_8 FILLER_76_2539 ();
 sg13g2_decap_8 FILLER_76_2546 ();
 sg13g2_decap_8 FILLER_76_2553 ();
 sg13g2_decap_8 FILLER_76_2560 ();
 sg13g2_decap_8 FILLER_76_2567 ();
 sg13g2_decap_8 FILLER_76_2574 ();
 sg13g2_decap_8 FILLER_76_2581 ();
 sg13g2_decap_8 FILLER_76_2588 ();
 sg13g2_decap_8 FILLER_76_2595 ();
 sg13g2_decap_8 FILLER_76_2602 ();
 sg13g2_decap_8 FILLER_76_2609 ();
 sg13g2_decap_8 FILLER_76_2616 ();
 sg13g2_decap_8 FILLER_76_2623 ();
 sg13g2_decap_8 FILLER_76_2630 ();
 sg13g2_decap_8 FILLER_76_2637 ();
 sg13g2_decap_8 FILLER_76_2644 ();
 sg13g2_decap_8 FILLER_76_2651 ();
 sg13g2_decap_8 FILLER_76_2658 ();
 sg13g2_decap_8 FILLER_76_2665 ();
 sg13g2_fill_2 FILLER_76_2672 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_fill_1 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_56 ();
 sg13g2_fill_1 FILLER_77_106 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_257 ();
 sg13g2_decap_4 FILLER_77_264 ();
 sg13g2_fill_2 FILLER_77_268 ();
 sg13g2_fill_2 FILLER_77_302 ();
 sg13g2_fill_1 FILLER_77_304 ();
 sg13g2_fill_2 FILLER_77_349 ();
 sg13g2_fill_1 FILLER_77_351 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_fill_2 FILLER_77_460 ();
 sg13g2_fill_2 FILLER_77_480 ();
 sg13g2_fill_1 FILLER_77_482 ();
 sg13g2_fill_2 FILLER_77_493 ();
 sg13g2_fill_1 FILLER_77_495 ();
 sg13g2_fill_1 FILLER_77_505 ();
 sg13g2_decap_4 FILLER_77_557 ();
 sg13g2_fill_1 FILLER_77_576 ();
 sg13g2_fill_2 FILLER_77_583 ();
 sg13g2_fill_1 FILLER_77_591 ();
 sg13g2_fill_2 FILLER_77_625 ();
 sg13g2_fill_1 FILLER_77_627 ();
 sg13g2_fill_1 FILLER_77_665 ();
 sg13g2_fill_1 FILLER_77_703 ();
 sg13g2_fill_1 FILLER_77_824 ();
 sg13g2_fill_2 FILLER_77_838 ();
 sg13g2_fill_1 FILLER_77_840 ();
 sg13g2_fill_2 FILLER_77_851 ();
 sg13g2_fill_1 FILLER_77_901 ();
 sg13g2_fill_1 FILLER_77_945 ();
 sg13g2_decap_4 FILLER_77_951 ();
 sg13g2_fill_1 FILLER_77_955 ();
 sg13g2_decap_8 FILLER_77_964 ();
 sg13g2_fill_2 FILLER_77_1003 ();
 sg13g2_fill_1 FILLER_77_1005 ();
 sg13g2_decap_8 FILLER_77_1042 ();
 sg13g2_fill_2 FILLER_77_1049 ();
 sg13g2_fill_2 FILLER_77_1074 ();
 sg13g2_fill_2 FILLER_77_1126 ();
 sg13g2_fill_2 FILLER_77_1196 ();
 sg13g2_fill_1 FILLER_77_1198 ();
 sg13g2_decap_4 FILLER_77_1219 ();
 sg13g2_fill_2 FILLER_77_1223 ();
 sg13g2_fill_1 FILLER_77_1253 ();
 sg13g2_decap_4 FILLER_77_1267 ();
 sg13g2_fill_2 FILLER_77_1299 ();
 sg13g2_decap_4 FILLER_77_1338 ();
 sg13g2_fill_1 FILLER_77_1355 ();
 sg13g2_fill_2 FILLER_77_1396 ();
 sg13g2_fill_1 FILLER_77_1398 ();
 sg13g2_fill_1 FILLER_77_1566 ();
 sg13g2_fill_2 FILLER_77_1734 ();
 sg13g2_fill_1 FILLER_77_1736 ();
 sg13g2_fill_1 FILLER_77_1751 ();
 sg13g2_fill_1 FILLER_77_1779 ();
 sg13g2_fill_1 FILLER_77_1916 ();
 sg13g2_fill_2 FILLER_77_1981 ();
 sg13g2_fill_2 FILLER_77_2037 ();
 sg13g2_fill_1 FILLER_77_2066 ();
 sg13g2_decap_8 FILLER_77_2132 ();
 sg13g2_decap_8 FILLER_77_2139 ();
 sg13g2_decap_8 FILLER_77_2146 ();
 sg13g2_decap_8 FILLER_77_2153 ();
 sg13g2_decap_8 FILLER_77_2160 ();
 sg13g2_decap_8 FILLER_77_2167 ();
 sg13g2_fill_1 FILLER_77_2174 ();
 sg13g2_fill_1 FILLER_77_2233 ();
 sg13g2_fill_2 FILLER_77_2285 ();
 sg13g2_decap_4 FILLER_77_2305 ();
 sg13g2_decap_8 FILLER_77_2313 ();
 sg13g2_fill_1 FILLER_77_2320 ();
 sg13g2_decap_8 FILLER_77_2353 ();
 sg13g2_decap_8 FILLER_77_2360 ();
 sg13g2_decap_8 FILLER_77_2367 ();
 sg13g2_decap_8 FILLER_77_2374 ();
 sg13g2_decap_8 FILLER_77_2381 ();
 sg13g2_decap_8 FILLER_77_2388 ();
 sg13g2_decap_8 FILLER_77_2395 ();
 sg13g2_decap_8 FILLER_77_2402 ();
 sg13g2_decap_8 FILLER_77_2409 ();
 sg13g2_decap_8 FILLER_77_2416 ();
 sg13g2_decap_8 FILLER_77_2423 ();
 sg13g2_decap_8 FILLER_77_2430 ();
 sg13g2_decap_8 FILLER_77_2437 ();
 sg13g2_decap_8 FILLER_77_2444 ();
 sg13g2_decap_8 FILLER_77_2451 ();
 sg13g2_decap_8 FILLER_77_2458 ();
 sg13g2_decap_8 FILLER_77_2465 ();
 sg13g2_decap_8 FILLER_77_2472 ();
 sg13g2_decap_8 FILLER_77_2479 ();
 sg13g2_decap_8 FILLER_77_2486 ();
 sg13g2_decap_8 FILLER_77_2493 ();
 sg13g2_decap_8 FILLER_77_2500 ();
 sg13g2_decap_8 FILLER_77_2507 ();
 sg13g2_decap_8 FILLER_77_2514 ();
 sg13g2_decap_8 FILLER_77_2521 ();
 sg13g2_decap_8 FILLER_77_2528 ();
 sg13g2_decap_8 FILLER_77_2535 ();
 sg13g2_decap_8 FILLER_77_2542 ();
 sg13g2_decap_8 FILLER_77_2549 ();
 sg13g2_decap_8 FILLER_77_2556 ();
 sg13g2_decap_8 FILLER_77_2563 ();
 sg13g2_decap_8 FILLER_77_2570 ();
 sg13g2_decap_8 FILLER_77_2577 ();
 sg13g2_decap_8 FILLER_77_2584 ();
 sg13g2_decap_8 FILLER_77_2591 ();
 sg13g2_decap_8 FILLER_77_2598 ();
 sg13g2_decap_8 FILLER_77_2605 ();
 sg13g2_decap_8 FILLER_77_2612 ();
 sg13g2_decap_8 FILLER_77_2619 ();
 sg13g2_decap_8 FILLER_77_2626 ();
 sg13g2_decap_8 FILLER_77_2633 ();
 sg13g2_decap_8 FILLER_77_2640 ();
 sg13g2_decap_8 FILLER_77_2647 ();
 sg13g2_decap_8 FILLER_77_2654 ();
 sg13g2_decap_8 FILLER_77_2661 ();
 sg13g2_decap_4 FILLER_77_2668 ();
 sg13g2_fill_2 FILLER_77_2672 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_fill_1 FILLER_78_104 ();
 sg13g2_fill_1 FILLER_78_165 ();
 sg13g2_decap_4 FILLER_78_194 ();
 sg13g2_fill_1 FILLER_78_198 ();
 sg13g2_fill_1 FILLER_78_259 ();
 sg13g2_fill_2 FILLER_78_300 ();
 sg13g2_fill_2 FILLER_78_311 ();
 sg13g2_fill_1 FILLER_78_313 ();
 sg13g2_fill_1 FILLER_78_368 ();
 sg13g2_fill_1 FILLER_78_397 ();
 sg13g2_fill_2 FILLER_78_403 ();
 sg13g2_fill_1 FILLER_78_445 ();
 sg13g2_fill_2 FILLER_78_507 ();
 sg13g2_fill_2 FILLER_78_522 ();
 sg13g2_decap_8 FILLER_78_556 ();
 sg13g2_decap_4 FILLER_78_563 ();
 sg13g2_fill_1 FILLER_78_580 ();
 sg13g2_fill_2 FILLER_78_596 ();
 sg13g2_fill_2 FILLER_78_715 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_fill_1 FILLER_78_791 ();
 sg13g2_fill_2 FILLER_78_842 ();
 sg13g2_fill_1 FILLER_78_844 ();
 sg13g2_fill_2 FILLER_78_921 ();
 sg13g2_fill_2 FILLER_78_933 ();
 sg13g2_fill_1 FILLER_78_953 ();
 sg13g2_decap_8 FILLER_78_963 ();
 sg13g2_fill_1 FILLER_78_970 ();
 sg13g2_fill_2 FILLER_78_977 ();
 sg13g2_decap_4 FILLER_78_1006 ();
 sg13g2_fill_2 FILLER_78_1043 ();
 sg13g2_fill_1 FILLER_78_1049 ();
 sg13g2_fill_2 FILLER_78_1080 ();
 sg13g2_fill_1 FILLER_78_1082 ();
 sg13g2_fill_2 FILLER_78_1147 ();
 sg13g2_fill_1 FILLER_78_1149 ();
 sg13g2_decap_8 FILLER_78_1250 ();
 sg13g2_fill_2 FILLER_78_1285 ();
 sg13g2_fill_1 FILLER_78_1287 ();
 sg13g2_fill_1 FILLER_78_1316 ();
 sg13g2_fill_2 FILLER_78_1349 ();
 sg13g2_fill_1 FILLER_78_1351 ();
 sg13g2_fill_2 FILLER_78_1392 ();
 sg13g2_fill_2 FILLER_78_1444 ();
 sg13g2_fill_2 FILLER_78_1451 ();
 sg13g2_fill_1 FILLER_78_1453 ();
 sg13g2_fill_1 FILLER_78_1490 ();
 sg13g2_fill_2 FILLER_78_1524 ();
 sg13g2_fill_1 FILLER_78_1665 ();
 sg13g2_fill_2 FILLER_78_1746 ();
 sg13g2_fill_2 FILLER_78_1802 ();
 sg13g2_fill_1 FILLER_78_1814 ();
 sg13g2_fill_2 FILLER_78_1847 ();
 sg13g2_fill_1 FILLER_78_1988 ();
 sg13g2_fill_2 FILLER_78_2035 ();
 sg13g2_fill_1 FILLER_78_2037 ();
 sg13g2_fill_2 FILLER_78_2066 ();
 sg13g2_fill_1 FILLER_78_2068 ();
 sg13g2_fill_1 FILLER_78_2101 ();
 sg13g2_decap_8 FILLER_78_2121 ();
 sg13g2_decap_8 FILLER_78_2128 ();
 sg13g2_decap_8 FILLER_78_2135 ();
 sg13g2_decap_8 FILLER_78_2142 ();
 sg13g2_decap_8 FILLER_78_2149 ();
 sg13g2_decap_8 FILLER_78_2156 ();
 sg13g2_decap_8 FILLER_78_2163 ();
 sg13g2_decap_8 FILLER_78_2170 ();
 sg13g2_decap_8 FILLER_78_2177 ();
 sg13g2_decap_4 FILLER_78_2184 ();
 sg13g2_fill_1 FILLER_78_2247 ();
 sg13g2_decap_8 FILLER_78_2303 ();
 sg13g2_decap_8 FILLER_78_2310 ();
 sg13g2_decap_8 FILLER_78_2317 ();
 sg13g2_decap_8 FILLER_78_2324 ();
 sg13g2_decap_8 FILLER_78_2331 ();
 sg13g2_decap_8 FILLER_78_2338 ();
 sg13g2_decap_8 FILLER_78_2345 ();
 sg13g2_decap_8 FILLER_78_2352 ();
 sg13g2_decap_8 FILLER_78_2359 ();
 sg13g2_decap_8 FILLER_78_2366 ();
 sg13g2_decap_8 FILLER_78_2373 ();
 sg13g2_decap_8 FILLER_78_2380 ();
 sg13g2_fill_2 FILLER_78_2387 ();
 sg13g2_decap_8 FILLER_78_2393 ();
 sg13g2_decap_8 FILLER_78_2400 ();
 sg13g2_decap_8 FILLER_78_2407 ();
 sg13g2_decap_8 FILLER_78_2414 ();
 sg13g2_decap_8 FILLER_78_2421 ();
 sg13g2_decap_8 FILLER_78_2428 ();
 sg13g2_decap_8 FILLER_78_2435 ();
 sg13g2_decap_8 FILLER_78_2442 ();
 sg13g2_decap_8 FILLER_78_2449 ();
 sg13g2_decap_8 FILLER_78_2456 ();
 sg13g2_decap_8 FILLER_78_2463 ();
 sg13g2_decap_8 FILLER_78_2470 ();
 sg13g2_decap_8 FILLER_78_2477 ();
 sg13g2_decap_8 FILLER_78_2484 ();
 sg13g2_decap_8 FILLER_78_2491 ();
 sg13g2_decap_8 FILLER_78_2498 ();
 sg13g2_decap_8 FILLER_78_2505 ();
 sg13g2_decap_8 FILLER_78_2512 ();
 sg13g2_decap_8 FILLER_78_2519 ();
 sg13g2_decap_8 FILLER_78_2526 ();
 sg13g2_decap_8 FILLER_78_2533 ();
 sg13g2_decap_8 FILLER_78_2540 ();
 sg13g2_decap_8 FILLER_78_2547 ();
 sg13g2_decap_8 FILLER_78_2554 ();
 sg13g2_decap_8 FILLER_78_2561 ();
 sg13g2_decap_8 FILLER_78_2568 ();
 sg13g2_decap_8 FILLER_78_2575 ();
 sg13g2_decap_8 FILLER_78_2582 ();
 sg13g2_decap_8 FILLER_78_2589 ();
 sg13g2_decap_8 FILLER_78_2596 ();
 sg13g2_decap_8 FILLER_78_2603 ();
 sg13g2_decap_8 FILLER_78_2610 ();
 sg13g2_decap_8 FILLER_78_2617 ();
 sg13g2_decap_8 FILLER_78_2624 ();
 sg13g2_decap_8 FILLER_78_2631 ();
 sg13g2_decap_8 FILLER_78_2638 ();
 sg13g2_decap_8 FILLER_78_2645 ();
 sg13g2_decap_8 FILLER_78_2652 ();
 sg13g2_decap_8 FILLER_78_2659 ();
 sg13g2_decap_8 FILLER_78_2666 ();
 sg13g2_fill_1 FILLER_78_2673 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_4 FILLER_79_42 ();
 sg13g2_fill_1 FILLER_79_103 ();
 sg13g2_fill_1 FILLER_79_157 ();
 sg13g2_fill_1 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_302 ();
 sg13g2_fill_2 FILLER_79_367 ();
 sg13g2_fill_2 FILLER_79_410 ();
 sg13g2_fill_2 FILLER_79_444 ();
 sg13g2_fill_2 FILLER_79_590 ();
 sg13g2_fill_2 FILLER_79_620 ();
 sg13g2_fill_1 FILLER_79_622 ();
 sg13g2_decap_4 FILLER_79_632 ();
 sg13g2_fill_1 FILLER_79_636 ();
 sg13g2_fill_1 FILLER_79_660 ();
 sg13g2_fill_2 FILLER_79_763 ();
 sg13g2_decap_8 FILLER_79_769 ();
 sg13g2_decap_8 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_783 ();
 sg13g2_decap_4 FILLER_79_790 ();
 sg13g2_fill_2 FILLER_79_794 ();
 sg13g2_fill_2 FILLER_79_884 ();
 sg13g2_fill_1 FILLER_79_914 ();
 sg13g2_decap_8 FILLER_79_940 ();
 sg13g2_decap_8 FILLER_79_947 ();
 sg13g2_decap_4 FILLER_79_954 ();
 sg13g2_fill_1 FILLER_79_958 ();
 sg13g2_decap_8 FILLER_79_964 ();
 sg13g2_decap_8 FILLER_79_971 ();
 sg13g2_decap_4 FILLER_79_978 ();
 sg13g2_decap_8 FILLER_79_995 ();
 sg13g2_decap_8 FILLER_79_1002 ();
 sg13g2_fill_2 FILLER_79_1009 ();
 sg13g2_fill_1 FILLER_79_1011 ();
 sg13g2_decap_4 FILLER_79_1018 ();
 sg13g2_decap_8 FILLER_79_1031 ();
 sg13g2_decap_8 FILLER_79_1038 ();
 sg13g2_decap_4 FILLER_79_1045 ();
 sg13g2_decap_8 FILLER_79_1072 ();
 sg13g2_decap_8 FILLER_79_1079 ();
 sg13g2_decap_4 FILLER_79_1086 ();
 sg13g2_fill_1 FILLER_79_1121 ();
 sg13g2_decap_8 FILLER_79_1237 ();
 sg13g2_fill_1 FILLER_79_1244 ();
 sg13g2_decap_4 FILLER_79_1311 ();
 sg13g2_fill_2 FILLER_79_1395 ();
 sg13g2_fill_1 FILLER_79_1397 ();
 sg13g2_fill_2 FILLER_79_1425 ();
 sg13g2_fill_1 FILLER_79_1427 ();
 sg13g2_fill_1 FILLER_79_1482 ();
 sg13g2_fill_1 FILLER_79_1546 ();
 sg13g2_fill_2 FILLER_79_1658 ();
 sg13g2_fill_2 FILLER_79_1807 ();
 sg13g2_fill_2 FILLER_79_1846 ();
 sg13g2_fill_2 FILLER_79_1888 ();
 sg13g2_fill_1 FILLER_79_1985 ();
 sg13g2_decap_8 FILLER_79_2027 ();
 sg13g2_fill_2 FILLER_79_2074 ();
 sg13g2_decap_8 FILLER_79_2112 ();
 sg13g2_decap_8 FILLER_79_2119 ();
 sg13g2_decap_8 FILLER_79_2126 ();
 sg13g2_decap_8 FILLER_79_2133 ();
 sg13g2_decap_8 FILLER_79_2140 ();
 sg13g2_decap_8 FILLER_79_2147 ();
 sg13g2_decap_8 FILLER_79_2154 ();
 sg13g2_decap_8 FILLER_79_2161 ();
 sg13g2_decap_8 FILLER_79_2168 ();
 sg13g2_decap_8 FILLER_79_2175 ();
 sg13g2_decap_8 FILLER_79_2182 ();
 sg13g2_fill_2 FILLER_79_2189 ();
 sg13g2_fill_1 FILLER_79_2191 ();
 sg13g2_decap_4 FILLER_79_2224 ();
 sg13g2_fill_1 FILLER_79_2228 ();
 sg13g2_fill_1 FILLER_79_2237 ();
 sg13g2_decap_4 FILLER_79_2243 ();
 sg13g2_fill_2 FILLER_79_2247 ();
 sg13g2_decap_8 FILLER_79_2294 ();
 sg13g2_decap_8 FILLER_79_2301 ();
 sg13g2_decap_8 FILLER_79_2308 ();
 sg13g2_decap_8 FILLER_79_2315 ();
 sg13g2_decap_8 FILLER_79_2322 ();
 sg13g2_decap_8 FILLER_79_2329 ();
 sg13g2_decap_8 FILLER_79_2336 ();
 sg13g2_decap_8 FILLER_79_2343 ();
 sg13g2_decap_8 FILLER_79_2350 ();
 sg13g2_decap_8 FILLER_79_2357 ();
 sg13g2_decap_8 FILLER_79_2364 ();
 sg13g2_decap_8 FILLER_79_2371 ();
 sg13g2_decap_4 FILLER_79_2378 ();
 sg13g2_fill_2 FILLER_79_2382 ();
 sg13g2_decap_8 FILLER_79_2437 ();
 sg13g2_decap_8 FILLER_79_2444 ();
 sg13g2_decap_8 FILLER_79_2451 ();
 sg13g2_decap_8 FILLER_79_2458 ();
 sg13g2_decap_8 FILLER_79_2465 ();
 sg13g2_decap_8 FILLER_79_2472 ();
 sg13g2_decap_8 FILLER_79_2479 ();
 sg13g2_decap_8 FILLER_79_2486 ();
 sg13g2_decap_8 FILLER_79_2493 ();
 sg13g2_decap_8 FILLER_79_2500 ();
 sg13g2_decap_8 FILLER_79_2507 ();
 sg13g2_decap_8 FILLER_79_2514 ();
 sg13g2_decap_8 FILLER_79_2521 ();
 sg13g2_decap_8 FILLER_79_2528 ();
 sg13g2_decap_8 FILLER_79_2535 ();
 sg13g2_decap_8 FILLER_79_2542 ();
 sg13g2_decap_8 FILLER_79_2549 ();
 sg13g2_decap_8 FILLER_79_2556 ();
 sg13g2_decap_8 FILLER_79_2563 ();
 sg13g2_decap_8 FILLER_79_2570 ();
 sg13g2_decap_8 FILLER_79_2577 ();
 sg13g2_decap_8 FILLER_79_2584 ();
 sg13g2_decap_8 FILLER_79_2591 ();
 sg13g2_decap_8 FILLER_79_2598 ();
 sg13g2_decap_8 FILLER_79_2605 ();
 sg13g2_decap_8 FILLER_79_2612 ();
 sg13g2_decap_8 FILLER_79_2619 ();
 sg13g2_decap_8 FILLER_79_2626 ();
 sg13g2_decap_8 FILLER_79_2633 ();
 sg13g2_decap_8 FILLER_79_2640 ();
 sg13g2_decap_8 FILLER_79_2647 ();
 sg13g2_decap_8 FILLER_79_2654 ();
 sg13g2_decap_8 FILLER_79_2661 ();
 sg13g2_decap_4 FILLER_79_2668 ();
 sg13g2_fill_2 FILLER_79_2672 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_4 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_85 ();
 sg13g2_fill_1 FILLER_80_96 ();
 sg13g2_decap_8 FILLER_80_152 ();
 sg13g2_decap_8 FILLER_80_159 ();
 sg13g2_fill_2 FILLER_80_166 ();
 sg13g2_decap_4 FILLER_80_199 ();
 sg13g2_decap_4 FILLER_80_238 ();
 sg13g2_fill_2 FILLER_80_270 ();
 sg13g2_fill_2 FILLER_80_282 ();
 sg13g2_fill_1 FILLER_80_284 ();
 sg13g2_fill_2 FILLER_80_305 ();
 sg13g2_fill_1 FILLER_80_307 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_4 FILLER_80_377 ();
 sg13g2_fill_2 FILLER_80_381 ();
 sg13g2_decap_4 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_469 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_fill_2 FILLER_80_483 ();
 sg13g2_fill_1 FILLER_80_485 ();
 sg13g2_fill_2 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_532 ();
 sg13g2_decap_4 FILLER_80_539 ();
 sg13g2_fill_2 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_fill_1 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_fill_2 FILLER_80_618 ();
 sg13g2_decap_4 FILLER_80_628 ();
 sg13g2_fill_2 FILLER_80_632 ();
 sg13g2_fill_2 FILLER_80_648 ();
 sg13g2_fill_2 FILLER_80_659 ();
 sg13g2_fill_1 FILLER_80_671 ();
 sg13g2_fill_1 FILLER_80_702 ();
 sg13g2_fill_1 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_4 FILLER_80_790 ();
 sg13g2_fill_1 FILLER_80_794 ();
 sg13g2_fill_2 FILLER_80_822 ();
 sg13g2_fill_1 FILLER_80_824 ();
 sg13g2_fill_2 FILLER_80_852 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_decap_4 FILLER_80_898 ();
 sg13g2_fill_2 FILLER_80_902 ();
 sg13g2_decap_4 FILLER_80_917 ();
 sg13g2_fill_2 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_932 ();
 sg13g2_decap_8 FILLER_80_939 ();
 sg13g2_decap_8 FILLER_80_946 ();
 sg13g2_decap_8 FILLER_80_953 ();
 sg13g2_decap_8 FILLER_80_960 ();
 sg13g2_decap_8 FILLER_80_967 ();
 sg13g2_decap_8 FILLER_80_974 ();
 sg13g2_decap_8 FILLER_80_981 ();
 sg13g2_decap_8 FILLER_80_988 ();
 sg13g2_decap_8 FILLER_80_995 ();
 sg13g2_decap_8 FILLER_80_1002 ();
 sg13g2_decap_8 FILLER_80_1009 ();
 sg13g2_decap_8 FILLER_80_1016 ();
 sg13g2_decap_8 FILLER_80_1023 ();
 sg13g2_decap_8 FILLER_80_1030 ();
 sg13g2_decap_8 FILLER_80_1037 ();
 sg13g2_decap_8 FILLER_80_1044 ();
 sg13g2_decap_4 FILLER_80_1051 ();
 sg13g2_decap_8 FILLER_80_1060 ();
 sg13g2_decap_8 FILLER_80_1067 ();
 sg13g2_decap_8 FILLER_80_1074 ();
 sg13g2_decap_8 FILLER_80_1081 ();
 sg13g2_decap_8 FILLER_80_1088 ();
 sg13g2_decap_4 FILLER_80_1095 ();
 sg13g2_fill_1 FILLER_80_1156 ();
 sg13g2_fill_2 FILLER_80_1237 ();
 sg13g2_fill_1 FILLER_80_1289 ();
 sg13g2_decap_4 FILLER_80_1306 ();
 sg13g2_fill_2 FILLER_80_1310 ();
 sg13g2_fill_2 FILLER_80_1321 ();
 sg13g2_fill_1 FILLER_80_1323 ();
 sg13g2_decap_4 FILLER_80_1349 ();
 sg13g2_fill_2 FILLER_80_1353 ();
 sg13g2_fill_1 FILLER_80_1368 ();
 sg13g2_fill_1 FILLER_80_1387 ();
 sg13g2_fill_1 FILLER_80_1418 ();
 sg13g2_fill_1 FILLER_80_1428 ();
 sg13g2_fill_2 FILLER_80_1442 ();
 sg13g2_fill_2 FILLER_80_1507 ();
 sg13g2_fill_2 FILLER_80_1593 ();
 sg13g2_fill_1 FILLER_80_1613 ();
 sg13g2_fill_2 FILLER_80_1628 ();
 sg13g2_fill_2 FILLER_80_1683 ();
 sg13g2_fill_1 FILLER_80_1685 ();
 sg13g2_fill_2 FILLER_80_1713 ();
 sg13g2_fill_1 FILLER_80_1715 ();
 sg13g2_fill_1 FILLER_80_1812 ();
 sg13g2_fill_2 FILLER_80_1845 ();
 sg13g2_fill_2 FILLER_80_1875 ();
 sg13g2_fill_2 FILLER_80_1903 ();
 sg13g2_fill_2 FILLER_80_1910 ();
 sg13g2_fill_1 FILLER_80_1957 ();
 sg13g2_fill_2 FILLER_80_1976 ();
 sg13g2_fill_1 FILLER_80_1978 ();
 sg13g2_decap_8 FILLER_80_2026 ();
 sg13g2_fill_2 FILLER_80_2033 ();
 sg13g2_fill_2 FILLER_80_2045 ();
 sg13g2_decap_8 FILLER_80_2111 ();
 sg13g2_decap_8 FILLER_80_2118 ();
 sg13g2_decap_8 FILLER_80_2125 ();
 sg13g2_decap_8 FILLER_80_2132 ();
 sg13g2_decap_8 FILLER_80_2139 ();
 sg13g2_decap_8 FILLER_80_2146 ();
 sg13g2_decap_8 FILLER_80_2153 ();
 sg13g2_decap_8 FILLER_80_2160 ();
 sg13g2_decap_8 FILLER_80_2167 ();
 sg13g2_decap_8 FILLER_80_2174 ();
 sg13g2_decap_8 FILLER_80_2181 ();
 sg13g2_decap_8 FILLER_80_2188 ();
 sg13g2_decap_8 FILLER_80_2195 ();
 sg13g2_fill_1 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2231 ();
 sg13g2_decap_8 FILLER_80_2238 ();
 sg13g2_decap_8 FILLER_80_2245 ();
 sg13g2_decap_8 FILLER_80_2252 ();
 sg13g2_fill_2 FILLER_80_2259 ();
 sg13g2_fill_2 FILLER_80_2265 ();
 sg13g2_decap_8 FILLER_80_2276 ();
 sg13g2_decap_8 FILLER_80_2283 ();
 sg13g2_decap_8 FILLER_80_2290 ();
 sg13g2_decap_8 FILLER_80_2297 ();
 sg13g2_decap_8 FILLER_80_2304 ();
 sg13g2_decap_8 FILLER_80_2311 ();
 sg13g2_decap_8 FILLER_80_2318 ();
 sg13g2_decap_8 FILLER_80_2325 ();
 sg13g2_decap_8 FILLER_80_2332 ();
 sg13g2_decap_8 FILLER_80_2339 ();
 sg13g2_decap_8 FILLER_80_2346 ();
 sg13g2_decap_8 FILLER_80_2353 ();
 sg13g2_decap_8 FILLER_80_2360 ();
 sg13g2_decap_8 FILLER_80_2367 ();
 sg13g2_decap_8 FILLER_80_2374 ();
 sg13g2_decap_8 FILLER_80_2381 ();
 sg13g2_decap_8 FILLER_80_2388 ();
 sg13g2_decap_8 FILLER_80_2395 ();
 sg13g2_decap_8 FILLER_80_2402 ();
 sg13g2_decap_8 FILLER_80_2409 ();
 sg13g2_decap_8 FILLER_80_2416 ();
 sg13g2_decap_8 FILLER_80_2423 ();
 sg13g2_decap_8 FILLER_80_2430 ();
 sg13g2_decap_8 FILLER_80_2437 ();
 sg13g2_decap_8 FILLER_80_2444 ();
 sg13g2_decap_8 FILLER_80_2451 ();
 sg13g2_decap_8 FILLER_80_2458 ();
 sg13g2_decap_8 FILLER_80_2465 ();
 sg13g2_decap_8 FILLER_80_2472 ();
 sg13g2_decap_8 FILLER_80_2479 ();
 sg13g2_decap_8 FILLER_80_2486 ();
 sg13g2_decap_8 FILLER_80_2493 ();
 sg13g2_decap_8 FILLER_80_2500 ();
 sg13g2_decap_8 FILLER_80_2507 ();
 sg13g2_decap_8 FILLER_80_2514 ();
 sg13g2_decap_8 FILLER_80_2521 ();
 sg13g2_decap_8 FILLER_80_2528 ();
 sg13g2_decap_8 FILLER_80_2535 ();
 sg13g2_decap_8 FILLER_80_2542 ();
 sg13g2_decap_8 FILLER_80_2549 ();
 sg13g2_decap_8 FILLER_80_2556 ();
 sg13g2_decap_8 FILLER_80_2563 ();
 sg13g2_decap_8 FILLER_80_2570 ();
 sg13g2_decap_8 FILLER_80_2577 ();
 sg13g2_decap_8 FILLER_80_2584 ();
 sg13g2_decap_8 FILLER_80_2591 ();
 sg13g2_decap_8 FILLER_80_2598 ();
 sg13g2_decap_8 FILLER_80_2605 ();
 sg13g2_decap_8 FILLER_80_2612 ();
 sg13g2_decap_8 FILLER_80_2619 ();
 sg13g2_decap_8 FILLER_80_2626 ();
 sg13g2_decap_8 FILLER_80_2633 ();
 sg13g2_decap_8 FILLER_80_2640 ();
 sg13g2_decap_8 FILLER_80_2647 ();
 sg13g2_decap_8 FILLER_80_2654 ();
 sg13g2_decap_8 FILLER_80_2661 ();
 sg13g2_decap_4 FILLER_80_2668 ();
 sg13g2_fill_2 FILLER_80_2672 ();
 assign uio_oe[0] = net76;
 assign uio_oe[3] = net77;
 assign uio_oe[6] = net78;
endmodule
