module tt_um_chrismoos_led_controller (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire clknet_leaf_0_clk;
 wire \led_controller.clock_divider[0] ;
 wire \led_controller.clock_divider[1] ;
 wire \led_controller.clock_divider[2] ;
 wire \led_controller.clock_divider[3] ;
 wire \led_controller.clock_divider[4] ;
 wire \led_controller.clock_divider[5] ;
 wire \led_controller.clock_divider[6] ;
 wire \led_controller.clock_divider[7] ;
 wire \led_controller.colors[0] ;
 wire \led_controller.colors[10] ;
 wire \led_controller.colors[11] ;
 wire \led_controller.colors[12] ;
 wire \led_controller.colors[13] ;
 wire \led_controller.colors[14] ;
 wire \led_controller.colors[15] ;
 wire \led_controller.colors[16] ;
 wire \led_controller.colors[17] ;
 wire \led_controller.colors[18] ;
 wire \led_controller.colors[19] ;
 wire \led_controller.colors[1] ;
 wire \led_controller.colors[20] ;
 wire \led_controller.colors[21] ;
 wire \led_controller.colors[22] ;
 wire \led_controller.colors[23] ;
 wire \led_controller.colors[24] ;
 wire \led_controller.colors[25] ;
 wire \led_controller.colors[26] ;
 wire \led_controller.colors[27] ;
 wire \led_controller.colors[28] ;
 wire \led_controller.colors[29] ;
 wire \led_controller.colors[2] ;
 wire \led_controller.colors[30] ;
 wire \led_controller.colors[31] ;
 wire \led_controller.colors[32] ;
 wire \led_controller.colors[33] ;
 wire \led_controller.colors[34] ;
 wire \led_controller.colors[35] ;
 wire \led_controller.colors[36] ;
 wire \led_controller.colors[37] ;
 wire \led_controller.colors[38] ;
 wire \led_controller.colors[39] ;
 wire \led_controller.colors[3] ;
 wire \led_controller.colors[40] ;
 wire \led_controller.colors[41] ;
 wire \led_controller.colors[42] ;
 wire \led_controller.colors[43] ;
 wire \led_controller.colors[44] ;
 wire \led_controller.colors[45] ;
 wire \led_controller.colors[46] ;
 wire \led_controller.colors[47] ;
 wire \led_controller.colors[48] ;
 wire \led_controller.colors[49] ;
 wire \led_controller.colors[4] ;
 wire \led_controller.colors[50] ;
 wire \led_controller.colors[51] ;
 wire \led_controller.colors[52] ;
 wire \led_controller.colors[53] ;
 wire \led_controller.colors[54] ;
 wire \led_controller.colors[55] ;
 wire \led_controller.colors[56] ;
 wire \led_controller.colors[57] ;
 wire \led_controller.colors[58] ;
 wire \led_controller.colors[59] ;
 wire \led_controller.colors[5] ;
 wire \led_controller.colors[60] ;
 wire \led_controller.colors[61] ;
 wire \led_controller.colors[62] ;
 wire \led_controller.colors[63] ;
 wire \led_controller.colors[64] ;
 wire \led_controller.colors[65] ;
 wire \led_controller.colors[66] ;
 wire \led_controller.colors[67] ;
 wire \led_controller.colors[68] ;
 wire \led_controller.colors[69] ;
 wire \led_controller.colors[6] ;
 wire \led_controller.colors[70] ;
 wire \led_controller.colors[71] ;
 wire \led_controller.colors[72] ;
 wire \led_controller.colors[73] ;
 wire \led_controller.colors[74] ;
 wire \led_controller.colors[75] ;
 wire \led_controller.colors[76] ;
 wire \led_controller.colors[77] ;
 wire \led_controller.colors[78] ;
 wire \led_controller.colors[79] ;
 wire \led_controller.colors[7] ;
 wire \led_controller.colors[80] ;
 wire \led_controller.colors[81] ;
 wire \led_controller.colors[82] ;
 wire \led_controller.colors[83] ;
 wire \led_controller.colors[84] ;
 wire \led_controller.colors[85] ;
 wire \led_controller.colors[86] ;
 wire \led_controller.colors[87] ;
 wire \led_controller.colors[88] ;
 wire \led_controller.colors[89] ;
 wire \led_controller.colors[8] ;
 wire \led_controller.colors[90] ;
 wire \led_controller.colors[91] ;
 wire \led_controller.colors[92] ;
 wire \led_controller.colors[93] ;
 wire \led_controller.colors[94] ;
 wire \led_controller.colors[95] ;
 wire \led_controller.colors[9] ;
 wire \led_controller.cpu.bus_hi_valid ;
 wire \led_controller.cpu.current_instruction[0] ;
 wire \led_controller.cpu.current_instruction[10] ;
 wire \led_controller.cpu.current_instruction[11] ;
 wire \led_controller.cpu.current_instruction[12] ;
 wire \led_controller.cpu.current_instruction[13] ;
 wire \led_controller.cpu.current_instruction[14] ;
 wire \led_controller.cpu.current_instruction[15] ;
 wire \led_controller.cpu.current_instruction[1] ;
 wire \led_controller.cpu.current_instruction[2] ;
 wire \led_controller.cpu.current_instruction[3] ;
 wire \led_controller.cpu.current_instruction[4] ;
 wire \led_controller.cpu.current_instruction[5] ;
 wire \led_controller.cpu.current_instruction[6] ;
 wire \led_controller.cpu.current_instruction[7] ;
 wire \led_controller.cpu.current_instruction[8] ;
 wire \led_controller.cpu.current_instruction[9] ;
 wire \led_controller.cpu.current_instruction_pc[0] ;
 wire \led_controller.cpu.current_instruction_pc[10] ;
 wire \led_controller.cpu.current_instruction_pc[11] ;
 wire \led_controller.cpu.current_instruction_pc[12] ;
 wire \led_controller.cpu.current_instruction_pc[13] ;
 wire \led_controller.cpu.current_instruction_pc[14] ;
 wire \led_controller.cpu.current_instruction_pc[15] ;
 wire \led_controller.cpu.current_instruction_pc[1] ;
 wire \led_controller.cpu.current_instruction_pc[2] ;
 wire \led_controller.cpu.current_instruction_pc[3] ;
 wire \led_controller.cpu.current_instruction_pc[4] ;
 wire \led_controller.cpu.current_instruction_pc[5] ;
 wire \led_controller.cpu.current_instruction_pc[6] ;
 wire \led_controller.cpu.current_instruction_pc[7] ;
 wire \led_controller.cpu.current_instruction_pc[8] ;
 wire \led_controller.cpu.current_instruction_pc[9] ;
 wire \led_controller.cpu.current_instruction_valid ;
 wire \led_controller.cpu.fetch_instruction[0] ;
 wire \led_controller.cpu.fetch_instruction[10] ;
 wire \led_controller.cpu.fetch_instruction[11] ;
 wire \led_controller.cpu.fetch_instruction[12] ;
 wire \led_controller.cpu.fetch_instruction[13] ;
 wire \led_controller.cpu.fetch_instruction[14] ;
 wire \led_controller.cpu.fetch_instruction[15] ;
 wire \led_controller.cpu.fetch_instruction[1] ;
 wire \led_controller.cpu.fetch_instruction[2] ;
 wire \led_controller.cpu.fetch_instruction[3] ;
 wire \led_controller.cpu.fetch_instruction[4] ;
 wire \led_controller.cpu.fetch_instruction[5] ;
 wire \led_controller.cpu.fetch_instruction[6] ;
 wire \led_controller.cpu.fetch_instruction[7] ;
 wire \led_controller.cpu.fetch_instruction[8] ;
 wire \led_controller.cpu.fetch_instruction[9] ;
 wire \led_controller.cpu.fetch_pc[0] ;
 wire \led_controller.cpu.fetch_pc[10] ;
 wire \led_controller.cpu.fetch_pc[11] ;
 wire \led_controller.cpu.fetch_pc[12] ;
 wire \led_controller.cpu.fetch_pc[13] ;
 wire \led_controller.cpu.fetch_pc[14] ;
 wire \led_controller.cpu.fetch_pc[15] ;
 wire \led_controller.cpu.fetch_pc[1] ;
 wire \led_controller.cpu.fetch_pc[2] ;
 wire \led_controller.cpu.fetch_pc[3] ;
 wire \led_controller.cpu.fetch_pc[4] ;
 wire \led_controller.cpu.fetch_pc[5] ;
 wire \led_controller.cpu.fetch_pc[6] ;
 wire \led_controller.cpu.fetch_pc[7] ;
 wire \led_controller.cpu.fetch_pc[8] ;
 wire \led_controller.cpu.fetch_pc[9] ;
 wire \led_controller.cpu.fetch_pc_valid ;
 wire \led_controller.cpu.i_bus_data[0] ;
 wire \led_controller.cpu.i_bus_data[1] ;
 wire \led_controller.cpu.i_bus_data[2] ;
 wire \led_controller.cpu.i_bus_data[3] ;
 wire \led_controller.cpu.i_bus_data[4] ;
 wire \led_controller.cpu.i_bus_data[5] ;
 wire \led_controller.cpu.i_bus_data[6] ;
 wire \led_controller.cpu.i_bus_data[7] ;
 wire \led_controller.cpu.i_bus_data_valid ;
 wire \led_controller.cpu.i_num_colors[0] ;
 wire \led_controller.cpu.i_num_colors[1] ;
 wire \led_controller.cpu.i_num_leds[0] ;
 wire \led_controller.cpu.i_num_leds[1] ;
 wire \led_controller.cpu.i_num_leds[2] ;
 wire \led_controller.cpu.i_num_leds[3] ;
 wire \led_controller.cpu.i_num_leds[4] ;
 wire \led_controller.cpu.i_num_leds[5] ;
 wire \led_controller.cpu.i_num_leds[6] ;
 wire \led_controller.cpu.i_num_leds[7] ;
 wire \led_controller.cpu.i_timer_100hz ;
 wire \led_controller.cpu.led_write_color[0] ;
 wire \led_controller.cpu.led_write_color[1] ;
 wire \led_controller.cpu.led_write_pending ;
 wire \led_controller.cpu.led_write_strb ;
 wire \led_controller.cpu.led_writing ;
 wire \led_controller.cpu.o_bus_addr[0] ;
 wire \led_controller.cpu.o_bus_addr[10] ;
 wire \led_controller.cpu.o_bus_addr[11] ;
 wire \led_controller.cpu.o_bus_addr[12] ;
 wire \led_controller.cpu.o_bus_addr[13] ;
 wire \led_controller.cpu.o_bus_addr[14] ;
 wire \led_controller.cpu.o_bus_addr[15] ;
 wire \led_controller.cpu.o_bus_addr[1] ;
 wire \led_controller.cpu.o_bus_addr[2] ;
 wire \led_controller.cpu.o_bus_addr[3] ;
 wire \led_controller.cpu.o_bus_addr[4] ;
 wire \led_controller.cpu.o_bus_addr[5] ;
 wire \led_controller.cpu.o_bus_addr[6] ;
 wire \led_controller.cpu.o_bus_addr[7] ;
 wire \led_controller.cpu.o_bus_addr[8] ;
 wire \led_controller.cpu.o_bus_addr[9] ;
 wire \led_controller.cpu.o_bus_addr_valid ;
 wire \led_controller.cpu.o_led_color[0] ;
 wire \led_controller.cpu.o_led_color[1] ;
 wire \led_controller.cpu.o_led_strb ;
 wire \led_controller.cpu.pc[0] ;
 wire \led_controller.cpu.pc[10] ;
 wire \led_controller.cpu.pc[11] ;
 wire \led_controller.cpu.pc[12] ;
 wire \led_controller.cpu.pc[13] ;
 wire \led_controller.cpu.pc[14] ;
 wire \led_controller.cpu.pc[15] ;
 wire \led_controller.cpu.pc[1] ;
 wire \led_controller.cpu.pc[2] ;
 wire \led_controller.cpu.pc[3] ;
 wire \led_controller.cpu.pc[4] ;
 wire \led_controller.cpu.pc[5] ;
 wire \led_controller.cpu.pc[6] ;
 wire \led_controller.cpu.pc[7] ;
 wire \led_controller.cpu.pc[8] ;
 wire \led_controller.cpu.pc[9] ;
 wire \led_controller.cpu.register_x[0] ;
 wire \led_controller.cpu.register_x[1] ;
 wire \led_controller.cpu.register_x[2] ;
 wire \led_controller.cpu.register_x[3] ;
 wire \led_controller.cpu.register_x[4] ;
 wire \led_controller.cpu.register_x[5] ;
 wire \led_controller.cpu.register_x[6] ;
 wire \led_controller.cpu.register_x[7] ;
 wire \led_controller.cpu.register_y[0] ;
 wire \led_controller.cpu.register_y[1] ;
 wire \led_controller.cpu.register_y[2] ;
 wire \led_controller.cpu.register_y[3] ;
 wire \led_controller.cpu.register_y[4] ;
 wire \led_controller.cpu.register_y[5] ;
 wire \led_controller.cpu.register_y[6] ;
 wire \led_controller.cpu.register_y[7] ;
 wire \led_controller.cpu.scratch_memory[0][0] ;
 wire \led_controller.cpu.scratch_memory[0][1] ;
 wire \led_controller.cpu.scratch_memory[0][2] ;
 wire \led_controller.cpu.scratch_memory[0][3] ;
 wire \led_controller.cpu.scratch_memory[0][4] ;
 wire \led_controller.cpu.scratch_memory[0][5] ;
 wire \led_controller.cpu.scratch_memory[0][6] ;
 wire \led_controller.cpu.scratch_memory[0][7] ;
 wire \led_controller.cpu.scratch_memory[10][0] ;
 wire \led_controller.cpu.scratch_memory[10][1] ;
 wire \led_controller.cpu.scratch_memory[10][2] ;
 wire \led_controller.cpu.scratch_memory[10][3] ;
 wire \led_controller.cpu.scratch_memory[10][4] ;
 wire \led_controller.cpu.scratch_memory[10][5] ;
 wire \led_controller.cpu.scratch_memory[10][6] ;
 wire \led_controller.cpu.scratch_memory[10][7] ;
 wire \led_controller.cpu.scratch_memory[11][0] ;
 wire \led_controller.cpu.scratch_memory[11][1] ;
 wire \led_controller.cpu.scratch_memory[11][2] ;
 wire \led_controller.cpu.scratch_memory[11][3] ;
 wire \led_controller.cpu.scratch_memory[11][4] ;
 wire \led_controller.cpu.scratch_memory[11][5] ;
 wire \led_controller.cpu.scratch_memory[11][6] ;
 wire \led_controller.cpu.scratch_memory[11][7] ;
 wire \led_controller.cpu.scratch_memory[12][0] ;
 wire \led_controller.cpu.scratch_memory[12][1] ;
 wire \led_controller.cpu.scratch_memory[12][2] ;
 wire \led_controller.cpu.scratch_memory[12][3] ;
 wire \led_controller.cpu.scratch_memory[12][4] ;
 wire \led_controller.cpu.scratch_memory[12][5] ;
 wire \led_controller.cpu.scratch_memory[12][6] ;
 wire \led_controller.cpu.scratch_memory[12][7] ;
 wire \led_controller.cpu.scratch_memory[13][0] ;
 wire \led_controller.cpu.scratch_memory[13][1] ;
 wire \led_controller.cpu.scratch_memory[13][2] ;
 wire \led_controller.cpu.scratch_memory[13][3] ;
 wire \led_controller.cpu.scratch_memory[13][4] ;
 wire \led_controller.cpu.scratch_memory[13][5] ;
 wire \led_controller.cpu.scratch_memory[13][6] ;
 wire \led_controller.cpu.scratch_memory[13][7] ;
 wire \led_controller.cpu.scratch_memory[14][0] ;
 wire \led_controller.cpu.scratch_memory[14][1] ;
 wire \led_controller.cpu.scratch_memory[14][2] ;
 wire \led_controller.cpu.scratch_memory[14][3] ;
 wire \led_controller.cpu.scratch_memory[14][4] ;
 wire \led_controller.cpu.scratch_memory[14][5] ;
 wire \led_controller.cpu.scratch_memory[14][6] ;
 wire \led_controller.cpu.scratch_memory[14][7] ;
 wire \led_controller.cpu.scratch_memory[15][0] ;
 wire \led_controller.cpu.scratch_memory[15][1] ;
 wire \led_controller.cpu.scratch_memory[15][2] ;
 wire \led_controller.cpu.scratch_memory[15][3] ;
 wire \led_controller.cpu.scratch_memory[15][4] ;
 wire \led_controller.cpu.scratch_memory[15][5] ;
 wire \led_controller.cpu.scratch_memory[15][6] ;
 wire \led_controller.cpu.scratch_memory[15][7] ;
 wire \led_controller.cpu.scratch_memory[1][0] ;
 wire \led_controller.cpu.scratch_memory[1][1] ;
 wire \led_controller.cpu.scratch_memory[1][2] ;
 wire \led_controller.cpu.scratch_memory[1][3] ;
 wire \led_controller.cpu.scratch_memory[1][4] ;
 wire \led_controller.cpu.scratch_memory[1][5] ;
 wire \led_controller.cpu.scratch_memory[1][6] ;
 wire \led_controller.cpu.scratch_memory[1][7] ;
 wire \led_controller.cpu.scratch_memory[2][0] ;
 wire \led_controller.cpu.scratch_memory[2][1] ;
 wire \led_controller.cpu.scratch_memory[2][2] ;
 wire \led_controller.cpu.scratch_memory[2][3] ;
 wire \led_controller.cpu.scratch_memory[2][4] ;
 wire \led_controller.cpu.scratch_memory[2][5] ;
 wire \led_controller.cpu.scratch_memory[2][6] ;
 wire \led_controller.cpu.scratch_memory[2][7] ;
 wire \led_controller.cpu.scratch_memory[3][0] ;
 wire \led_controller.cpu.scratch_memory[3][1] ;
 wire \led_controller.cpu.scratch_memory[3][2] ;
 wire \led_controller.cpu.scratch_memory[3][3] ;
 wire \led_controller.cpu.scratch_memory[3][4] ;
 wire \led_controller.cpu.scratch_memory[3][5] ;
 wire \led_controller.cpu.scratch_memory[3][6] ;
 wire \led_controller.cpu.scratch_memory[3][7] ;
 wire \led_controller.cpu.scratch_memory[4][0] ;
 wire \led_controller.cpu.scratch_memory[4][1] ;
 wire \led_controller.cpu.scratch_memory[4][2] ;
 wire \led_controller.cpu.scratch_memory[4][3] ;
 wire \led_controller.cpu.scratch_memory[4][4] ;
 wire \led_controller.cpu.scratch_memory[4][5] ;
 wire \led_controller.cpu.scratch_memory[4][6] ;
 wire \led_controller.cpu.scratch_memory[4][7] ;
 wire \led_controller.cpu.scratch_memory[5][0] ;
 wire \led_controller.cpu.scratch_memory[5][1] ;
 wire \led_controller.cpu.scratch_memory[5][2] ;
 wire \led_controller.cpu.scratch_memory[5][3] ;
 wire \led_controller.cpu.scratch_memory[5][4] ;
 wire \led_controller.cpu.scratch_memory[5][5] ;
 wire \led_controller.cpu.scratch_memory[5][6] ;
 wire \led_controller.cpu.scratch_memory[5][7] ;
 wire \led_controller.cpu.scratch_memory[6][0] ;
 wire \led_controller.cpu.scratch_memory[6][1] ;
 wire \led_controller.cpu.scratch_memory[6][2] ;
 wire \led_controller.cpu.scratch_memory[6][3] ;
 wire \led_controller.cpu.scratch_memory[6][4] ;
 wire \led_controller.cpu.scratch_memory[6][5] ;
 wire \led_controller.cpu.scratch_memory[6][6] ;
 wire \led_controller.cpu.scratch_memory[6][7] ;
 wire \led_controller.cpu.scratch_memory[7][0] ;
 wire \led_controller.cpu.scratch_memory[7][1] ;
 wire \led_controller.cpu.scratch_memory[7][2] ;
 wire \led_controller.cpu.scratch_memory[7][3] ;
 wire \led_controller.cpu.scratch_memory[7][4] ;
 wire \led_controller.cpu.scratch_memory[7][5] ;
 wire \led_controller.cpu.scratch_memory[7][6] ;
 wire \led_controller.cpu.scratch_memory[7][7] ;
 wire \led_controller.cpu.scratch_memory[8][0] ;
 wire \led_controller.cpu.scratch_memory[8][1] ;
 wire \led_controller.cpu.scratch_memory[8][2] ;
 wire \led_controller.cpu.scratch_memory[8][3] ;
 wire \led_controller.cpu.scratch_memory[8][4] ;
 wire \led_controller.cpu.scratch_memory[8][5] ;
 wire \led_controller.cpu.scratch_memory[8][6] ;
 wire \led_controller.cpu.scratch_memory[8][7] ;
 wire \led_controller.cpu.scratch_memory[9][0] ;
 wire \led_controller.cpu.scratch_memory[9][1] ;
 wire \led_controller.cpu.scratch_memory[9][2] ;
 wire \led_controller.cpu.scratch_memory[9][3] ;
 wire \led_controller.cpu.scratch_memory[9][4] ;
 wire \led_controller.cpu.scratch_memory[9][5] ;
 wire \led_controller.cpu.scratch_memory[9][6] ;
 wire \led_controller.cpu.scratch_memory[9][7] ;
 wire \led_controller.cpu.stall_counter[0] ;
 wire \led_controller.cpu.stall_counter[1] ;
 wire \led_controller.cpu.stall_counter[2] ;
 wire \led_controller.cpu.stall_counter[3] ;
 wire \led_controller.cpu.stall_counter[4] ;
 wire \led_controller.cpu.stall_counter[5] ;
 wire \led_controller.cpu.stall_counter[6] ;
 wire \led_controller.cpu.stall_counter[7] ;
 wire \led_controller.cpu.status_negative ;
 wire \led_controller.cpu.status_zero ;
 wire \led_controller.cpu_reset_counter[0] ;
 wire \led_controller.cpu_reset_counter[1] ;
 wire \led_controller.cpu_reset_counter[2] ;
 wire \led_controller.cpu_reset_counter[3] ;
 wire \led_controller.effect[0] ;
 wire \led_controller.effect[1] ;
 wire \led_controller.effect[2] ;
 wire \led_controller.effect[3] ;
 wire \led_controller.effect_chase_led_color[0] ;
 wire \led_controller.effect_chase_led_color[1] ;
 wire \led_controller.effect_chase_led_strb ;
 wire \led_controller.effect_pulse_led_color[0] ;
 wire \led_controller.effect_pulse_led_color[10] ;
 wire \led_controller.effect_pulse_led_color[11] ;
 wire \led_controller.effect_pulse_led_color[12] ;
 wire \led_controller.effect_pulse_led_color[13] ;
 wire \led_controller.effect_pulse_led_color[14] ;
 wire \led_controller.effect_pulse_led_color[15] ;
 wire \led_controller.effect_pulse_led_color[16] ;
 wire \led_controller.effect_pulse_led_color[17] ;
 wire \led_controller.effect_pulse_led_color[18] ;
 wire \led_controller.effect_pulse_led_color[19] ;
 wire \led_controller.effect_pulse_led_color[1] ;
 wire \led_controller.effect_pulse_led_color[20] ;
 wire \led_controller.effect_pulse_led_color[21] ;
 wire \led_controller.effect_pulse_led_color[22] ;
 wire \led_controller.effect_pulse_led_color[23] ;
 wire \led_controller.effect_pulse_led_color[24] ;
 wire \led_controller.effect_pulse_led_color[25] ;
 wire \led_controller.effect_pulse_led_color[26] ;
 wire \led_controller.effect_pulse_led_color[27] ;
 wire \led_controller.effect_pulse_led_color[28] ;
 wire \led_controller.effect_pulse_led_color[29] ;
 wire \led_controller.effect_pulse_led_color[2] ;
 wire \led_controller.effect_pulse_led_color[30] ;
 wire \led_controller.effect_pulse_led_color[31] ;
 wire \led_controller.effect_pulse_led_color[3] ;
 wire \led_controller.effect_pulse_led_color[4] ;
 wire \led_controller.effect_pulse_led_color[5] ;
 wire \led_controller.effect_pulse_led_color[6] ;
 wire \led_controller.effect_pulse_led_color[7] ;
 wire \led_controller.effect_pulse_led_color[8] ;
 wire \led_controller.effect_pulse_led_color[9] ;
 wire \led_controller.effect_pulse_led_strb ;
 wire \led_controller.flash.addr[0] ;
 wire \led_controller.flash.addr[10] ;
 wire \led_controller.flash.addr[11] ;
 wire \led_controller.flash.addr[12] ;
 wire \led_controller.flash.addr[13] ;
 wire \led_controller.flash.addr[14] ;
 wire \led_controller.flash.addr[15] ;
 wire \led_controller.flash.addr[1] ;
 wire \led_controller.flash.addr[2] ;
 wire \led_controller.flash.addr[3] ;
 wire \led_controller.flash.addr[4] ;
 wire \led_controller.flash.addr[5] ;
 wire \led_controller.flash.addr[6] ;
 wire \led_controller.flash.addr[7] ;
 wire \led_controller.flash.addr[8] ;
 wire \led_controller.flash.addr[9] ;
 wire \led_controller.flash.cs_delay_counter[0] ;
 wire \led_controller.flash.cs_delay_counter[1] ;
 wire \led_controller.flash.cs_delay_counter[2] ;
 wire \led_controller.flash.cs_delay_counter[3] ;
 wire \led_controller.flash.cs_delay_counter[4] ;
 wire \led_controller.flash.cs_delay_counter[5] ;
 wire \led_controller.flash.cs_delay_counter[6] ;
 wire \led_controller.flash.cs_delay_counter[7] ;
 wire \led_controller.flash.i_addr_width_24 ;
 wire \led_controller.flash.master.active ;
 wire \led_controller.flash.master.bit_counter[0] ;
 wire \led_controller.flash.master.bit_counter[1] ;
 wire \led_controller.flash.master.bit_counter[2] ;
 wire \led_controller.flash.master.bit_counter[3] ;
 wire \led_controller.flash.master.i_tx_data[0] ;
 wire \led_controller.flash.master.i_tx_data[1] ;
 wire \led_controller.flash.master.i_tx_data[2] ;
 wire \led_controller.flash.master.i_tx_data[3] ;
 wire \led_controller.flash.master.i_tx_data[4] ;
 wire \led_controller.flash.master.i_tx_data[5] ;
 wire \led_controller.flash.master.i_tx_data[6] ;
 wire \led_controller.flash.master.i_tx_data[7] ;
 wire \led_controller.flash.master.o_busy ;
 wire \led_controller.flash.master.o_mosi ;
 wire \led_controller.flash.master.o_rx_data_valid ;
 wire \led_controller.flash.master.o_sck ;
 wire \led_controller.flash.master.sck ;
 wire \led_controller.flash.master.sck_counter[0] ;
 wire \led_controller.flash.master.sck_counter[1] ;
 wire \led_controller.flash.master.sck_counter[2] ;
 wire \led_controller.flash.master.sck_counter[3] ;
 wire \led_controller.flash.master.sck_counter[4] ;
 wire \led_controller.flash.master.sck_counter[5] ;
 wire \led_controller.flash.master.sck_counter[6] ;
 wire \led_controller.flash.master.sck_counter[7] ;
 wire \led_controller.flash.master.tx_data[0] ;
 wire \led_controller.flash.master.tx_data[1] ;
 wire \led_controller.flash.master.tx_data[2] ;
 wire \led_controller.flash.master.tx_data[3] ;
 wire \led_controller.flash.master.tx_data[4] ;
 wire \led_controller.flash.master.tx_data[5] ;
 wire \led_controller.flash.master.tx_data[6] ;
 wire \led_controller.flash.master.tx_data[7] ;
 wire \led_controller.flash.o_cs_n ;
 wire \led_controller.flash.state[0] ;
 wire \led_controller.flash.state[1] ;
 wire \led_controller.flash.state[2] ;
 wire \led_controller.flash.state[3] ;
 wire \led_controller.flash.state[4] ;
 wire \led_controller.flash.state[5] ;
 wire \led_controller.flash.state[6] ;
 wire \led_controller.led_effect_chase.current_led[0] ;
 wire \led_controller.led_effect_chase.current_led[1] ;
 wire \led_controller.led_effect_chase.current_led[2] ;
 wire \led_controller.led_effect_chase.current_led[3] ;
 wire \led_controller.led_effect_chase.current_led[4] ;
 wire \led_controller.led_effect_chase.current_led[5] ;
 wire \led_controller.led_effect_chase.current_led[6] ;
 wire \led_controller.led_effect_chase.current_led[7] ;
 wire \led_controller.led_effect_chase.finished ;
 wire \led_controller.led_effect_chase.i_reset_n ;
 wire \led_controller.led_effect_pulse.brightness[0] ;
 wire \led_controller.led_effect_pulse.brightness[1] ;
 wire \led_controller.led_effect_pulse.brightness[2] ;
 wire \led_controller.led_effect_pulse.brightness[3] ;
 wire \led_controller.led_effect_pulse.brightness[4] ;
 wire \led_controller.led_effect_pulse.calc_color_out[0] ;
 wire \led_controller.led_effect_pulse.calc_color_out[10] ;
 wire \led_controller.led_effect_pulse.calc_color_out[11] ;
 wire \led_controller.led_effect_pulse.calc_color_out[12] ;
 wire \led_controller.led_effect_pulse.calc_color_out[13] ;
 wire \led_controller.led_effect_pulse.calc_color_out[14] ;
 wire \led_controller.led_effect_pulse.calc_color_out[15] ;
 wire \led_controller.led_effect_pulse.calc_color_out[16] ;
 wire \led_controller.led_effect_pulse.calc_color_out[17] ;
 wire \led_controller.led_effect_pulse.calc_color_out[18] ;
 wire \led_controller.led_effect_pulse.calc_color_out[19] ;
 wire \led_controller.led_effect_pulse.calc_color_out[1] ;
 wire \led_controller.led_effect_pulse.calc_color_out[20] ;
 wire \led_controller.led_effect_pulse.calc_color_out[21] ;
 wire \led_controller.led_effect_pulse.calc_color_out[22] ;
 wire \led_controller.led_effect_pulse.calc_color_out[23] ;
 wire \led_controller.led_effect_pulse.calc_color_out[24] ;
 wire \led_controller.led_effect_pulse.calc_color_out[25] ;
 wire \led_controller.led_effect_pulse.calc_color_out[26] ;
 wire \led_controller.led_effect_pulse.calc_color_out[27] ;
 wire \led_controller.led_effect_pulse.calc_color_out[28] ;
 wire \led_controller.led_effect_pulse.calc_color_out[29] ;
 wire \led_controller.led_effect_pulse.calc_color_out[2] ;
 wire \led_controller.led_effect_pulse.calc_color_out[30] ;
 wire \led_controller.led_effect_pulse.calc_color_out[31] ;
 wire \led_controller.led_effect_pulse.calc_color_out[3] ;
 wire \led_controller.led_effect_pulse.calc_color_out[4] ;
 wire \led_controller.led_effect_pulse.calc_color_out[5] ;
 wire \led_controller.led_effect_pulse.calc_color_out[6] ;
 wire \led_controller.led_effect_pulse.calc_color_out[7] ;
 wire \led_controller.led_effect_pulse.calc_color_out[8] ;
 wire \led_controller.led_effect_pulse.calc_color_out[9] ;
 wire \led_controller.led_effect_pulse.calc_color_valid ;
 wire \led_controller.led_effect_pulse.color_1.active ;
 wire \led_controller.led_effect_pulse.color_1.counter[0] ;
 wire \led_controller.led_effect_pulse.color_1.counter[1] ;
 wire \led_controller.led_effect_pulse.color_1.i_strb ;
 wire \led_controller.led_effect_pulse.color_index[0] ;
 wire \led_controller.led_effect_pulse.color_index[1] ;
 wire \led_controller.led_effect_pulse.current_led[0] ;
 wire \led_controller.led_effect_pulse.current_led[1] ;
 wire \led_controller.led_effect_pulse.current_led[2] ;
 wire \led_controller.led_effect_pulse.current_led[3] ;
 wire \led_controller.led_effect_pulse.current_led[4] ;
 wire \led_controller.led_effect_pulse.current_led[5] ;
 wire \led_controller.led_effect_pulse.current_led[6] ;
 wire \led_controller.led_effect_pulse.current_led[7] ;
 wire \led_controller.led_effect_pulse.fade_out ;
 wire \led_controller.led_effect_pulse.finished ;
 wire \led_controller.led_effect_pulse.state[0] ;
 wire \led_controller.led_effect_pulse.state[1] ;
 wire \led_controller.o_data ;
 wire \led_controller.o_spi_miso ;
 wire \led_controller.register_address[0] ;
 wire \led_controller.register_address[1] ;
 wire \led_controller.register_address[2] ;
 wire \led_controller.register_address[3] ;
 wire \led_controller.register_address[4] ;
 wire \led_controller.register_address[5] ;
 wire \led_controller.register_address[6] ;
 wire \led_controller.register_address[7] ;
 wire \led_controller.register_data[0] ;
 wire \led_controller.register_data[1] ;
 wire \led_controller.register_data[2] ;
 wire \led_controller.register_data[3] ;
 wire \led_controller.register_data[4] ;
 wire \led_controller.register_data[5] ;
 wire \led_controller.register_data[6] ;
 wire \led_controller.register_data[7] ;
 wire \led_controller.reset.reset1 ;
 wire \led_controller.rgbw.color[0] ;
 wire \led_controller.rgbw.color[10] ;
 wire \led_controller.rgbw.color[11] ;
 wire \led_controller.rgbw.color[12] ;
 wire \led_controller.rgbw.color[13] ;
 wire \led_controller.rgbw.color[14] ;
 wire \led_controller.rgbw.color[15] ;
 wire \led_controller.rgbw.color[16] ;
 wire \led_controller.rgbw.color[17] ;
 wire \led_controller.rgbw.color[18] ;
 wire \led_controller.rgbw.color[19] ;
 wire \led_controller.rgbw.color[1] ;
 wire \led_controller.rgbw.color[20] ;
 wire \led_controller.rgbw.color[21] ;
 wire \led_controller.rgbw.color[22] ;
 wire \led_controller.rgbw.color[23] ;
 wire \led_controller.rgbw.color[24] ;
 wire \led_controller.rgbw.color[25] ;
 wire \led_controller.rgbw.color[26] ;
 wire \led_controller.rgbw.color[27] ;
 wire \led_controller.rgbw.color[28] ;
 wire \led_controller.rgbw.color[29] ;
 wire \led_controller.rgbw.color[2] ;
 wire \led_controller.rgbw.color[30] ;
 wire \led_controller.rgbw.color[31] ;
 wire \led_controller.rgbw.color[3] ;
 wire \led_controller.rgbw.color[4] ;
 wire \led_controller.rgbw.color[5] ;
 wire \led_controller.rgbw.color[6] ;
 wire \led_controller.rgbw.color[7] ;
 wire \led_controller.rgbw.color[8] ;
 wire \led_controller.rgbw.color[9] ;
 wire \led_controller.rgbw.counter[0] ;
 wire \led_controller.rgbw.counter[1] ;
 wire \led_controller.rgbw.counter[2] ;
 wire \led_controller.rgbw.counter[3] ;
 wire \led_controller.rgbw.counter[4] ;
 wire \led_controller.rgbw.counter[5] ;
 wire \led_controller.rgbw.counter[6] ;
 wire \led_controller.rgbw.counter[7] ;
 wire \led_controller.rgbw.high_cycles[0] ;
 wire \led_controller.rgbw.high_cycles[1] ;
 wire \led_controller.rgbw.high_cycles[2] ;
 wire \led_controller.rgbw.low_cycles[0] ;
 wire \led_controller.rgbw.low_cycles[1] ;
 wire \led_controller.rgbw.low_cycles[2] ;
 wire \led_controller.rgbw.low_cycles[3] ;
 wire \led_controller.rgbw.low_cycles[4] ;
 wire \led_controller.rgbw.low_cycles[5] ;
 wire \led_controller.rgbw.low_cycles[6] ;
 wire \led_controller.rgbw.low_cycles[7] ;
 wire \led_controller.rgbw.low_cycles[8] ;
 wire \led_controller.rgbw.low_cycles[9] ;
 wire \led_controller.rgbw.pixel_counter[0] ;
 wire \led_controller.rgbw.pixel_counter[1] ;
 wire \led_controller.rgbw.pixel_counter[2] ;
 wire \led_controller.rgbw.pixel_counter[3] ;
 wire \led_controller.rgbw.pixel_counter[4] ;
 wire \led_controller.rgbw.pixel_counter[5] ;
 wire \led_controller.rgbw.state[0] ;
 wire \led_controller.rgbw.state[1] ;
 wire \led_controller.rgbw.state[2] ;
 wire \led_controller.spi_data[0] ;
 wire \led_controller.spi_data[1] ;
 wire \led_controller.spi_data[2] ;
 wire \led_controller.spi_data[3] ;
 wire \led_controller.spi_data[4] ;
 wire \led_controller.spi_data[5] ;
 wire \led_controller.spi_data[6] ;
 wire \led_controller.spi_data[7] ;
 wire \led_controller.spi_data_write[0] ;
 wire \led_controller.spi_data_write[1] ;
 wire \led_controller.spi_data_write[2] ;
 wire \led_controller.spi_data_write[3] ;
 wire \led_controller.spi_data_write[4] ;
 wire \led_controller.spi_data_write[5] ;
 wire \led_controller.spi_data_write[6] ;
 wire \led_controller.spi_data_write[7] ;
 wire \led_controller.spi_data_write_strb ;
 wire \led_controller.spi_slave.data_bits[0] ;
 wire \led_controller.spi_slave.data_bits[1] ;
 wire \led_controller.spi_slave.data_bits[2] ;
 wire \led_controller.spi_slave.data_bits[3] ;
 wire \led_controller.spi_slave.last_sck ;
 wire \led_controller.spi_slave.last_ss ;
 wire \led_controller.spi_slave.mosi ;
 wire \led_controller.spi_slave.o_tx_start_strb ;
 wire \led_controller.spi_slave.output_register[0] ;
 wire \led_controller.spi_slave.output_register[1] ;
 wire \led_controller.spi_slave.output_register[2] ;
 wire \led_controller.spi_slave.output_register[3] ;
 wire \led_controller.spi_slave.output_register[4] ;
 wire \led_controller.spi_slave.output_register[5] ;
 wire \led_controller.spi_slave.output_register[6] ;
 wire \led_controller.spi_slave.output_register[7] ;
 wire \led_controller.spi_slave.sck ;
 wire \led_controller.spi_slave.ss_n ;
 wire \led_controller.spi_slave.sync_mosi.data ;
 wire \led_controller.spi_slave.sync_sck.data ;
 wire \led_controller.spi_slave.sync_ss_n.data ;
 wire \led_controller.spi_state[0] ;
 wire \led_controller.spi_state[1] ;
 wire \led_controller.spi_state[2] ;
 wire \led_controller.timer_100hz.counter[0] ;
 wire \led_controller.timer_100hz.counter[10] ;
 wire \led_controller.timer_100hz.counter[11] ;
 wire \led_controller.timer_100hz.counter[12] ;
 wire \led_controller.timer_100hz.counter[13] ;
 wire \led_controller.timer_100hz.counter[14] ;
 wire \led_controller.timer_100hz.counter[15] ;
 wire \led_controller.timer_100hz.counter[16] ;
 wire \led_controller.timer_100hz.counter[17] ;
 wire \led_controller.timer_100hz.counter[18] ;
 wire \led_controller.timer_100hz.counter[19] ;
 wire \led_controller.timer_100hz.counter[1] ;
 wire \led_controller.timer_100hz.counter[20] ;
 wire \led_controller.timer_100hz.counter[21] ;
 wire \led_controller.timer_100hz.counter[22] ;
 wire \led_controller.timer_100hz.counter[23] ;
 wire \led_controller.timer_100hz.counter[24] ;
 wire \led_controller.timer_100hz.counter[25] ;
 wire \led_controller.timer_100hz.counter[26] ;
 wire \led_controller.timer_100hz.counter[27] ;
 wire \led_controller.timer_100hz.counter[28] ;
 wire \led_controller.timer_100hz.counter[29] ;
 wire \led_controller.timer_100hz.counter[2] ;
 wire \led_controller.timer_100hz.counter[30] ;
 wire \led_controller.timer_100hz.counter[31] ;
 wire \led_controller.timer_100hz.counter[3] ;
 wire \led_controller.timer_100hz.counter[4] ;
 wire \led_controller.timer_100hz.counter[5] ;
 wire \led_controller.timer_100hz.counter[6] ;
 wire \led_controller.timer_100hz.counter[7] ;
 wire \led_controller.timer_100hz.counter[8] ;
 wire \led_controller.timer_100hz.counter[9] ;
 wire \led_controller.timer_100hz.div_counter[0] ;
 wire \led_controller.timer_100hz.div_counter[1] ;
 wire \led_controller.timer_100hz.div_counter[2] ;
 wire \led_controller.timer_100hz.div_counter[3] ;
 wire \led_controller.timer_100hz.div_counter[4] ;
 wire \led_controller.timer_100hz.div_counter[5] ;
 wire \led_controller.timer_100hz.div_counter[6] ;
 wire \led_controller.timer_100hz.div_counter[7] ;
 wire \led_controller.timer_10hz.counter[0] ;
 wire \led_controller.timer_10hz.counter[1] ;
 wire \led_controller.timer_10hz.counter[2] ;
 wire \led_controller.timer_10hz.counter[3] ;
 wire \led_controller.timer_2hz.counter[0] ;
 wire \led_controller.timer_2hz.counter[1] ;
 wire \led_controller.timer_2hz.counter[2] ;
 wire \led_controller.timer_2hz.counter[3] ;
 wire \led_controller.timer_2hz.counter[4] ;
 wire \led_controller.timer_2hz.counter[5] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;

 sg13g2_inv_4 _4340_ (.A(net2042),
    .Y(_0740_));
 sg13g2_inv_4 _4341_ (.A(net2140),
    .Y(_0741_));
 sg13g2_inv_4 _4342_ (.A(net1948),
    .Y(_0742_));
 sg13g2_inv_4 _4343_ (.A(net2047),
    .Y(_0743_));
 sg13g2_inv_4 _4344_ (.A(net2000),
    .Y(_0744_));
 sg13g2_inv_4 _4345_ (.A(net2091),
    .Y(_0745_));
 sg13g2_inv_4 _4346_ (.A(net2124),
    .Y(_0746_));
 sg13g2_inv_4 _4347_ (.A(net2314),
    .Y(_0747_));
 sg13g2_inv_1 _4348_ (.Y(_0748_),
    .A(net2162));
 sg13g2_inv_1 _4349_ (.Y(_0749_),
    .A(\led_controller.cpu.i_num_leds[1] ));
 sg13g2_inv_2 _4350_ (.Y(_0750_),
    .A(net2128));
 sg13g2_inv_1 _4351_ (.Y(_0751_),
    .A(net2082));
 sg13g2_inv_1 _4352_ (.Y(_0752_),
    .A(\led_controller.register_address[1] ));
 sg13g2_inv_1 _4353_ (.Y(_0753_),
    .A(net1633));
 sg13g2_inv_1 _4354_ (.Y(_0754_),
    .A(net1952));
 sg13g2_inv_1 _4355_ (.Y(_0755_),
    .A(net1194));
 sg13g2_inv_2 _4356_ (.Y(_0756_),
    .A(\led_controller.cpu.i_bus_data_valid ));
 sg13g2_inv_1 _4357_ (.Y(_0757_),
    .A(net1170));
 sg13g2_inv_1 _4358_ (.Y(_0758_),
    .A(net1172));
 sg13g2_inv_1 _4359_ (.Y(_0759_),
    .A(net1175));
 sg13g2_inv_1 _4360_ (.Y(_0760_),
    .A(net1738));
 sg13g2_inv_1 _4361_ (.Y(_0761_),
    .A(net1921));
 sg13g2_inv_2 _4362_ (.Y(_0762_),
    .A(net1535));
 sg13g2_inv_1 _4363_ (.Y(_0763_),
    .A(net1414));
 sg13g2_inv_1 _4364_ (.Y(_0764_),
    .A(net1472));
 sg13g2_inv_2 _4365_ (.Y(_0765_),
    .A(net1619));
 sg13g2_inv_1 _4366_ (.Y(_0766_),
    .A(net1481));
 sg13g2_inv_1 _4367_ (.Y(_0767_),
    .A(net1457));
 sg13g2_inv_2 _4368_ (.Y(_0768_),
    .A(net1512));
 sg13g2_inv_2 _4369_ (.Y(_0769_),
    .A(net1549));
 sg13g2_inv_1 _4370_ (.Y(_0770_),
    .A(net1402));
 sg13g2_inv_1 _4371_ (.Y(_0771_),
    .A(net1391));
 sg13g2_inv_1 _4372_ (.Y(_0772_),
    .A(net1366));
 sg13g2_inv_1 _4373_ (.Y(_0773_),
    .A(net1375));
 sg13g2_inv_1 _4374_ (.Y(_0774_),
    .A(net1468));
 sg13g2_inv_1 _4375_ (.Y(_0775_),
    .A(net1587));
 sg13g2_inv_2 _4376_ (.Y(_0776_),
    .A(net1466));
 sg13g2_inv_2 _4377_ (.Y(_0777_),
    .A(net1487));
 sg13g2_inv_2 _4378_ (.Y(_0778_),
    .A(net1570));
 sg13g2_inv_2 _4379_ (.Y(_0779_),
    .A(net1643));
 sg13g2_inv_2 _4380_ (.Y(_0780_),
    .A(net1480));
 sg13g2_inv_2 _4381_ (.Y(_0781_),
    .A(net1604));
 sg13g2_inv_2 _4382_ (.Y(_0782_),
    .A(net1442));
 sg13g2_inv_2 _4383_ (.Y(_0783_),
    .A(net1447));
 sg13g2_inv_1 _4384_ (.Y(_0784_),
    .A(net1420));
 sg13g2_inv_2 _4385_ (.Y(_0785_),
    .A(net1511));
 sg13g2_inv_1 _4386_ (.Y(_0786_),
    .A(net1368));
 sg13g2_inv_1 _4387_ (.Y(_0787_),
    .A(net1432));
 sg13g2_inv_1 _4388_ (.Y(_0788_),
    .A(net1424));
 sg13g2_inv_1 _4389_ (.Y(_0789_),
    .A(net1422));
 sg13g2_inv_1 _4390_ (.Y(_0790_),
    .A(net1412));
 sg13g2_inv_1 _4391_ (.Y(_0791_),
    .A(net1396));
 sg13g2_inv_1 _4392_ (.Y(_0792_),
    .A(net1509));
 sg13g2_inv_2 _4393_ (.Y(_0793_),
    .A(net1426));
 sg13g2_inv_1 _4394_ (.Y(_0794_),
    .A(net1845));
 sg13g2_inv_1 _4395_ (.Y(_0795_),
    .A(net1653));
 sg13g2_inv_1 _4396_ (.Y(_0796_),
    .A(net2107));
 sg13g2_inv_1 _4397_ (.Y(_0797_),
    .A(net1265));
 sg13g2_inv_2 _4398_ (.Y(_0798_),
    .A(net1333));
 sg13g2_inv_1 _4399_ (.Y(_0799_),
    .A(net1734));
 sg13g2_inv_1 _4400_ (.Y(_0800_),
    .A(net1796));
 sg13g2_inv_1 _4401_ (.Y(_0801_),
    .A(net1628));
 sg13g2_inv_1 _4402_ (.Y(_0802_),
    .A(net1706));
 sg13g2_inv_1 _4403_ (.Y(_0803_),
    .A(net1850));
 sg13g2_inv_1 _4404_ (.Y(_0804_),
    .A(net2370));
 sg13g2_inv_1 _4405_ (.Y(_0805_),
    .A(\led_controller.flash.master.bit_counter[3] ));
 sg13g2_inv_1 _4406_ (.Y(_0806_),
    .A(net1389));
 sg13g2_inv_1 _4407_ (.Y(_0807_),
    .A(net1321));
 sg13g2_inv_1 _4408_ (.Y(_0808_),
    .A(net1356));
 sg13g2_inv_1 _4409_ (.Y(_0809_),
    .A(net1329));
 sg13g2_inv_1 _4410_ (.Y(_0810_),
    .A(net1325));
 sg13g2_inv_1 _4411_ (.Y(_0811_),
    .A(net1378));
 sg13g2_inv_1 _4412_ (.Y(_0812_),
    .A(net1602));
 sg13g2_inv_1 _4413_ (.Y(_0813_),
    .A(net1384));
 sg13g2_inv_1 _4414_ (.Y(_0814_),
    .A(net1343));
 sg13g2_inv_1 _4415_ (.Y(_0815_),
    .A(net1370));
 sg13g2_inv_1 _4416_ (.Y(_0816_),
    .A(net1398));
 sg13g2_inv_1 _4417_ (.Y(_0817_),
    .A(net1382));
 sg13g2_inv_1 _4418_ (.Y(_0818_),
    .A(net1430));
 sg13g2_inv_1 _4419_ (.Y(_0819_),
    .A(net1492));
 sg13g2_inv_1 _4420_ (.Y(_0820_),
    .A(net1474));
 sg13g2_inv_1 _4421_ (.Y(_0821_),
    .A(net1400));
 sg13g2_inv_1 _4422_ (.Y(_0822_),
    .A(net1437));
 sg13g2_inv_1 _4423_ (.Y(_0823_),
    .A(net1836));
 sg13g2_inv_1 _4424_ (.Y(_0824_),
    .A(net1434));
 sg13g2_inv_1 _4425_ (.Y(_0825_),
    .A(net1445));
 sg13g2_inv_1 _4426_ (.Y(_0826_),
    .A(net1485));
 sg13g2_inv_1 _4427_ (.Y(_0827_),
    .A(net1449));
 sg13g2_inv_1 _4428_ (.Y(_0828_),
    .A(net1476));
 sg13g2_inv_1 _4429_ (.Y(_0829_),
    .A(net1517));
 sg13g2_inv_1 _4430_ (.Y(_0830_),
    .A(net1461));
 sg13g2_inv_1 _4431_ (.Y(_0831_),
    .A(net1503));
 sg13g2_inv_1 _4432_ (.Y(_0832_),
    .A(net1505));
 sg13g2_inv_1 _4433_ (.Y(_0833_),
    .A(net1834));
 sg13g2_inv_1 _4434_ (.Y(_0834_),
    .A(net1553));
 sg13g2_inv_1 _4435_ (.Y(_0835_),
    .A(net1496));
 sg13g2_inv_1 _4436_ (.Y(_0836_),
    .A(net1561));
 sg13g2_inv_1 _4437_ (.Y(_0837_),
    .A(\led_controller.cpu.fetch_pc[4] ));
 sg13g2_inv_1 _4438_ (.Y(_0838_),
    .A(net1451));
 sg13g2_inv_1 _4439_ (.Y(_0839_),
    .A(net1483));
 sg13g2_inv_1 _4440_ (.Y(_0840_),
    .A(net1345));
 sg13g2_inv_1 _4441_ (.Y(_0841_),
    .A(net1359));
 sg13g2_inv_1 _4442_ (.Y(_0842_),
    .A(net1339));
 sg13g2_inv_1 _4443_ (.Y(_0843_),
    .A(net1807));
 sg13g2_inv_1 _4444_ (.Y(_0844_),
    .A(net1941));
 sg13g2_inv_2 _4445_ (.Y(_0845_),
    .A(net1840));
 sg13g2_inv_2 _4446_ (.Y(_0846_),
    .A(net2055));
 sg13g2_inv_2 _4447_ (.Y(_0847_),
    .A(net2192));
 sg13g2_inv_1 _4448_ (.Y(_0848_),
    .A(net1507));
 sg13g2_inv_1 _4449_ (.Y(_0849_),
    .A(net1443));
 sg13g2_inv_2 _4450_ (.Y(_0850_),
    .A(net1597));
 sg13g2_inv_2 _4451_ (.Y(_0851_),
    .A(net1624));
 sg13g2_inv_2 _4452_ (.Y(_0852_),
    .A(net2270));
 sg13g2_inv_2 _4453_ (.Y(_0853_),
    .A(net2292));
 sg13g2_inv_1 _4454_ (.Y(_0854_),
    .A(net2266));
 sg13g2_inv_2 _4455_ (.Y(_0855_),
    .A(net2304));
 sg13g2_inv_1 _4456_ (.Y(_0856_),
    .A(net2315));
 sg13g2_inv_1 _4457_ (.Y(_0857_),
    .A(net1531));
 sg13g2_inv_1 _4458_ (.Y(_0858_),
    .A(\led_controller.cpu.status_zero ));
 sg13g2_inv_2 _4459_ (.Y(_0859_),
    .A(net2318));
 sg13g2_inv_4 _4460_ (.A(net2247),
    .Y(_0860_));
 sg13g2_inv_1 _4461_ (.Y(_0861_),
    .A(net2210));
 sg13g2_inv_2 _4462_ (.Y(_0862_),
    .A(\led_controller.cpu.register_x[6] ));
 sg13g2_inv_1 _4463_ (.Y(_0863_),
    .A(net1182));
 sg13g2_inv_2 _4464_ (.Y(_0864_),
    .A(\led_controller.cpu.register_x[3] ));
 sg13g2_inv_1 _4465_ (.Y(_0865_),
    .A(net1183));
 sg13g2_inv_1 _4466_ (.Y(_0866_),
    .A(\led_controller.cpu.pc[11] ));
 sg13g2_inv_1 _4467_ (.Y(_0867_),
    .A(\led_controller.cpu.pc[8] ));
 sg13g2_inv_1 _4468_ (.Y(_0868_),
    .A(\led_controller.cpu.pc[6] ));
 sg13g2_inv_2 _4469_ (.Y(_0869_),
    .A(\led_controller.cpu.pc[4] ));
 sg13g2_inv_1 _4470_ (.Y(_0870_),
    .A(net1635));
 sg13g2_inv_1 _4471_ (.Y(_0871_),
    .A(net1435));
 sg13g2_inv_1 _4472_ (.Y(_0872_),
    .A(net1478));
 sg13g2_inv_1 _4473_ (.Y(_0873_),
    .A(\led_controller.cpu.o_led_strb ));
 sg13g2_inv_1 _4474_ (.Y(_0874_),
    .A(net1646));
 sg13g2_inv_1 _4475_ (.Y(_0875_),
    .A(net1732));
 sg13g2_inv_1 _4476_ (.Y(_0876_),
    .A(net2213));
 sg13g2_inv_1 _4477_ (.Y(_0877_),
    .A(net2324));
 sg13g2_inv_1 _4478_ (.Y(_0878_),
    .A(net2104));
 sg13g2_inv_1 _4479_ (.Y(_0879_),
    .A(net2063));
 sg13g2_inv_1 _4480_ (.Y(_0880_),
    .A(net2328));
 sg13g2_inv_1 _4481_ (.Y(_0881_),
    .A(\led_controller.timer_2hz.counter[1] ));
 sg13g2_inv_1 _4482_ (.Y(_0882_),
    .A(net2283));
 sg13g2_inv_1 _4483_ (.Y(_0883_),
    .A(net1191));
 sg13g2_inv_1 _4484_ (.Y(_0884_),
    .A(net1153));
 sg13g2_inv_2 _4485_ (.Y(_0885_),
    .A(net1165));
 sg13g2_inv_1 _4486_ (.Y(_0886_),
    .A(\led_controller.flash.cs_delay_counter[1] ));
 sg13g2_inv_1 _4487_ (.Y(_0887_),
    .A(net1993));
 sg13g2_inv_1 _4488_ (.Y(_0888_),
    .A(net1665));
 sg13g2_inv_1 _4489_ (.Y(_0889_),
    .A(net2077));
 sg13g2_inv_1 _4490_ (.Y(_0890_),
    .A(\led_controller.led_effect_chase.finished ));
 sg13g2_inv_2 _4491_ (.Y(uio_oe[0]),
    .A(net3));
 sg13g2_inv_1 _4492_ (.Y(_0891_),
    .A(net1903));
 sg13g2_inv_1 _4493_ (.Y(_0892_),
    .A(net783));
 sg13g2_inv_1 _4494_ (.Y(_0893_),
    .A(\led_controller.spi_slave.output_register[7] ));
 sg13g2_inv_1 _4495_ (.Y(_0894_),
    .A(net1196));
 sg13g2_inv_4 _4496_ (.A(net1195),
    .Y(_0895_));
 sg13g2_inv_1 _4497_ (.Y(_0896_),
    .A(\led_controller.cpu.scratch_memory[4][2] ));
 sg13g2_inv_1 _4498_ (.Y(_0897_),
    .A(\led_controller.cpu.scratch_memory[12][4] ));
 sg13g2_inv_1 _4499_ (.Y(_0898_),
    .A(\led_controller.cpu.scratch_memory[12][5] ));
 sg13g2_inv_1 _4500_ (.Y(_0899_),
    .A(\led_controller.cpu.scratch_memory[12][6] ));
 sg13g2_inv_1 _4501_ (.Y(_0900_),
    .A(\led_controller.cpu.scratch_memory[4][7] ));
 sg13g2_inv_1 _4502_ (.Y(_0901_),
    .A(\led_controller.cpu.scratch_memory[14][7] ));
 sg13g2_inv_2 _4503_ (.Y(_0902_),
    .A(net1164));
 sg13g2_nor4_1 _4504_ (.A(net2295),
    .B(\led_controller.cpu_reset_counter[1] ),
    .C(\led_controller.cpu_reset_counter[3] ),
    .D(\led_controller.cpu_reset_counter[2] ),
    .Y(_0903_));
 sg13g2_and2_1 _4505_ (.A(net1144),
    .B(_0903_),
    .X(_0904_));
 sg13g2_nand2_1 _4506_ (.Y(_0905_),
    .A(net1144),
    .B(_0903_));
 sg13g2_nand2_1 _4507_ (.Y(_0906_),
    .A(net2315),
    .B(net1056));
 sg13g2_nor2_2 _4508_ (.A(net2355),
    .B(_0906_),
    .Y(_0907_));
 sg13g2_and2_1 _4509_ (.A(net2355),
    .B(net1057),
    .X(_0908_));
 sg13g2_a22oi_1 _4510_ (.Y(_0909_),
    .B1(_0908_),
    .B2(net1192),
    .A2(_0907_),
    .A1(net1193));
 sg13g2_inv_1 _4511_ (.Y(_0005_),
    .A(_0909_));
 sg13g2_nor2_2 _4512_ (.A(net2059),
    .B(net2118),
    .Y(_0910_));
 sg13g2_nand2_1 _4513_ (.Y(_0911_),
    .A(\led_controller.effect[1] ),
    .B(_0910_));
 sg13g2_nor2_1 _4514_ (.A(\led_controller.effect[0] ),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_nand3_1 _4515_ (.B(_0748_),
    .C(_0910_),
    .A(\led_controller.effect[1] ),
    .Y(_0913_));
 sg13g2_a21oi_2 _4516_ (.B1(net1121),
    .Y(_0914_),
    .A2(_0913_),
    .A1(\led_controller.led_effect_pulse.finished ));
 sg13g2_a21o_2 _4517_ (.A2(_0913_),
    .A1(net2238),
    .B1(net1121),
    .X(_0915_));
 sg13g2_nor2_2 _4518_ (.A(net1876),
    .B(net1191),
    .Y(_0916_));
 sg13g2_or2_1 _4519_ (.X(_0917_),
    .B(net1191),
    .A(\led_controller.rgbw.state[0] ));
 sg13g2_nor3_2 _4520_ (.A(\led_controller.led_effect_pulse.finished ),
    .B(_0794_),
    .C(net1098),
    .Y(_0918_));
 sg13g2_nand2_1 _4521_ (.Y(_0919_),
    .A(net994),
    .B(_0918_));
 sg13g2_nand3_1 _4522_ (.B(net994),
    .C(_0918_),
    .A(net1380),
    .Y(_0920_));
 sg13g2_o21ai_1 _4523_ (.B1(net1708),
    .Y(_0921_),
    .A1(_0887_),
    .A2(_0913_));
 sg13g2_nand3_1 _4524_ (.B(_0920_),
    .C(net1709),
    .A(net985),
    .Y(_0011_));
 sg13g2_nand2_1 _4525_ (.Y(_0922_),
    .A(net1380),
    .B(_0919_));
 sg13g2_nand3_1 _4526_ (.B(\led_controller.led_effect_pulse.calc_color_valid ),
    .C(net994),
    .A(\led_controller.led_effect_pulse.state[0] ),
    .Y(_0923_));
 sg13g2_a21oi_1 _4527_ (.A1(_0922_),
    .A2(_0923_),
    .Y(_0012_),
    .B1(_0915_));
 sg13g2_nor2_1 _4528_ (.A(net1704),
    .B(\led_controller.rgbw.low_cycles[0] ),
    .Y(_0924_));
 sg13g2_nor3_1 _4529_ (.A(net2112),
    .B(net1704),
    .C(\led_controller.rgbw.low_cycles[0] ),
    .Y(_0925_));
 sg13g2_nand2b_1 _4530_ (.Y(_0926_),
    .B(_0925_),
    .A_N(net2028));
 sg13g2_nand2b_2 _4531_ (.Y(_0927_),
    .B(_0874_),
    .A_N(_0926_));
 sg13g2_inv_1 _4532_ (.Y(_0928_),
    .A(_0927_));
 sg13g2_nor3_2 _4533_ (.A(net2096),
    .B(\led_controller.rgbw.low_cycles[5] ),
    .C(_0927_),
    .Y(_0929_));
 sg13g2_nand2b_2 _4534_ (.Y(_0930_),
    .B(_0929_),
    .A_N(\led_controller.rgbw.low_cycles[7] ));
 sg13g2_nor2_1 _4535_ (.A(net2099),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_nor3_2 _4536_ (.A(net1890),
    .B(net2099),
    .C(_0930_),
    .Y(_0932_));
 sg13g2_nand2b_2 _4537_ (.Y(_0933_),
    .B(_0931_),
    .A_N(net1890));
 sg13g2_a21o_1 _4538_ (.A2(_0933_),
    .A1(net1876),
    .B1(net1117),
    .X(_0013_));
 sg13g2_nand3_1 _4539_ (.B(\led_controller.effect[0] ),
    .C(_0910_),
    .A(\led_controller.effect[1] ),
    .Y(_0934_));
 sg13g2_nor2_1 _4540_ (.A(_0873_),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_a221oi_1 _4541_ (.B2(\led_controller.effect_pulse_led_strb ),
    .C1(_0935_),
    .B1(net993),
    .A1(\led_controller.effect_chase_led_strb ),
    .Y(_0936_),
    .A2(_0911_));
 sg13g2_nand2b_1 _4542_ (.Y(_0937_),
    .B(net1098),
    .A_N(_0936_));
 sg13g2_inv_1 _4543_ (.Y(_0938_),
    .A(_0937_));
 sg13g2_a22oi_1 _4544_ (.Y(_0939_),
    .B1(_0937_),
    .B2(net2373),
    .A2(_0932_),
    .A1(net1876));
 sg13g2_or3_1 _4545_ (.A(\led_controller.clock_divider[2] ),
    .B(\led_controller.clock_divider[1] ),
    .C(\led_controller.clock_divider[0] ),
    .X(_0940_));
 sg13g2_or2_1 _4546_ (.X(_0941_),
    .B(_0940_),
    .A(\led_controller.clock_divider[3] ));
 sg13g2_nor3_2 _4547_ (.A(\led_controller.clock_divider[5] ),
    .B(\led_controller.clock_divider[4] ),
    .C(_0941_),
    .Y(_0942_));
 sg13g2_nor2b_1 _4548_ (.A(\led_controller.clock_divider[6] ),
    .B_N(_0942_),
    .Y(_0943_));
 sg13g2_xnor2_1 _4549_ (.Y(_0944_),
    .A(\led_controller.clock_divider[6] ),
    .B(_0942_));
 sg13g2_nand2b_2 _4550_ (.Y(_0945_),
    .B(\led_controller.clock_divider[7] ),
    .A_N(_0943_));
 sg13g2_xnor2_1 _4551_ (.Y(_0946_),
    .A(\led_controller.rgbw.counter[7] ),
    .B(_0945_));
 sg13g2_nor2b_2 _4552_ (.A(net2111),
    .B_N(_0943_),
    .Y(_0947_));
 sg13g2_xor2_1 _4553_ (.B(_0940_),
    .A(\led_controller.clock_divider[3] ),
    .X(_0948_));
 sg13g2_xnor2_1 _4554_ (.Y(_0949_),
    .A(\led_controller.rgbw.counter[3] ),
    .B(_0948_));
 sg13g2_xor2_1 _4555_ (.B(\led_controller.clock_divider[0] ),
    .A(\led_controller.clock_divider[1] ),
    .X(_0950_));
 sg13g2_xnor2_1 _4556_ (.Y(_0951_),
    .A(\led_controller.clock_divider[0] ),
    .B(\led_controller.rgbw.counter[0] ));
 sg13g2_xnor2_1 _4557_ (.Y(_0952_),
    .A(\led_controller.rgbw.counter[1] ),
    .B(_0950_));
 sg13g2_o21ai_1 _4558_ (.B1(\led_controller.clock_divider[2] ),
    .Y(_0953_),
    .A1(\led_controller.clock_divider[1] ),
    .A2(\led_controller.clock_divider[0] ));
 sg13g2_and2_1 _4559_ (.A(_0940_),
    .B(_0953_),
    .X(_0954_));
 sg13g2_xnor2_1 _4560_ (.Y(_0955_),
    .A(\led_controller.rgbw.counter[2] ),
    .B(_0954_));
 sg13g2_nor4_1 _4561_ (.A(_0949_),
    .B(_0951_),
    .C(_0952_),
    .D(_0955_),
    .Y(_0956_));
 sg13g2_o21ai_1 _4562_ (.B1(\led_controller.clock_divider[5] ),
    .Y(_0957_),
    .A1(\led_controller.clock_divider[4] ),
    .A2(_0941_));
 sg13g2_nor2b_2 _4563_ (.A(_0942_),
    .B_N(_0957_),
    .Y(_0958_));
 sg13g2_xor2_1 _4564_ (.B(_0941_),
    .A(\led_controller.clock_divider[4] ),
    .X(_0959_));
 sg13g2_xor2_1 _4565_ (.B(_0959_),
    .A(\led_controller.rgbw.counter[4] ),
    .X(_0960_));
 sg13g2_xor2_1 _4566_ (.B(_0944_),
    .A(\led_controller.rgbw.counter[6] ),
    .X(_0961_));
 sg13g2_nand3_1 _4567_ (.B(_0960_),
    .C(_0961_),
    .A(_0956_),
    .Y(_0962_));
 sg13g2_xnor2_1 _4568_ (.Y(_0963_),
    .A(\led_controller.rgbw.counter[5] ),
    .B(_0958_));
 sg13g2_nor4_2 _4569_ (.A(_0946_),
    .B(_0947_),
    .C(_0962_),
    .Y(_0964_),
    .D(_0963_));
 sg13g2_nor2_2 _4570_ (.A(net1189),
    .B(net1190),
    .Y(_0965_));
 sg13g2_nor3_1 _4571_ (.A(\led_controller.rgbw.pixel_counter[2] ),
    .B(net1189),
    .C(net1190),
    .Y(_0966_));
 sg13g2_nor2b_2 _4572_ (.A(net1978),
    .B_N(_0966_),
    .Y(_0967_));
 sg13g2_and3_2 _4573_ (.X(_0968_),
    .A(_0875_),
    .B(_0876_),
    .C(_0967_));
 sg13g2_nand3_1 _4574_ (.B(_0964_),
    .C(_0968_),
    .A(_0932_),
    .Y(_0969_));
 sg13g2_o21ai_1 _4575_ (.B1(_0939_),
    .Y(_0970_),
    .A1(_0883_),
    .A2(_0969_));
 sg13g2_and2_1 _4576_ (.A(net1152),
    .B(_0970_),
    .X(_0014_));
 sg13g2_nand2_1 _4577_ (.Y(_0971_),
    .A(\led_controller.rgbw.state[1] ),
    .B(_0938_));
 sg13g2_nand2_1 _4578_ (.Y(_0972_),
    .A(net1191),
    .B(_0969_));
 sg13g2_a21oi_1 _4579_ (.A1(net856),
    .A2(_0972_),
    .Y(_0015_),
    .B1(net1117));
 sg13g2_nor4_2 _4580_ (.A(net1966),
    .B(net1494),
    .C(net1887),
    .Y(_0973_),
    .D(_0888_));
 sg13g2_a21oi_1 _4581_ (.A1(net1825),
    .A2(\led_controller.spi_state[1] ),
    .Y(_0974_),
    .B1(\led_controller.spi_state[0] ));
 sg13g2_o21ai_1 _4582_ (.B1(net1150),
    .Y(_0016_),
    .A1(_0973_),
    .A2(net1826));
 sg13g2_nand2_2 _4583_ (.Y(_0975_),
    .A(net2317),
    .B(_0973_));
 sg13g2_nand3_1 _4584_ (.B(net2317),
    .C(_0973_),
    .A(net1916),
    .Y(_0976_));
 sg13g2_nand2b_1 _4585_ (.Y(_0977_),
    .B(net2014),
    .A_N(net1825));
 sg13g2_o21ai_1 _4586_ (.B1(_0976_),
    .Y(_0978_),
    .A1(_0973_),
    .A2(_0977_));
 sg13g2_o21ai_1 _4587_ (.B1(net1145),
    .Y(_0979_),
    .A1(net1194),
    .A2(_0978_));
 sg13g2_inv_1 _4588_ (.Y(_0017_),
    .A(_0979_));
 sg13g2_nand2_2 _4589_ (.Y(_0980_),
    .A(net2014),
    .B(_0973_));
 sg13g2_o21ai_1 _4590_ (.B1(net984),
    .Y(_0981_),
    .A1(net1916),
    .A2(_0975_));
 sg13g2_and2_1 _4591_ (.A(net1145),
    .B(_0981_),
    .X(_0018_));
 sg13g2_or2_1 _4592_ (.X(_0982_),
    .B(net764),
    .A(net2343));
 sg13g2_or2_1 _4593_ (.X(_0983_),
    .B(_0982_),
    .A(net1555));
 sg13g2_nor2_1 _4594_ (.A(\led_controller.flash.cs_delay_counter[3] ),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_nor3_1 _4595_ (.A(\led_controller.flash.cs_delay_counter[3] ),
    .B(\led_controller.flash.cs_delay_counter[4] ),
    .C(_0983_),
    .Y(_0985_));
 sg13g2_nand2b_1 _4596_ (.Y(_0986_),
    .B(_0985_),
    .A_N(net1718));
 sg13g2_or2_1 _4597_ (.X(_0987_),
    .B(_0986_),
    .A(net1605));
 sg13g2_nor2_1 _4598_ (.A(\led_controller.flash.cs_delay_counter[7] ),
    .B(_0987_),
    .Y(_0988_));
 sg13g2_nor3_2 _4599_ (.A(net1608),
    .B(net1566),
    .C(_0987_),
    .Y(_0989_));
 sg13g2_nor2_1 _4600_ (.A(_0889_),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_nor4_2 _4601_ (.A(net1936),
    .B(net1192),
    .C(net1500),
    .Y(_0991_),
    .D(net1528));
 sg13g2_nor2_1 _4602_ (.A(net1353),
    .B(net1041),
    .Y(_0992_));
 sg13g2_o21ai_1 _4603_ (.B1(_0992_),
    .Y(_0993_),
    .A1(\led_controller.flash.master.o_rx_data_valid ),
    .A2(_0991_));
 sg13g2_o21ai_1 _4604_ (.B1(_0906_),
    .Y(_0994_),
    .A1(_0990_),
    .A2(_0993_));
 sg13g2_nand3_1 _4605_ (.B(\led_controller.cpu.o_bus_addr_valid ),
    .C(_0989_),
    .A(\led_controller.flash.o_cs_n ),
    .Y(_0995_));
 sg13g2_nand3_1 _4606_ (.B(net1056),
    .C(_0995_),
    .A(net1575),
    .Y(_0996_));
 sg13g2_nor2_1 _4607_ (.A(net1176),
    .B(net1942),
    .Y(_0997_));
 sg13g2_nand2_1 _4608_ (.Y(_0004_),
    .A(_0994_),
    .B(net1576));
 sg13g2_nand2_1 _4609_ (.Y(_0998_),
    .A(net1500),
    .B(_0907_));
 sg13g2_nand4_1 _4610_ (.B(\led_controller.flash.state[4] ),
    .C(net1056),
    .A(\led_controller.flash.i_addr_width_24 ),
    .Y(_0999_),
    .D(_0989_));
 sg13g2_nand2_1 _4611_ (.Y(_0006_),
    .A(net1501),
    .B(_0999_));
 sg13g2_a22oi_1 _4612_ (.Y(_1000_),
    .B1(_0908_),
    .B2(net1500),
    .A2(_0907_),
    .A1(net1192));
 sg13g2_nand3b_1 _4613_ (.B(net1056),
    .C(_0989_),
    .Y(_1001_),
    .A_N(\led_controller.flash.i_addr_width_24 ));
 sg13g2_o21ai_1 _4614_ (.B1(_1000_),
    .Y(_0010_),
    .A1(_0889_),
    .A2(_1001_));
 sg13g2_a22oi_1 _4615_ (.Y(_1002_),
    .B1(_0908_),
    .B2(net1936),
    .A2(_0907_),
    .A1(net1528));
 sg13g2_inv_1 _4616_ (.Y(_0009_),
    .A(net1937));
 sg13g2_nand2b_1 _4617_ (.Y(_1003_),
    .B(_0990_),
    .A_N(_0906_));
 sg13g2_nand4_1 _4618_ (.B(net2361),
    .C(net1575),
    .A(net1942),
    .Y(_1004_),
    .D(_0989_));
 sg13g2_o21ai_1 _4619_ (.B1(_1003_),
    .Y(_0008_),
    .A1(net1041),
    .A2(net854));
 sg13g2_nand2_1 _4620_ (.Y(_1005_),
    .A(net1528),
    .B(_0908_));
 sg13g2_nand2_1 _4621_ (.Y(_1006_),
    .A(\led_controller.cpu.o_bus_addr_valid ),
    .B(net1353));
 sg13g2_o21ai_1 _4622_ (.B1(net1529),
    .Y(_0007_),
    .A1(net1040),
    .A2(_1006_));
 sg13g2_nor4_1 _4623_ (.A(net1823),
    .B(net1525),
    .C(net1899),
    .D(net1563),
    .Y(_1007_));
 sg13g2_nor4_1 _4624_ (.A(net2161),
    .B(net1926),
    .C(net1519),
    .D(net2167),
    .Y(_1008_));
 sg13g2_and2_1 _4625_ (.A(_1007_),
    .B(_1008_),
    .X(_1009_));
 sg13g2_and2_1 _4626_ (.A(_0991_),
    .B(_1006_),
    .X(_1010_));
 sg13g2_a21oi_1 _4627_ (.A1(_1009_),
    .A2(_1010_),
    .Y(\led_controller.flash.master.o_sck ),
    .B1(_0798_));
 sg13g2_nand2_1 _4628_ (.Y(_1011_),
    .A(net1982),
    .B(net1961));
 sg13g2_nor3_1 _4629_ (.A(net1558),
    .B(net1697),
    .C(_1011_),
    .Y(_1012_));
 sg13g2_nor2_2 _4630_ (.A(net1708),
    .B(_0913_),
    .Y(_1013_));
 sg13g2_and2_1 _4631_ (.A(_1012_),
    .B(_1013_),
    .X(_1014_));
 sg13g2_and2_1 _4632_ (.A(net2238),
    .B(_1014_),
    .X(_1015_));
 sg13g2_nand2_2 _4633_ (.Y(_1016_),
    .A(net2238),
    .B(_1014_));
 sg13g2_nor2_2 _4634_ (.A(net1174),
    .B(net1175),
    .Y(_1017_));
 sg13g2_nand3_1 _4635_ (.B(_0758_),
    .C(_1017_),
    .A(_0757_),
    .Y(_1018_));
 sg13g2_nor2_1 _4636_ (.A(net951),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_nor3_1 _4637_ (.A(net1168),
    .B(net951),
    .C(_1018_),
    .Y(_1020_));
 sg13g2_o21ai_1 _4638_ (.B1(net986),
    .Y(_1021_),
    .A1(net2283),
    .A2(_1019_));
 sg13g2_nor2_1 _4639_ (.A(_1020_),
    .B(_1021_),
    .Y(_0019_));
 sg13g2_xor2_1 _4640_ (.B(\led_controller.cpu.pc[1] ),
    .A(\led_controller.cpu.fetch_pc[1] ),
    .X(_1022_));
 sg13g2_xnor2_1 _4641_ (.Y(_1023_),
    .A(\led_controller.cpu.fetch_pc[14] ),
    .B(\led_controller.cpu.pc[14] ));
 sg13g2_xnor2_1 _4642_ (.Y(_1024_),
    .A(\led_controller.cpu.fetch_pc[15] ),
    .B(\led_controller.cpu.pc[15] ));
 sg13g2_xnor2_1 _4643_ (.Y(_1025_),
    .A(\led_controller.cpu.fetch_pc[11] ),
    .B(\led_controller.cpu.pc[11] ));
 sg13g2_xnor2_1 _4644_ (.Y(_1026_),
    .A(\led_controller.cpu.fetch_pc[0] ),
    .B(\led_controller.cpu.pc[0] ));
 sg13g2_xor2_1 _4645_ (.B(\led_controller.cpu.pc[13] ),
    .A(\led_controller.cpu.fetch_pc[13] ),
    .X(_1027_));
 sg13g2_xor2_1 _4646_ (.B(\led_controller.cpu.pc[2] ),
    .A(\led_controller.cpu.fetch_pc[2] ),
    .X(_1028_));
 sg13g2_xnor2_1 _4647_ (.Y(_1029_),
    .A(\led_controller.cpu.fetch_pc[10] ),
    .B(\led_controller.cpu.pc[10] ));
 sg13g2_xor2_1 _4648_ (.B(\led_controller.cpu.pc[9] ),
    .A(\led_controller.cpu.fetch_pc[9] ),
    .X(_1030_));
 sg13g2_xor2_1 _4649_ (.B(\led_controller.cpu.pc[8] ),
    .A(\led_controller.cpu.fetch_pc[8] ),
    .X(_1031_));
 sg13g2_xor2_1 _4650_ (.B(\led_controller.cpu.pc[6] ),
    .A(\led_controller.cpu.fetch_pc[6] ),
    .X(_1032_));
 sg13g2_xor2_1 _4651_ (.B(\led_controller.cpu.pc[5] ),
    .A(\led_controller.cpu.fetch_pc[5] ),
    .X(_1033_));
 sg13g2_nor3_1 _4652_ (.A(_1027_),
    .B(_1030_),
    .C(_1033_),
    .Y(_1034_));
 sg13g2_xor2_1 _4653_ (.B(\led_controller.cpu.pc[7] ),
    .A(\led_controller.cpu.fetch_pc[7] ),
    .X(_1035_));
 sg13g2_nor3_1 _4654_ (.A(_1022_),
    .B(_1028_),
    .C(_1035_),
    .Y(_1036_));
 sg13g2_xnor2_1 _4655_ (.Y(_1037_),
    .A(\led_controller.cpu.fetch_pc[12] ),
    .B(\led_controller.cpu.pc[12] ));
 sg13g2_nand4_1 _4656_ (.B(_1024_),
    .C(_1025_),
    .A(_1023_),
    .Y(_1038_),
    .D(_1037_));
 sg13g2_xnor2_1 _4657_ (.Y(_1039_),
    .A(\led_controller.cpu.fetch_pc[3] ),
    .B(\led_controller.cpu.pc[3] ));
 sg13g2_xnor2_1 _4658_ (.Y(_1040_),
    .A(\led_controller.cpu.fetch_pc[4] ),
    .B(\led_controller.cpu.pc[4] ));
 sg13g2_nand4_1 _4659_ (.B(_1029_),
    .C(_1039_),
    .A(_1026_),
    .Y(_1041_),
    .D(_1040_));
 sg13g2_nor4_1 _4660_ (.A(_1031_),
    .B(_1032_),
    .C(_1038_),
    .D(_1041_),
    .Y(_1042_));
 sg13g2_nand3_1 _4661_ (.B(_1036_),
    .C(_1042_),
    .A(_1034_),
    .Y(_1043_));
 sg13g2_nor2_2 _4662_ (.A(_0823_),
    .B(_1043_),
    .Y(_1044_));
 sg13g2_or2_1 _4663_ (.X(_1045_),
    .B(_1043_),
    .A(_0823_));
 sg13g2_o21ai_1 _4664_ (.B1(net1059),
    .Y(_1046_),
    .A1(net1954),
    .A2(net945));
 sg13g2_a21oi_1 _4665_ (.A1(_0855_),
    .A2(net945),
    .Y(_0020_),
    .B1(_1046_));
 sg13g2_o21ai_1 _4666_ (.B1(net1059),
    .Y(_1047_),
    .A1(net1756),
    .A2(net945));
 sg13g2_a21oi_1 _4667_ (.A1(_0854_),
    .A2(net947),
    .Y(_0021_),
    .B1(_1047_));
 sg13g2_o21ai_1 _4668_ (.B1(net1059),
    .Y(_1048_),
    .A1(net1969),
    .A2(net946));
 sg13g2_a21oi_1 _4669_ (.A1(_0853_),
    .A2(net946),
    .Y(_0022_),
    .B1(_1048_));
 sg13g2_o21ai_1 _4670_ (.B1(net1059),
    .Y(_1049_),
    .A1(net1767),
    .A2(net945));
 sg13g2_a21oi_1 _4671_ (.A1(_0852_),
    .A2(net946),
    .Y(_0023_),
    .B1(_1049_));
 sg13g2_nor2_2 _4672_ (.A(_0854_),
    .B(net2304),
    .Y(_1050_));
 sg13g2_nand2_2 _4673_ (.Y(_1051_),
    .A(\led_controller.cpu.current_instruction[1] ),
    .B(_0855_));
 sg13g2_nor2_2 _4674_ (.A(\led_controller.cpu.current_instruction[1] ),
    .B(\led_controller.cpu.current_instruction[0] ),
    .Y(_1052_));
 sg13g2_or2_1 _4675_ (.X(_1053_),
    .B(\led_controller.cpu.current_instruction[0] ),
    .A(\led_controller.cpu.current_instruction[1] ));
 sg13g2_nor2_1 _4676_ (.A(\led_controller.cpu.current_instruction[3] ),
    .B(net2389),
    .Y(_1054_));
 sg13g2_or3_1 _4677_ (.A(\led_controller.cpu.current_instruction[4] ),
    .B(\led_controller.cpu.current_instruction[3] ),
    .C(\led_controller.cpu.current_instruction[2] ),
    .X(_1055_));
 sg13g2_o21ai_1 _4678_ (.B1(\led_controller.cpu.current_instruction[5] ),
    .Y(_1056_),
    .A1(_1053_),
    .A2(_1055_));
 sg13g2_nor2_1 _4679_ (.A(net1507),
    .B(net1443),
    .Y(_1057_));
 sg13g2_nand2_1 _4680_ (.Y(_1058_),
    .A(_0850_),
    .B(_0851_));
 sg13g2_and3_2 _4681_ (.X(_1059_),
    .A(_1056_),
    .B(_1057_),
    .C(_1058_));
 sg13g2_nand3_1 _4682_ (.B(_1057_),
    .C(_1058_),
    .A(_1056_),
    .Y(_1060_));
 sg13g2_nor3_1 _4683_ (.A(\led_controller.cpu.current_instruction[15] ),
    .B(\led_controller.cpu.current_instruction[14] ),
    .C(\led_controller.cpu.current_instruction[13] ),
    .Y(_1061_));
 sg13g2_and2_1 _4684_ (.A(_0843_),
    .B(_1061_),
    .X(_1062_));
 sg13g2_nand2_2 _4685_ (.Y(_1063_),
    .A(_0843_),
    .B(_1061_));
 sg13g2_nand4_1 _4686_ (.B(net1840),
    .C(net2055),
    .A(net1941),
    .Y(_1064_),
    .D(_1062_));
 sg13g2_xnor2_1 _4687_ (.Y(_1065_),
    .A(\led_controller.cpu.current_instruction_pc[11] ),
    .B(\led_controller.cpu.pc[11] ));
 sg13g2_xor2_1 _4688_ (.B(\led_controller.cpu.pc[7] ),
    .A(\led_controller.cpu.current_instruction_pc[7] ),
    .X(_1066_));
 sg13g2_xnor2_1 _4689_ (.Y(_1067_),
    .A(\led_controller.cpu.current_instruction_pc[8] ),
    .B(\led_controller.cpu.pc[8] ));
 sg13g2_xor2_1 _4690_ (.B(\led_controller.cpu.pc[2] ),
    .A(\led_controller.cpu.current_instruction_pc[2] ),
    .X(_1068_));
 sg13g2_xnor2_1 _4691_ (.Y(_1069_),
    .A(\led_controller.cpu.current_instruction_pc[12] ),
    .B(\led_controller.cpu.pc[12] ));
 sg13g2_xor2_1 _4692_ (.B(\led_controller.cpu.pc[5] ),
    .A(\led_controller.cpu.current_instruction_pc[5] ),
    .X(_1070_));
 sg13g2_xor2_1 _4693_ (.B(\led_controller.cpu.pc[10] ),
    .A(\led_controller.cpu.current_instruction_pc[10] ),
    .X(_1071_));
 sg13g2_xor2_1 _4694_ (.B(\led_controller.cpu.pc[1] ),
    .A(\led_controller.cpu.current_instruction_pc[1] ),
    .X(_1072_));
 sg13g2_xor2_1 _4695_ (.B(\led_controller.cpu.pc[13] ),
    .A(\led_controller.cpu.current_instruction_pc[13] ),
    .X(_1073_));
 sg13g2_xor2_1 _4696_ (.B(\led_controller.cpu.pc[14] ),
    .A(\led_controller.cpu.current_instruction_pc[14] ),
    .X(_1074_));
 sg13g2_nor4_1 _4697_ (.A(_1066_),
    .B(_1070_),
    .C(_1071_),
    .D(_1073_),
    .Y(_1075_));
 sg13g2_xor2_1 _4698_ (.B(\led_controller.cpu.pc[3] ),
    .A(\led_controller.cpu.current_instruction_pc[3] ),
    .X(_1076_));
 sg13g2_nor4_1 _4699_ (.A(_1068_),
    .B(_1072_),
    .C(_1074_),
    .D(_1076_),
    .Y(_1077_));
 sg13g2_a22oi_1 _4700_ (.Y(_1078_),
    .B1(\led_controller.cpu.pc[4] ),
    .B2(_0836_),
    .A2(\led_controller.cpu.pc[6] ),
    .A1(_0834_));
 sg13g2_xnor2_1 _4701_ (.Y(_1079_),
    .A(\led_controller.cpu.current_instruction_pc[0] ),
    .B(\led_controller.cpu.pc[0] ));
 sg13g2_nand4_1 _4702_ (.B(_1067_),
    .C(_1078_),
    .A(_1065_),
    .Y(_1080_),
    .D(_1079_));
 sg13g2_xnor2_1 _4703_ (.Y(_1081_),
    .A(\led_controller.cpu.current_instruction_pc[15] ),
    .B(\led_controller.cpu.pc[15] ));
 sg13g2_xnor2_1 _4704_ (.Y(_1082_),
    .A(\led_controller.cpu.current_instruction_pc[9] ),
    .B(\led_controller.cpu.pc[9] ));
 sg13g2_a22oi_1 _4705_ (.Y(_1083_),
    .B1(_0869_),
    .B2(\led_controller.cpu.current_instruction_pc[4] ),
    .A2(_0868_),
    .A1(\led_controller.cpu.current_instruction_pc[6] ));
 sg13g2_nand4_1 _4706_ (.B(_1081_),
    .C(_1082_),
    .A(_1069_),
    .Y(_1084_),
    .D(_1083_));
 sg13g2_nor2_1 _4707_ (.A(_1080_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nand3_1 _4708_ (.B(_1077_),
    .C(_1085_),
    .A(_1075_),
    .Y(_1086_));
 sg13g2_nor2_1 _4709_ (.A(net2138),
    .B(net1635),
    .Y(_1087_));
 sg13g2_nand2_2 _4710_ (.Y(_1088_),
    .A(net1434),
    .B(_1087_));
 sg13g2_nor3_1 _4711_ (.A(net2142),
    .B(\led_controller.cpu.stall_counter[1] ),
    .C(\led_controller.cpu.stall_counter[0] ),
    .Y(_1089_));
 sg13g2_nor2b_1 _4712_ (.A(net1626),
    .B_N(_1089_),
    .Y(_1090_));
 sg13g2_nor3_1 _4713_ (.A(\led_controller.cpu.stall_counter[6] ),
    .B(\led_controller.cpu.stall_counter[5] ),
    .C(\led_controller.cpu.stall_counter[4] ),
    .Y(_1091_));
 sg13g2_nand2_1 _4714_ (.Y(_1092_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_nand3_1 _4715_ (.B(_1090_),
    .C(_1091_),
    .A(_0857_),
    .Y(_1093_));
 sg13g2_nor4_2 _4716_ (.A(net2364),
    .B(_1086_),
    .C(_1088_),
    .Y(_1094_),
    .D(_1093_));
 sg13g2_inv_4 _4717_ (.A(_1094_),
    .Y(_1095_));
 sg13g2_nor4_1 _4718_ (.A(net1031),
    .B(_1060_),
    .C(_1064_),
    .D(_1095_),
    .Y(_1096_));
 sg13g2_nand3_1 _4719_ (.B(\led_controller.cpu.current_instruction[2] ),
    .C(_1096_),
    .A(\led_controller.cpu.current_instruction[3] ),
    .Y(_1097_));
 sg13g2_nor4_2 _4720_ (.A(\led_controller.cpu.led_write_strb ),
    .B(_1086_),
    .C(_1088_),
    .Y(_1098_),
    .D(_1093_));
 sg13g2_nand2b_1 _4721_ (.Y(_1099_),
    .B(_1098_),
    .A_N(_1064_));
 sg13g2_nor3_1 _4722_ (.A(net1031),
    .B(_1060_),
    .C(_1099_),
    .Y(_1100_));
 sg13g2_nand3_1 _4723_ (.B(net2389),
    .C(_1100_),
    .A(\led_controller.cpu.current_instruction[3] ),
    .Y(_1101_));
 sg13g2_or2_1 _4724_ (.X(_1102_),
    .B(_1101_),
    .A(_1051_));
 sg13g2_or4_1 _4725_ (.A(\led_controller.cpu.led_write_strb ),
    .B(_1086_),
    .C(_1088_),
    .D(_1093_),
    .X(_1103_));
 sg13g2_or4_1 _4726_ (.A(net1033),
    .B(_1060_),
    .C(_1064_),
    .D(net876),
    .X(_1104_));
 sg13g2_and2_1 _4727_ (.A(net1060),
    .B(_1102_),
    .X(_1105_));
 sg13g2_nand2_1 _4728_ (.Y(_1106_),
    .A(net1274),
    .B(_1105_));
 sg13g2_nor2_2 _4729_ (.A(\led_controller.cpu.current_instruction[8] ),
    .B(_1064_),
    .Y(_1107_));
 sg13g2_nor2_2 _4730_ (.A(_0847_),
    .B(_1064_),
    .Y(_1108_));
 sg13g2_a22oi_1 _4731_ (.Y(_1109_),
    .B1(_1108_),
    .B2(net1185),
    .A2(_1107_),
    .A1(\led_controller.cpu.register_y[0] ));
 sg13g2_o21ai_1 _4732_ (.B1(_1106_),
    .Y(_0024_),
    .A1(_1102_),
    .A2(net934));
 sg13g2_nand2_1 _4733_ (.Y(_1110_),
    .A(net802),
    .B(_1105_));
 sg13g2_a22oi_1 _4734_ (.Y(_1111_),
    .B1(_1108_),
    .B2(net1184),
    .A2(_1107_),
    .A1(net1180));
 sg13g2_o21ai_1 _4735_ (.B1(_1110_),
    .Y(_0025_),
    .A1(_1102_),
    .A2(net933));
 sg13g2_nand2_1 _4736_ (.Y(_1112_),
    .A(net1404),
    .B(_1105_));
 sg13g2_a22oi_1 _4737_ (.Y(_1113_),
    .B1(_1108_),
    .B2(net1183),
    .A2(_1107_),
    .A1(\led_controller.cpu.register_y[2] ));
 sg13g2_o21ai_1 _4738_ (.B1(_1112_),
    .Y(_0026_),
    .A1(_1102_),
    .A2(net929));
 sg13g2_nand2_1 _4739_ (.Y(_1114_),
    .A(net780),
    .B(_1105_));
 sg13g2_a22oi_1 _4740_ (.Y(_1115_),
    .B1(_1108_),
    .B2(\led_controller.cpu.register_x[3] ),
    .A2(_1107_),
    .A1(\led_controller.cpu.register_y[3] ));
 sg13g2_o21ai_1 _4741_ (.B1(_1114_),
    .Y(_0027_),
    .A1(_1102_),
    .A2(net926));
 sg13g2_nand2_1 _4742_ (.Y(_1116_),
    .A(net775),
    .B(_1105_));
 sg13g2_a22oi_1 _4743_ (.Y(_1117_),
    .B1(_1108_),
    .B2(net1182),
    .A2(_1107_),
    .A1(\led_controller.cpu.register_y[4] ));
 sg13g2_o21ai_1 _4744_ (.B1(_1116_),
    .Y(_0028_),
    .A1(_1102_),
    .A2(net925));
 sg13g2_a22oi_1 _4745_ (.Y(_1118_),
    .B1(_1108_),
    .B2(\led_controller.cpu.register_x[5] ),
    .A2(_1107_),
    .A1(net1178));
 sg13g2_nor3_1 _4746_ (.A(_1051_),
    .B(_1097_),
    .C(net922),
    .Y(_1119_));
 sg13g2_a21o_1 _4747_ (.A2(_1105_),
    .A1(net1533),
    .B1(_1119_),
    .X(_0029_));
 sg13g2_nand2_1 _4748_ (.Y(_1120_),
    .A(net1292),
    .B(_1105_));
 sg13g2_a22oi_1 _4749_ (.Y(_1121_),
    .B1(_1108_),
    .B2(net2392),
    .A2(_1107_),
    .A1(\led_controller.cpu.register_y[6] ));
 sg13g2_o21ai_1 _4750_ (.B1(_1120_),
    .Y(_0030_),
    .A1(_1102_),
    .A2(net918));
 sg13g2_nand2_1 _4751_ (.Y(_1122_),
    .A(net787),
    .B(_1105_));
 sg13g2_a22oi_1 _4752_ (.Y(_1123_),
    .B1(_1108_),
    .B2(\led_controller.cpu.register_x[7] ),
    .A2(_1107_),
    .A1(\led_controller.cpu.register_y[7] ));
 sg13g2_o21ai_1 _4753_ (.B1(_1122_),
    .Y(_0031_),
    .A1(_1102_),
    .A2(net917));
 sg13g2_nor2_2 _4754_ (.A(\led_controller.cpu.current_instruction[1] ),
    .B(_0855_),
    .Y(_1124_));
 sg13g2_and3_2 _4755_ (.X(_1125_),
    .A(\led_controller.cpu.current_instruction[3] ),
    .B(_0853_),
    .C(_1096_));
 sg13g2_nand2_2 _4756_ (.Y(_1126_),
    .A(_1124_),
    .B(_1125_));
 sg13g2_nor3_2 _4757_ (.A(_0852_),
    .B(\led_controller.cpu.current_instruction[2] ),
    .C(_1104_),
    .Y(_1127_));
 sg13g2_a21oi_2 _4758_ (.B1(net1031),
    .Y(_1128_),
    .A2(_1127_),
    .A1(_1124_));
 sg13g2_nand2_1 _4759_ (.Y(_1129_),
    .A(net1310),
    .B(_1128_));
 sg13g2_o21ai_1 _4760_ (.B1(_1129_),
    .Y(_0032_),
    .A1(net934),
    .A2(_1126_));
 sg13g2_nand2_1 _4761_ (.Y(_1130_),
    .A(net1239),
    .B(_1128_));
 sg13g2_o21ai_1 _4762_ (.B1(_1130_),
    .Y(_0033_),
    .A1(net931),
    .A2(_1126_));
 sg13g2_nand2_1 _4763_ (.Y(_1131_),
    .A(net800),
    .B(_1128_));
 sg13g2_o21ai_1 _4764_ (.B1(_1131_),
    .Y(_0034_),
    .A1(net929),
    .A2(_1126_));
 sg13g2_nand2_1 _4765_ (.Y(_1132_),
    .A(net1241),
    .B(_1128_));
 sg13g2_o21ai_1 _4766_ (.B1(_1132_),
    .Y(_0035_),
    .A1(net927),
    .A2(_1126_));
 sg13g2_nand2_1 _4767_ (.Y(_1133_),
    .A(net1284),
    .B(_1128_));
 sg13g2_o21ai_1 _4768_ (.B1(_1133_),
    .Y(_0036_),
    .A1(net924),
    .A2(_1126_));
 sg13g2_nand2_1 _4769_ (.Y(_1134_),
    .A(net1250),
    .B(_1128_));
 sg13g2_o21ai_1 _4770_ (.B1(_1134_),
    .Y(_0037_),
    .A1(net921),
    .A2(_1126_));
 sg13g2_nand2_1 _4771_ (.Y(_1135_),
    .A(net1290),
    .B(_1128_));
 sg13g2_o21ai_1 _4772_ (.B1(_1135_),
    .Y(_0038_),
    .A1(net918),
    .A2(_1126_));
 sg13g2_nand2_1 _4773_ (.Y(_1136_),
    .A(net793),
    .B(_1128_));
 sg13g2_o21ai_1 _4774_ (.B1(_1136_),
    .Y(_0039_),
    .A1(net916),
    .A2(_1126_));
 sg13g2_nand2_2 _4775_ (.Y(_1137_),
    .A(\led_controller.cpu.current_instruction[1] ),
    .B(\led_controller.cpu.current_instruction[0] ));
 sg13g2_nand3_1 _4776_ (.B(\led_controller.cpu.current_instruction[0] ),
    .C(_1127_),
    .A(\led_controller.cpu.current_instruction[1] ),
    .Y(_1138_));
 sg13g2_and2_1 _4777_ (.A(net1060),
    .B(_1138_),
    .X(_1139_));
 sg13g2_nand2_1 _4778_ (.Y(_1140_),
    .A(net1297),
    .B(_1139_));
 sg13g2_o21ai_1 _4779_ (.B1(_1140_),
    .Y(_0040_),
    .A1(net935),
    .A2(net831));
 sg13g2_nand2_1 _4780_ (.Y(_1141_),
    .A(net1226),
    .B(_1139_));
 sg13g2_o21ai_1 _4781_ (.B1(_1141_),
    .Y(_0041_),
    .A1(net932),
    .A2(net831));
 sg13g2_nand2_1 _4782_ (.Y(_1142_),
    .A(net803),
    .B(_1139_));
 sg13g2_o21ai_1 _4783_ (.B1(_1142_),
    .Y(_0042_),
    .A1(net929),
    .A2(net831));
 sg13g2_nand2_1 _4784_ (.Y(_1143_),
    .A(net1263),
    .B(_1139_));
 sg13g2_o21ai_1 _4785_ (.B1(_1143_),
    .Y(_0043_),
    .A1(net926),
    .A2(net831));
 sg13g2_nand2_1 _4786_ (.Y(_1144_),
    .A(net812),
    .B(_1139_));
 sg13g2_o21ai_1 _4787_ (.B1(_1144_),
    .Y(_0044_),
    .A1(net924),
    .A2(net831));
 sg13g2_nand2_1 _4788_ (.Y(_1145_),
    .A(net1361),
    .B(_1139_));
 sg13g2_o21ai_1 _4789_ (.B1(_1145_),
    .Y(_0045_),
    .A1(net921),
    .A2(net831));
 sg13g2_nand2_1 _4790_ (.Y(_1146_),
    .A(net1364),
    .B(_1139_));
 sg13g2_o21ai_1 _4791_ (.B1(_1146_),
    .Y(_0046_),
    .A1(net918),
    .A2(net831));
 sg13g2_nand2_1 _4792_ (.Y(_1147_),
    .A(net1301),
    .B(_1139_));
 sg13g2_o21ai_1 _4793_ (.B1(_1147_),
    .Y(_0047_),
    .A1(net916),
    .A2(net831));
 sg13g2_nand2_2 _4794_ (.Y(_1148_),
    .A(_1050_),
    .B(_1125_));
 sg13g2_a21oi_2 _4795_ (.B1(net1031),
    .Y(_1149_),
    .A2(_1127_),
    .A1(_1050_));
 sg13g2_nand2_1 _4796_ (.Y(_1150_),
    .A(net806),
    .B(_1149_));
 sg13g2_o21ai_1 _4797_ (.B1(_1150_),
    .Y(_0048_),
    .A1(net935),
    .A2(_1148_));
 sg13g2_nand2_1 _4798_ (.Y(_1151_),
    .A(net1327),
    .B(_1149_));
 sg13g2_o21ai_1 _4799_ (.B1(_1151_),
    .Y(_0049_),
    .A1(net932),
    .A2(_1148_));
 sg13g2_nand2_1 _4800_ (.Y(_1152_),
    .A(net767),
    .B(_1149_));
 sg13g2_o21ai_1 _4801_ (.B1(_1152_),
    .Y(_0050_),
    .A1(net929),
    .A2(_1148_));
 sg13g2_nand2_1 _4802_ (.Y(_1153_),
    .A(net777),
    .B(_1149_));
 sg13g2_o21ai_1 _4803_ (.B1(_1153_),
    .Y(_0051_),
    .A1(net926),
    .A2(_1148_));
 sg13g2_nand2_1 _4804_ (.Y(_1154_),
    .A(net1331),
    .B(_1149_));
 sg13g2_o21ai_1 _4805_ (.B1(_1154_),
    .Y(_0052_),
    .A1(net924),
    .A2(_1148_));
 sg13g2_nand2_1 _4806_ (.Y(_1155_),
    .A(net1387),
    .B(_1149_));
 sg13g2_o21ai_1 _4807_ (.B1(_1155_),
    .Y(_0053_),
    .A1(net921),
    .A2(_1148_));
 sg13g2_nand2_1 _4808_ (.Y(_1156_),
    .A(net796),
    .B(_1149_));
 sg13g2_o21ai_1 _4809_ (.B1(_1156_),
    .Y(_0054_),
    .A1(net918),
    .A2(_1148_));
 sg13g2_nand2_1 _4810_ (.Y(_1157_),
    .A(net773),
    .B(_1149_));
 sg13g2_o21ai_1 _4811_ (.B1(_1157_),
    .Y(_0055_),
    .A1(net916),
    .A2(_1148_));
 sg13g2_nor3_2 _4812_ (.A(\led_controller.cpu.current_instruction[3] ),
    .B(_0853_),
    .C(_1104_),
    .Y(_1158_));
 sg13g2_nand2_2 _4813_ (.Y(_1159_),
    .A(_1124_),
    .B(_1158_));
 sg13g2_a21oi_2 _4814_ (.B1(net1031),
    .Y(_1160_),
    .A2(_1158_),
    .A1(_1124_));
 sg13g2_nand2_1 _4815_ (.Y(_1161_),
    .A(net1317),
    .B(_1160_));
 sg13g2_o21ai_1 _4816_ (.B1(_1161_),
    .Y(_0056_),
    .A1(net934),
    .A2(_1159_));
 sg13g2_nand2_1 _4817_ (.Y(_1162_),
    .A(net1254),
    .B(_1160_));
 sg13g2_o21ai_1 _4818_ (.B1(_1162_),
    .Y(_0057_),
    .A1(net931),
    .A2(_1159_));
 sg13g2_nand2_1 _4819_ (.Y(_1163_),
    .A(net1337),
    .B(_1160_));
 sg13g2_o21ai_1 _4820_ (.B1(_1163_),
    .Y(_0058_),
    .A1(net930),
    .A2(_1159_));
 sg13g2_nand2_1 _4821_ (.Y(_1164_),
    .A(net1271),
    .B(_1160_));
 sg13g2_o21ai_1 _4822_ (.B1(_1164_),
    .Y(_0059_),
    .A1(net926),
    .A2(_1159_));
 sg13g2_nand2_1 _4823_ (.Y(_1165_),
    .A(net1300),
    .B(_1160_));
 sg13g2_o21ai_1 _4824_ (.B1(_1165_),
    .Y(_0060_),
    .A1(net925),
    .A2(_1159_));
 sg13g2_nand2_1 _4825_ (.Y(_1166_),
    .A(net798),
    .B(_1160_));
 sg13g2_o21ai_1 _4826_ (.B1(_1166_),
    .Y(_0061_),
    .A1(net921),
    .A2(_1159_));
 sg13g2_nand2_1 _4827_ (.Y(_1167_),
    .A(net1238),
    .B(_1160_));
 sg13g2_o21ai_1 _4828_ (.B1(_1167_),
    .Y(_0062_),
    .A1(net918),
    .A2(_1159_));
 sg13g2_nand2_1 _4829_ (.Y(_1168_),
    .A(net1282),
    .B(_1160_));
 sg13g2_o21ai_1 _4830_ (.B1(_1168_),
    .Y(_0063_),
    .A1(net917),
    .A2(_1159_));
 sg13g2_nor2_1 _4831_ (.A(net2095),
    .B(_0945_),
    .Y(_1169_));
 sg13g2_nor2_1 _4832_ (.A(\led_controller.timer_100hz.div_counter[1] ),
    .B(_0950_),
    .Y(_1170_));
 sg13g2_a22oi_1 _4833_ (.Y(_1171_),
    .B1(\led_controller.timer_100hz.div_counter[1] ),
    .B2(_0950_),
    .A2(\led_controller.timer_100hz.div_counter[0] ),
    .A1(\led_controller.clock_divider[0] ));
 sg13g2_o21ai_1 _4834_ (.B1(_1171_),
    .Y(_1172_),
    .A1(\led_controller.clock_divider[0] ),
    .A2(\led_controller.timer_100hz.div_counter[0] ));
 sg13g2_xnor2_1 _4835_ (.Y(_1173_),
    .A(\led_controller.timer_100hz.div_counter[2] ),
    .B(_0954_));
 sg13g2_xnor2_1 _4836_ (.Y(_1174_),
    .A(\led_controller.timer_100hz.div_counter[3] ),
    .B(_0948_));
 sg13g2_nor4_1 _4837_ (.A(_1170_),
    .B(_1172_),
    .C(_1173_),
    .D(_1174_),
    .Y(_1175_));
 sg13g2_xor2_1 _4838_ (.B(_0959_),
    .A(net1793),
    .X(_1176_));
 sg13g2_xnor2_1 _4839_ (.Y(_1177_),
    .A(\led_controller.timer_100hz.div_counter[6] ),
    .B(_0944_));
 sg13g2_a21o_1 _4840_ (.A2(_0945_),
    .A1(net2095),
    .B1(_1177_),
    .X(_1178_));
 sg13g2_xor2_1 _4841_ (.B(_0958_),
    .A(net1878),
    .X(_1179_));
 sg13g2_nand3_1 _4842_ (.B(_1176_),
    .C(_1179_),
    .A(_1175_),
    .Y(_1180_));
 sg13g2_nor4_2 _4843_ (.A(_0947_),
    .B(_1169_),
    .C(_1178_),
    .Y(_1181_),
    .D(_1180_));
 sg13g2_nand2b_2 _4844_ (.Y(_1182_),
    .B(net1158),
    .A_N(_1181_));
 sg13g2_nor2_1 _4845_ (.A(net1280),
    .B(_1182_),
    .Y(_0064_));
 sg13g2_xnor2_1 _4846_ (.Y(_1183_),
    .A(net1280),
    .B(net1930));
 sg13g2_nor2_1 _4847_ (.A(_1182_),
    .B(_1183_),
    .Y(_0065_));
 sg13g2_and3_1 _4848_ (.X(_1184_),
    .A(net1280),
    .B(net2391),
    .C(net1514));
 sg13g2_a21oi_1 _4849_ (.A1(net1280),
    .A2(\led_controller.timer_100hz.div_counter[1] ),
    .Y(_1185_),
    .B1(net1514));
 sg13g2_nor3_1 _4850_ (.A(_1182_),
    .B(_1184_),
    .C(net1515),
    .Y(_0066_));
 sg13g2_and2_1 _4851_ (.A(net1843),
    .B(_1184_),
    .X(_1186_));
 sg13g2_nor2_1 _4852_ (.A(net1843),
    .B(_1184_),
    .Y(_1187_));
 sg13g2_nor3_1 _4853_ (.A(_1182_),
    .B(_1186_),
    .C(net1844),
    .Y(_0067_));
 sg13g2_and2_1 _4854_ (.A(net1793),
    .B(_1186_),
    .X(_1188_));
 sg13g2_nor2_1 _4855_ (.A(net1793),
    .B(_1186_),
    .Y(_1189_));
 sg13g2_nor3_1 _4856_ (.A(_1182_),
    .B(_1188_),
    .C(net1794),
    .Y(_0068_));
 sg13g2_and2_1 _4857_ (.A(net1878),
    .B(_1188_),
    .X(_1190_));
 sg13g2_nor2_1 _4858_ (.A(net1878),
    .B(_1188_),
    .Y(_1191_));
 sg13g2_nor3_1 _4859_ (.A(_1182_),
    .B(_1190_),
    .C(_1191_),
    .Y(_0069_));
 sg13g2_nand2_1 _4860_ (.Y(_1192_),
    .A(net1974),
    .B(_1190_));
 sg13g2_xnor2_1 _4861_ (.Y(_1193_),
    .A(net1974),
    .B(_1190_));
 sg13g2_nor2_1 _4862_ (.A(_1182_),
    .B(_1193_),
    .Y(_0070_));
 sg13g2_xor2_1 _4863_ (.B(_1192_),
    .A(net2095),
    .X(_1194_));
 sg13g2_nor2_1 _4864_ (.A(_1182_),
    .B(_1194_),
    .Y(_0071_));
 sg13g2_nand2_2 _4865_ (.Y(_1195_),
    .A(_1052_),
    .B(_1158_));
 sg13g2_a21oi_2 _4866_ (.B1(net1031),
    .Y(_1196_),
    .A2(_1158_),
    .A1(_1052_));
 sg13g2_nand2_1 _4867_ (.Y(_1197_),
    .A(net788),
    .B(_1196_));
 sg13g2_o21ai_1 _4868_ (.B1(_1197_),
    .Y(_0072_),
    .A1(net934),
    .A2(_1195_));
 sg13g2_nand2_1 _4869_ (.Y(_1198_),
    .A(net1341),
    .B(_1196_));
 sg13g2_o21ai_1 _4870_ (.B1(_1198_),
    .Y(_0073_),
    .A1(net931),
    .A2(_1195_));
 sg13g2_nand2_1 _4871_ (.Y(_1199_),
    .A(net1255),
    .B(_1196_));
 sg13g2_o21ai_1 _4872_ (.B1(_1199_),
    .Y(_0074_),
    .A1(net930),
    .A2(_1195_));
 sg13g2_nand2_1 _4873_ (.Y(_1200_),
    .A(net819),
    .B(_1196_));
 sg13g2_o21ai_1 _4874_ (.B1(_1200_),
    .Y(_0075_),
    .A1(net926),
    .A2(_1195_));
 sg13g2_nand2_1 _4875_ (.Y(_1201_),
    .A(net1275),
    .B(_1196_));
 sg13g2_o21ai_1 _4876_ (.B1(_1201_),
    .Y(_0076_),
    .A1(net925),
    .A2(_1195_));
 sg13g2_nand2_1 _4877_ (.Y(_1202_),
    .A(net1308),
    .B(_1196_));
 sg13g2_o21ai_1 _4878_ (.B1(_1202_),
    .Y(_0077_),
    .A1(net921),
    .A2(_1195_));
 sg13g2_nand2_1 _4879_ (.Y(_1203_),
    .A(net795),
    .B(_1196_));
 sg13g2_o21ai_1 _4880_ (.B1(_1203_),
    .Y(_0078_),
    .A1(net918),
    .A2(_1195_));
 sg13g2_nand2_1 _4881_ (.Y(_1204_),
    .A(net1262),
    .B(_1196_));
 sg13g2_o21ai_1 _4882_ (.B1(_1204_),
    .Y(_0079_),
    .A1(net916),
    .A2(_1195_));
 sg13g2_and2_1 _4883_ (.A(_1054_),
    .B(_1100_),
    .X(_1205_));
 sg13g2_nand2b_2 _4884_ (.Y(_1206_),
    .B(_1205_),
    .A_N(_1137_));
 sg13g2_and2_1 _4885_ (.A(net1059),
    .B(net825),
    .X(_1207_));
 sg13g2_nand2_1 _4886_ (.Y(_1208_),
    .A(net1347),
    .B(_1207_));
 sg13g2_o21ai_1 _4887_ (.B1(_1208_),
    .Y(_0080_),
    .A1(net936),
    .A2(_1206_));
 sg13g2_nand2_1 _4888_ (.Y(_1209_),
    .A(net1395),
    .B(_1207_));
 sg13g2_o21ai_1 _4889_ (.B1(_1209_),
    .Y(_0081_),
    .A1(net931),
    .A2(net825));
 sg13g2_nand2_1 _4890_ (.Y(_1210_),
    .A(net1377),
    .B(_1207_));
 sg13g2_o21ai_1 _4891_ (.B1(_1210_),
    .Y(_0082_),
    .A1(net930),
    .A2(net825));
 sg13g2_nand2_1 _4892_ (.Y(_1211_),
    .A(net1299),
    .B(_1207_));
 sg13g2_o21ai_1 _4893_ (.B1(_1211_),
    .Y(_0083_),
    .A1(net928),
    .A2(net825));
 sg13g2_nand2_1 _4894_ (.Y(_1212_),
    .A(net1270),
    .B(_1207_));
 sg13g2_o21ai_1 _4895_ (.B1(_1212_),
    .Y(_0084_),
    .A1(net924),
    .A2(net825));
 sg13g2_nand2_1 _4896_ (.Y(_1213_),
    .A(net1324),
    .B(_1207_));
 sg13g2_o21ai_1 _4897_ (.B1(_1213_),
    .Y(_0085_),
    .A1(net923),
    .A2(net825));
 sg13g2_nand2_1 _4898_ (.Y(_1214_),
    .A(net1273),
    .B(_1207_));
 sg13g2_o21ai_1 _4899_ (.B1(_1214_),
    .Y(_0086_),
    .A1(net920),
    .A2(net825));
 sg13g2_nand2_1 _4900_ (.Y(_1215_),
    .A(net1338),
    .B(_1207_));
 sg13g2_o21ai_1 _4901_ (.B1(_1215_),
    .Y(_0087_),
    .A1(net916),
    .A2(net825));
 sg13g2_or2_1 _4902_ (.X(_1216_),
    .B(net2390),
    .A(_1053_));
 sg13g2_and2_1 _4903_ (.A(net1060),
    .B(net824),
    .X(_1217_));
 sg13g2_nand2_1 _4904_ (.Y(_1218_),
    .A(net1228),
    .B(_1217_));
 sg13g2_o21ai_1 _4905_ (.B1(_1218_),
    .Y(_0088_),
    .A1(net935),
    .A2(net824));
 sg13g2_nand2_1 _4906_ (.Y(_1219_),
    .A(net784),
    .B(_1217_));
 sg13g2_o21ai_1 _4907_ (.B1(_1219_),
    .Y(_0089_),
    .A1(net933),
    .A2(_1216_));
 sg13g2_nand2_1 _4908_ (.Y(_1220_),
    .A(net1349),
    .B(_1217_));
 sg13g2_o21ai_1 _4909_ (.B1(_1220_),
    .Y(_0090_),
    .A1(net929),
    .A2(net824));
 sg13g2_nand2_1 _4910_ (.Y(_1221_),
    .A(net1267),
    .B(_1217_));
 sg13g2_o21ai_1 _4911_ (.B1(_1221_),
    .Y(_0091_),
    .A1(net927),
    .A2(net824));
 sg13g2_nand2_1 _4912_ (.Y(_1222_),
    .A(net1372),
    .B(_1217_));
 sg13g2_o21ai_1 _4913_ (.B1(_1222_),
    .Y(_0092_),
    .A1(net925),
    .A2(net824));
 sg13g2_nand2_1 _4914_ (.Y(_1223_),
    .A(net811),
    .B(_1217_));
 sg13g2_o21ai_1 _4915_ (.B1(_1223_),
    .Y(_0093_),
    .A1(net922),
    .A2(net824));
 sg13g2_nand2_1 _4916_ (.Y(_1224_),
    .A(net1260),
    .B(_1217_));
 sg13g2_o21ai_1 _4917_ (.B1(_1224_),
    .Y(_0094_),
    .A1(net918),
    .A2(net824));
 sg13g2_nand2_1 _4918_ (.Y(_1225_),
    .A(net1287),
    .B(_1217_));
 sg13g2_o21ai_1 _4919_ (.B1(_1225_),
    .Y(_0095_),
    .A1(net917),
    .A2(net824));
 sg13g2_and2_1 _4920_ (.A(_0856_),
    .B(_1086_),
    .X(_1226_));
 sg13g2_and2_1 _4921_ (.A(_1043_),
    .B(_1226_),
    .X(_1227_));
 sg13g2_nand2_1 _4922_ (.Y(_1228_),
    .A(net1186),
    .B(net848));
 sg13g2_nand2_1 _4923_ (.Y(_1229_),
    .A(net2339),
    .B(net948));
 sg13g2_nor2b_1 _4924_ (.A(net848),
    .B_N(_1229_),
    .Y(_1230_));
 sg13g2_o21ai_1 _4925_ (.B1(_1230_),
    .Y(_1231_),
    .A1(net2339),
    .A2(net948));
 sg13g2_a21oi_1 _4926_ (.A1(_1228_),
    .A2(_1231_),
    .Y(_0096_),
    .B1(net1039));
 sg13g2_xor2_1 _4927_ (.B(\led_controller.cpu.fetch_pc[1] ),
    .A(net2216),
    .X(_1232_));
 sg13g2_a22oi_1 _4928_ (.Y(_1233_),
    .B1(_1232_),
    .B2(net949),
    .A2(net848),
    .A1(\led_controller.cpu.pc[2] ));
 sg13g2_nor2_1 _4929_ (.A(net1039),
    .B(_1233_),
    .Y(_1234_));
 sg13g2_nor2_1 _4930_ (.A(net950),
    .B(net847),
    .Y(_1235_));
 sg13g2_or2_1 _4931_ (.X(_1236_),
    .B(net847),
    .A(net950));
 sg13g2_nor2_1 _4932_ (.A(net1038),
    .B(_1236_),
    .Y(_1237_));
 sg13g2_a21o_1 _4933_ (.A2(net829),
    .A1(net2216),
    .B1(_1234_),
    .X(_0097_));
 sg13g2_nand3_1 _4934_ (.B(\led_controller.cpu.fetch_pc[2] ),
    .C(\led_controller.cpu.fetch_pc[1] ),
    .A(\led_controller.cpu.fetch_pc[3] ),
    .Y(_1238_));
 sg13g2_a21o_1 _4935_ (.A2(\led_controller.cpu.fetch_pc[1] ),
    .A1(\led_controller.cpu.fetch_pc[2] ),
    .B1(\led_controller.cpu.fetch_pc[3] ),
    .X(_1239_));
 sg13g2_and2_1 _4936_ (.A(_1238_),
    .B(_1239_),
    .X(_1240_));
 sg13g2_a22oi_1 _4937_ (.Y(_1241_),
    .B1(_1240_),
    .B2(net949),
    .A2(net848),
    .A1(\led_controller.cpu.pc[3] ));
 sg13g2_nor2_1 _4938_ (.A(net1039),
    .B(_1241_),
    .Y(_1242_));
 sg13g2_a21o_1 _4939_ (.A2(net829),
    .A1(net2009),
    .B1(_1242_),
    .X(_0098_));
 sg13g2_nor2_1 _4940_ (.A(_0837_),
    .B(_1238_),
    .Y(_1243_));
 sg13g2_xnor2_1 _4941_ (.Y(_1244_),
    .A(net2155),
    .B(_1238_));
 sg13g2_a22oi_1 _4942_ (.Y(_1245_),
    .B1(_1244_),
    .B2(net949),
    .A2(net849),
    .A1(\led_controller.cpu.pc[4] ));
 sg13g2_nor2_1 _4943_ (.A(net1037),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_a21o_1 _4944_ (.A2(net830),
    .A1(net2155),
    .B1(_1246_),
    .X(_0099_));
 sg13g2_xor2_1 _4945_ (.B(_1243_),
    .A(net2226),
    .X(_1247_));
 sg13g2_a22oi_1 _4946_ (.Y(_1248_),
    .B1(_1247_),
    .B2(net948),
    .A2(net848),
    .A1(\led_controller.cpu.pc[5] ));
 sg13g2_nor2_1 _4947_ (.A(net1037),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_a21o_1 _4948_ (.A2(net829),
    .A1(net2226),
    .B1(_1249_),
    .X(_0100_));
 sg13g2_a21oi_1 _4949_ (.A1(\led_controller.cpu.fetch_pc[5] ),
    .A2(_1243_),
    .Y(_1250_),
    .B1(net1924));
 sg13g2_nand3_1 _4950_ (.B(\led_controller.cpu.fetch_pc[5] ),
    .C(_1243_),
    .A(\led_controller.cpu.fetch_pc[6] ),
    .Y(_1251_));
 sg13g2_nor2b_1 _4951_ (.A(_1250_),
    .B_N(_1251_),
    .Y(_1252_));
 sg13g2_a22oi_1 _4952_ (.Y(_1253_),
    .B1(_1252_),
    .B2(net949),
    .A2(net848),
    .A1(\led_controller.cpu.pc[6] ));
 sg13g2_nand2_1 _4953_ (.Y(_1254_),
    .A(net1924),
    .B(net835));
 sg13g2_a21oi_1 _4954_ (.A1(_1253_),
    .A2(_1254_),
    .Y(_0101_),
    .B1(net1038));
 sg13g2_nor2_1 _4955_ (.A(_0833_),
    .B(_1251_),
    .Y(_1255_));
 sg13g2_xnor2_1 _4956_ (.Y(_1256_),
    .A(net1834),
    .B(_1251_));
 sg13g2_a22oi_1 _4957_ (.Y(_1257_),
    .B1(_1256_),
    .B2(net950),
    .A2(net848),
    .A1(\led_controller.cpu.pc[7] ));
 sg13g2_nand2_1 _4958_ (.Y(_1258_),
    .A(net1834),
    .B(net835));
 sg13g2_a21oi_1 _4959_ (.A1(_1257_),
    .A2(_1258_),
    .Y(_0102_),
    .B1(net1038));
 sg13g2_nor2_1 _4960_ (.A(net1904),
    .B(_1255_),
    .Y(_1259_));
 sg13g2_and2_1 _4961_ (.A(\led_controller.cpu.fetch_pc[8] ),
    .B(_1255_),
    .X(_1260_));
 sg13g2_nor3_1 _4962_ (.A(net940),
    .B(_1259_),
    .C(_1260_),
    .Y(_1261_));
 sg13g2_a21oi_1 _4963_ (.A1(net1907),
    .A2(net849),
    .Y(_1262_),
    .B1(_1261_));
 sg13g2_nand2_1 _4964_ (.Y(_1263_),
    .A(net1904),
    .B(net835));
 sg13g2_a21oi_1 _4965_ (.A1(_1262_),
    .A2(_1263_),
    .Y(_0103_),
    .B1(net1027));
 sg13g2_and2_1 _4966_ (.A(\led_controller.cpu.fetch_pc[9] ),
    .B(_1260_),
    .X(_1264_));
 sg13g2_o21ai_1 _4967_ (.B1(net950),
    .Y(_1265_),
    .A1(net1874),
    .A2(_1260_));
 sg13g2_nor2_1 _4968_ (.A(_1264_),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_a21oi_1 _4969_ (.A1(\led_controller.cpu.pc[9] ),
    .A2(net849),
    .Y(_1267_),
    .B1(_1266_));
 sg13g2_nand2_1 _4970_ (.Y(_1268_),
    .A(net1874),
    .B(net834));
 sg13g2_a21oi_1 _4971_ (.A1(_1267_),
    .A2(_1268_),
    .Y(_0104_),
    .B1(net1037));
 sg13g2_o21ai_1 _4972_ (.B1(net950),
    .Y(_1269_),
    .A1(\led_controller.cpu.fetch_pc[10] ),
    .A2(_1264_));
 sg13g2_a21oi_1 _4973_ (.A1(net2267),
    .A2(_1264_),
    .Y(_1270_),
    .B1(_1269_));
 sg13g2_a21o_2 _4974_ (.A2(net849),
    .A1(net2203),
    .B1(_1270_),
    .X(_1271_));
 sg13g2_a22oi_1 _4975_ (.Y(_1272_),
    .B1(_1271_),
    .B2(net1052),
    .A2(net829),
    .A1(net2267));
 sg13g2_inv_1 _4976_ (.Y(_0105_),
    .A(_1272_));
 sg13g2_nand2_1 _4977_ (.Y(_1273_),
    .A(net1838),
    .B(net834));
 sg13g2_and3_1 _4978_ (.X(_1274_),
    .A(net1838),
    .B(\led_controller.cpu.fetch_pc[10] ),
    .C(_1264_));
 sg13g2_a21oi_1 _4979_ (.A1(\led_controller.cpu.fetch_pc[10] ),
    .A2(_1264_),
    .Y(_1275_),
    .B1(net1838));
 sg13g2_nor3_1 _4980_ (.A(net939),
    .B(_1274_),
    .C(_1275_),
    .Y(_1276_));
 sg13g2_a21oi_1 _4981_ (.A1(net2056),
    .A2(net847),
    .Y(_1277_),
    .B1(_1276_));
 sg13g2_a21oi_1 _4982_ (.A1(_1273_),
    .A2(_1277_),
    .Y(_0106_),
    .B1(net1037));
 sg13g2_nand2_1 _4983_ (.Y(_1278_),
    .A(\led_controller.cpu.pc[12] ),
    .B(net847));
 sg13g2_a22oi_1 _4984_ (.Y(_1279_),
    .B1(net834),
    .B2(net2272),
    .A2(net847),
    .A1(net2248));
 sg13g2_and2_1 _4985_ (.A(\led_controller.cpu.fetch_pc[12] ),
    .B(_1274_),
    .X(_1280_));
 sg13g2_nor2_1 _4986_ (.A(net939),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_o21ai_1 _4987_ (.B1(_1281_),
    .Y(_1282_),
    .A1(net2272),
    .A2(_1274_));
 sg13g2_a21oi_1 _4988_ (.A1(_1279_),
    .A2(_1282_),
    .Y(_0107_),
    .B1(net1037));
 sg13g2_o21ai_1 _4989_ (.B1(net950),
    .Y(_1283_),
    .A1(\led_controller.cpu.fetch_pc[13] ),
    .A2(_1280_));
 sg13g2_a21oi_1 _4990_ (.A1(net2224),
    .A2(_1280_),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_a21oi_1 _4991_ (.A1(\led_controller.cpu.pc[13] ),
    .A2(net847),
    .Y(_1285_),
    .B1(_1284_));
 sg13g2_nor2_1 _4992_ (.A(net1037),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_a21o_1 _4993_ (.A2(net829),
    .A1(net2224),
    .B1(_1286_),
    .X(_0108_));
 sg13g2_a21o_1 _4994_ (.A2(_1280_),
    .A1(\led_controller.cpu.fetch_pc[13] ),
    .B1(net1917),
    .X(_1287_));
 sg13g2_nand3_1 _4995_ (.B(\led_controller.cpu.fetch_pc[13] ),
    .C(_1280_),
    .A(net1917),
    .Y(_1288_));
 sg13g2_and2_1 _4996_ (.A(net950),
    .B(_1288_),
    .X(_1289_));
 sg13g2_a22oi_1 _4997_ (.Y(_1290_),
    .B1(_1287_),
    .B2(_1289_),
    .A2(net847),
    .A1(\led_controller.cpu.pc[14] ));
 sg13g2_nand2_1 _4998_ (.Y(_1291_),
    .A(net1917),
    .B(net834));
 sg13g2_a21oi_1 _4999_ (.A1(_1290_),
    .A2(_1291_),
    .Y(_0109_),
    .B1(net1037));
 sg13g2_nor3_1 _5000_ (.A(net2034),
    .B(net939),
    .C(_1288_),
    .Y(_1292_));
 sg13g2_a22oi_1 _5001_ (.Y(_1293_),
    .B1(_1289_),
    .B2(net2034),
    .A2(net847),
    .A1(\led_controller.cpu.pc[15] ));
 sg13g2_nand2b_1 _5002_ (.Y(_1294_),
    .B(_1293_),
    .A_N(_1292_));
 sg13g2_a21oi_1 _5003_ (.A1(net2034),
    .A2(net834),
    .Y(_1295_),
    .B1(_1294_));
 sg13g2_nor2_1 _5004_ (.A(net1027),
    .B(net2035),
    .Y(_0110_));
 sg13g2_nand2_2 _5005_ (.Y(_1296_),
    .A(_1050_),
    .B(_1158_));
 sg13g2_a21oi_2 _5006_ (.B1(net1031),
    .Y(_1297_),
    .A2(_1158_),
    .A1(_1050_));
 sg13g2_nand2_1 _5007_ (.Y(_1298_),
    .A(net779),
    .B(_1297_));
 sg13g2_o21ai_1 _5008_ (.B1(_1298_),
    .Y(_0111_),
    .A1(net934),
    .A2(_1296_));
 sg13g2_nand2_1 _5009_ (.Y(_1299_),
    .A(net815),
    .B(_1297_));
 sg13g2_o21ai_1 _5010_ (.B1(_1299_),
    .Y(_0112_),
    .A1(net931),
    .A2(_1296_));
 sg13g2_nand2_1 _5011_ (.Y(_1300_),
    .A(net770),
    .B(_1297_));
 sg13g2_o21ai_1 _5012_ (.B1(_1300_),
    .Y(_0113_),
    .A1(net929),
    .A2(_1296_));
 sg13g2_nand2_1 _5013_ (.Y(_1301_),
    .A(net776),
    .B(_1297_));
 sg13g2_o21ai_1 _5014_ (.B1(_1301_),
    .Y(_0114_),
    .A1(net926),
    .A2(_1296_));
 sg13g2_nand2_1 _5015_ (.Y(_1302_),
    .A(net766),
    .B(_1297_));
 sg13g2_o21ai_1 _5016_ (.B1(_1302_),
    .Y(_0115_),
    .A1(net925),
    .A2(_1296_));
 sg13g2_nand2_1 _5017_ (.Y(_1303_),
    .A(net769),
    .B(_1297_));
 sg13g2_o21ai_1 _5018_ (.B1(_1303_),
    .Y(_0116_),
    .A1(net921),
    .A2(_1296_));
 sg13g2_nand2_1 _5019_ (.Y(_1304_),
    .A(net791),
    .B(_1297_));
 sg13g2_o21ai_1 _5020_ (.B1(_1304_),
    .Y(_0117_),
    .A1(net919),
    .A2(_1296_));
 sg13g2_nand2_1 _5021_ (.Y(_1305_),
    .A(net771),
    .B(_1297_));
 sg13g2_o21ai_1 _5022_ (.B1(_1305_),
    .Y(_0118_),
    .A1(net917),
    .A2(_1296_));
 sg13g2_nand2_2 _5023_ (.Y(_1306_),
    .A(_1124_),
    .B(_1205_));
 sg13g2_a21oi_2 _5024_ (.B1(net1033),
    .Y(_1307_),
    .A2(_1205_),
    .A1(_1124_));
 sg13g2_nand2_1 _5025_ (.Y(_1308_),
    .A(net816),
    .B(_1307_));
 sg13g2_o21ai_1 _5026_ (.B1(_1308_),
    .Y(_0119_),
    .A1(net936),
    .A2(_1306_));
 sg13g2_nand2_1 _5027_ (.Y(_1309_),
    .A(net1281),
    .B(_1307_));
 sg13g2_o21ai_1 _5028_ (.B1(_1309_),
    .Y(_0120_),
    .A1(net931),
    .A2(_1306_));
 sg13g2_nand2_1 _5029_ (.Y(_1310_),
    .A(net1245),
    .B(_1307_));
 sg13g2_o21ai_1 _5030_ (.B1(_1310_),
    .Y(_0121_),
    .A1(net930),
    .A2(_1306_));
 sg13g2_nand2_1 _5031_ (.Y(_1311_),
    .A(net1237),
    .B(_1307_));
 sg13g2_o21ai_1 _5032_ (.B1(_1311_),
    .Y(_0122_),
    .A1(net928),
    .A2(_1306_));
 sg13g2_nand2_1 _5033_ (.Y(_1312_),
    .A(net810),
    .B(_1307_));
 sg13g2_o21ai_1 _5034_ (.B1(_1312_),
    .Y(_0123_),
    .A1(net924),
    .A2(_1306_));
 sg13g2_nand2_1 _5035_ (.Y(_1313_),
    .A(net1249),
    .B(_1307_));
 sg13g2_o21ai_1 _5036_ (.B1(_1313_),
    .Y(_0124_),
    .A1(net923),
    .A2(_1306_));
 sg13g2_nand2_1 _5037_ (.Y(_1314_),
    .A(net1235),
    .B(_1307_));
 sg13g2_o21ai_1 _5038_ (.B1(_1314_),
    .Y(_0125_),
    .A1(net920),
    .A2(_1306_));
 sg13g2_nand2_1 _5039_ (.Y(_1315_),
    .A(net1279),
    .B(_1307_));
 sg13g2_o21ai_1 _5040_ (.B1(_1315_),
    .Y(_0126_),
    .A1(net916),
    .A2(_1306_));
 sg13g2_nand2b_2 _5041_ (.Y(_1316_),
    .B(net1161),
    .A_N(_0964_));
 sg13g2_nor2_1 _5042_ (.A(net785),
    .B(_1316_),
    .Y(_0127_));
 sg13g2_xnor2_1 _5043_ (.Y(_1317_),
    .A(net785),
    .B(net1872));
 sg13g2_nor2_1 _5044_ (.A(_1316_),
    .B(_1317_),
    .Y(_0128_));
 sg13g2_and3_1 _5045_ (.X(_1318_),
    .A(net785),
    .B(\led_controller.rgbw.counter[1] ),
    .C(net1588));
 sg13g2_a21oi_1 _5046_ (.A1(net785),
    .A2(\led_controller.rgbw.counter[1] ),
    .Y(_1319_),
    .B1(net1588));
 sg13g2_nor3_1 _5047_ (.A(_1316_),
    .B(_1318_),
    .C(net1589),
    .Y(_0129_));
 sg13g2_and2_1 _5048_ (.A(net1723),
    .B(_1318_),
    .X(_1320_));
 sg13g2_nor2_1 _5049_ (.A(net1723),
    .B(_1318_),
    .Y(_1321_));
 sg13g2_nor3_1 _5050_ (.A(_1316_),
    .B(_1320_),
    .C(net1724),
    .Y(_0130_));
 sg13g2_and2_1 _5051_ (.A(net1800),
    .B(_1320_),
    .X(_1322_));
 sg13g2_nor2_1 _5052_ (.A(net1800),
    .B(_1320_),
    .Y(_1323_));
 sg13g2_nor3_1 _5053_ (.A(_1316_),
    .B(_1322_),
    .C(net1801),
    .Y(_0131_));
 sg13g2_and2_1 _5054_ (.A(net1828),
    .B(_1322_),
    .X(_1324_));
 sg13g2_nor2_1 _5055_ (.A(net1828),
    .B(_1322_),
    .Y(_1325_));
 sg13g2_nor3_1 _5056_ (.A(_1316_),
    .B(_1324_),
    .C(_1325_),
    .Y(_0132_));
 sg13g2_nand2_1 _5057_ (.Y(_1326_),
    .A(net1928),
    .B(_1324_));
 sg13g2_xnor2_1 _5058_ (.Y(_1327_),
    .A(net1928),
    .B(_1324_));
 sg13g2_nor2_1 _5059_ (.A(_1316_),
    .B(_1327_),
    .Y(_0133_));
 sg13g2_xor2_1 _5060_ (.B(_1326_),
    .A(net2081),
    .X(_1328_));
 sg13g2_nor2_1 _5061_ (.A(_1316_),
    .B(_1328_),
    .Y(_0134_));
 sg13g2_nand2_1 _5062_ (.Y(_0161_),
    .A(net1150),
    .B(_0891_));
 sg13g2_nand2_1 _5063_ (.Y(_1329_),
    .A(net1470),
    .B(_0891_));
 sg13g2_nor2_1 _5064_ (.A(net1103),
    .B(net1471),
    .Y(_0135_));
 sg13g2_and3_1 _5065_ (.X(_1330_),
    .A(_0891_),
    .B(\led_controller.spi_slave.last_sck ),
    .C(_0892_));
 sg13g2_and2_1 _5066_ (.A(net1145),
    .B(_1330_),
    .X(_1331_));
 sg13g2_inv_1 _5067_ (.Y(_1332_),
    .A(_1331_));
 sg13g2_nand3_1 _5068_ (.B(net1489),
    .C(net1471),
    .A(net1150),
    .Y(_1333_));
 sg13g2_a22oi_1 _5069_ (.Y(_0136_),
    .B1(_1332_),
    .B2(_1333_),
    .A2(_1330_),
    .A1(_0893_));
 sg13g2_nor3_1 _5070_ (.A(\led_controller.spi_slave.ss_n ),
    .B(net1783),
    .C(_0892_),
    .Y(_1334_));
 sg13g2_a21oi_1 _5071_ (.A1(net1470),
    .A2(_0891_),
    .Y(_1335_),
    .B1(net1022));
 sg13g2_inv_1 _5072_ (.Y(_1336_),
    .A(_1335_));
 sg13g2_o21ai_1 _5073_ (.B1(net1150),
    .Y(_1337_),
    .A1(net1494),
    .A2(net1022));
 sg13g2_a21oi_1 _5074_ (.A1(net1494),
    .A2(_1336_),
    .Y(_0137_),
    .B1(_1337_));
 sg13g2_and2_1 _5075_ (.A(\led_controller.spi_slave.data_bits[1] ),
    .B(net1494),
    .X(_1338_));
 sg13g2_xor2_1 _5076_ (.B(net1494),
    .A(net1966),
    .X(_1339_));
 sg13g2_a22oi_1 _5077_ (.Y(_1340_),
    .B1(_1339_),
    .B2(net1022),
    .A2(_1335_),
    .A1(net1966));
 sg13g2_nor2_1 _5078_ (.A(net1110),
    .B(_1340_),
    .Y(_0138_));
 sg13g2_nand2_1 _5079_ (.Y(_1341_),
    .A(net1887),
    .B(_1338_));
 sg13g2_nand2_1 _5080_ (.Y(_1342_),
    .A(net1022),
    .B(_1341_));
 sg13g2_nand2_1 _5081_ (.Y(_1343_),
    .A(net1887),
    .B(_1335_));
 sg13g2_o21ai_1 _5082_ (.B1(net1150),
    .Y(_1344_),
    .A1(net1887),
    .A2(_1338_));
 sg13g2_a21oi_1 _5083_ (.A1(_1342_),
    .A2(net1888),
    .Y(_0139_),
    .B1(_1344_));
 sg13g2_nand3_1 _5084_ (.B(net1022),
    .C(_1338_),
    .A(\led_controller.spi_slave.data_bits[2] ),
    .Y(_1345_));
 sg13g2_nor2_1 _5085_ (.A(_0973_),
    .B(_1336_),
    .Y(_1346_));
 sg13g2_nand2_1 _5086_ (.Y(_1347_),
    .A(net1665),
    .B(_1342_));
 sg13g2_o21ai_1 _5087_ (.B1(net1150),
    .Y(_1348_),
    .A1(_1346_),
    .A2(_1347_));
 sg13g2_a21oi_1 _5088_ (.A1(_0888_),
    .A2(_1345_),
    .Y(_0140_),
    .B1(_1348_));
 sg13g2_a22oi_1 _5089_ (.Y(_1349_),
    .B1(net915),
    .B2(\led_controller.spi_data[0] ),
    .A2(net1021),
    .A1(net1748));
 sg13g2_nor2_1 _5090_ (.A(net1103),
    .B(net1749),
    .Y(_0141_));
 sg13g2_a22oi_1 _5091_ (.Y(_1350_),
    .B1(net915),
    .B2(net1952),
    .A2(net1021),
    .A1(net1994));
 sg13g2_nor2_1 _5092_ (.A(net1103),
    .B(_1350_),
    .Y(_0142_));
 sg13g2_a22oi_1 _5093_ (.Y(_1351_),
    .B1(net915),
    .B2(net1785),
    .A2(net1021),
    .A1(net1952));
 sg13g2_nor2_1 _5094_ (.A(net1103),
    .B(_1351_),
    .Y(_0143_));
 sg13g2_a22oi_1 _5095_ (.Y(_1352_),
    .B1(net915),
    .B2(net1797),
    .A2(net1021),
    .A1(net1785));
 sg13g2_nor2_1 _5096_ (.A(net1103),
    .B(_1352_),
    .Y(_0144_));
 sg13g2_a22oi_1 _5097_ (.Y(_1353_),
    .B1(net915),
    .B2(net1906),
    .A2(net1021),
    .A1(net1797));
 sg13g2_nor2_1 _5098_ (.A(net1103),
    .B(_1353_),
    .Y(_0145_));
 sg13g2_a22oi_1 _5099_ (.Y(_1354_),
    .B1(net915),
    .B2(net1695),
    .A2(net1021),
    .A1(\led_controller.spi_data[4] ));
 sg13g2_nor2_1 _5100_ (.A(net1104),
    .B(net1696),
    .Y(_0146_));
 sg13g2_a22oi_1 _5101_ (.Y(_1355_),
    .B1(net915),
    .B2(net1633),
    .A2(net1021),
    .A1(net1695));
 sg13g2_nor2_1 _5102_ (.A(net1103),
    .B(_1355_),
    .Y(_0147_));
 sg13g2_a22oi_1 _5103_ (.Y(_1356_),
    .B1(net915),
    .B2(net1916),
    .A2(net1021),
    .A1(net1633));
 sg13g2_nor2_1 _5104_ (.A(net1103),
    .B(_1356_),
    .Y(_0148_));
 sg13g2_nand3b_1 _5105_ (.B(net1150),
    .C(_1329_),
    .Y(_1357_),
    .A_N(_1330_));
 sg13g2_nor2b_1 _5106_ (.A(net1142),
    .B_N(net1428),
    .Y(_1358_));
 sg13g2_a21oi_1 _5107_ (.A1(net1498),
    .A2(net1143),
    .Y(_1359_),
    .B1(_1358_));
 sg13g2_nor2_1 _5108_ (.A(_1357_),
    .B(_1359_),
    .Y(_0149_));
 sg13g2_nand2_1 _5109_ (.Y(_1360_),
    .A(net1428),
    .B(_1331_));
 sg13g2_nand2b_1 _5110_ (.Y(_1361_),
    .B(net1142),
    .A_N(\led_controller.spi_data_write[1] ));
 sg13g2_o21ai_1 _5111_ (.B1(_1361_),
    .Y(_1362_),
    .A1(net1142),
    .A2(net1233));
 sg13g2_o21ai_1 _5112_ (.B1(_1360_),
    .Y(_0150_),
    .A1(_1357_),
    .A2(_1362_));
 sg13g2_nand2_1 _5113_ (.Y(_1363_),
    .A(net1233),
    .B(_1331_));
 sg13g2_nand2b_1 _5114_ (.Y(_1364_),
    .B(net1142),
    .A_N(\led_controller.spi_data_write[2] ));
 sg13g2_o21ai_1 _5115_ (.B1(_1364_),
    .Y(_1365_),
    .A1(net1142),
    .A2(\led_controller.spi_slave.output_register[2] ));
 sg13g2_o21ai_1 _5116_ (.B1(_1363_),
    .Y(_0151_),
    .A1(_1357_),
    .A2(_1365_));
 sg13g2_nand2_1 _5117_ (.Y(_1366_),
    .A(net1351),
    .B(_1331_));
 sg13g2_nand2b_1 _5118_ (.Y(_1367_),
    .B(net1142),
    .A_N(\led_controller.spi_data_write[3] ));
 sg13g2_o21ai_1 _5119_ (.B1(_1367_),
    .Y(_1368_),
    .A1(net1142),
    .A2(net1312));
 sg13g2_o21ai_1 _5120_ (.B1(_1366_),
    .Y(_0152_),
    .A1(_1357_),
    .A2(_1368_));
 sg13g2_nand2_1 _5121_ (.Y(_1369_),
    .A(net1312),
    .B(_1331_));
 sg13g2_nand2b_1 _5122_ (.Y(_1370_),
    .B(net1143),
    .A_N(\led_controller.spi_data_write[4] ));
 sg13g2_o21ai_1 _5123_ (.B1(_1370_),
    .Y(_1371_),
    .A1(net1142),
    .A2(net781));
 sg13g2_o21ai_1 _5124_ (.B1(_1369_),
    .Y(_0153_),
    .A1(_1357_),
    .A2(_1371_));
 sg13g2_nand2_1 _5125_ (.Y(_1372_),
    .A(net781),
    .B(_1331_));
 sg13g2_nand2b_1 _5126_ (.Y(_1373_),
    .B(net1143),
    .A_N(\led_controller.spi_data_write[5] ));
 sg13g2_o21ai_1 _5127_ (.B1(_1373_),
    .Y(_1374_),
    .A1(net1143),
    .A2(\led_controller.spi_slave.output_register[5] ));
 sg13g2_o21ai_1 _5128_ (.B1(_1372_),
    .Y(_0154_),
    .A1(_1357_),
    .A2(_1374_));
 sg13g2_nand2_1 _5129_ (.Y(_1375_),
    .A(net1393),
    .B(_1331_));
 sg13g2_nand2b_1 _5130_ (.Y(_1376_),
    .B(net1143),
    .A_N(\led_controller.spi_data_write[6] ));
 sg13g2_o21ai_1 _5131_ (.B1(_1376_),
    .Y(_1377_),
    .A1(net1143),
    .A2(net1335));
 sg13g2_o21ai_1 _5132_ (.B1(_1375_),
    .Y(_0155_),
    .A1(_1357_),
    .A2(_1377_));
 sg13g2_nand2_1 _5133_ (.Y(_1378_),
    .A(net1335),
    .B(_1331_));
 sg13g2_nand2b_1 _5134_ (.Y(_1379_),
    .B(net1143),
    .A_N(\led_controller.spi_data_write[7] ));
 sg13g2_o21ai_1 _5135_ (.B1(_1379_),
    .Y(_1380_),
    .A1(\led_controller.spi_data_write_strb ),
    .A2(\led_controller.spi_slave.output_register[7] ));
 sg13g2_o21ai_1 _5136_ (.B1(_1378_),
    .Y(_0156_),
    .A1(_1357_),
    .A2(_1380_));
 sg13g2_nor2_1 _5137_ (.A(net1110),
    .B(_0892_),
    .Y(_0157_));
 sg13g2_and2_1 _5138_ (.A(net1152),
    .B(net763),
    .X(_0158_));
 sg13g2_and2_1 _5139_ (.A(net1152),
    .B(net4),
    .X(_0159_));
 sg13g2_and2_1 _5140_ (.A(net1151),
    .B(net762),
    .X(_0160_));
 sg13g2_and2_1 _5141_ (.A(net1153),
    .B(net761),
    .X(_0162_));
 sg13g2_and2_1 _5142_ (.A(net1154),
    .B(net2),
    .X(_0163_));
 sg13g2_nor4_1 _5143_ (.A(\led_controller.timer_2hz.counter[3] ),
    .B(\led_controller.timer_2hz.counter[2] ),
    .C(_0881_),
    .D(\led_controller.timer_2hz.counter[0] ),
    .Y(_1381_));
 sg13g2_nand3_1 _5144_ (.B(\led_controller.timer_2hz.counter[4] ),
    .C(_1381_),
    .A(\led_controller.timer_2hz.counter[5] ),
    .Y(_1382_));
 sg13g2_nand2_2 _5145_ (.Y(_1383_),
    .A(net1158),
    .B(_1382_));
 sg13g2_xnor2_1 _5146_ (.Y(_1384_),
    .A(\led_controller.cpu.i_timer_100hz ),
    .B(net1713));
 sg13g2_nor2_1 _5147_ (.A(_1383_),
    .B(net1714),
    .Y(_0164_));
 sg13g2_and3_1 _5148_ (.X(_1385_),
    .A(\led_controller.cpu.i_timer_100hz ),
    .B(net1405),
    .C(\led_controller.timer_2hz.counter[0] ));
 sg13g2_a21oi_1 _5149_ (.A1(\led_controller.cpu.i_timer_100hz ),
    .A2(\led_controller.timer_2hz.counter[0] ),
    .Y(_1386_),
    .B1(net1405));
 sg13g2_nor3_1 _5150_ (.A(_1383_),
    .B(_1385_),
    .C(net1406),
    .Y(_0165_));
 sg13g2_and2_1 _5151_ (.A(net1630),
    .B(_1385_),
    .X(_1387_));
 sg13g2_nor2_1 _5152_ (.A(net1630),
    .B(_1385_),
    .Y(_1388_));
 sg13g2_nor3_1 _5153_ (.A(_1383_),
    .B(_1387_),
    .C(net1631),
    .Y(_0166_));
 sg13g2_nor2_1 _5154_ (.A(net1675),
    .B(_1387_),
    .Y(_1389_));
 sg13g2_and2_1 _5155_ (.A(net1675),
    .B(_1387_),
    .X(_1390_));
 sg13g2_nor3_1 _5156_ (.A(_1383_),
    .B(net1676),
    .C(_1390_),
    .Y(_0167_));
 sg13g2_nor2_1 _5157_ (.A(net1790),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_and2_1 _5158_ (.A(net1790),
    .B(_1390_),
    .X(_1392_));
 sg13g2_nor3_1 _5159_ (.A(_1383_),
    .B(_1391_),
    .C(_1392_),
    .Y(_0168_));
 sg13g2_a21oi_1 _5160_ (.A1(net2094),
    .A2(_1392_),
    .Y(_1393_),
    .B1(_1383_));
 sg13g2_o21ai_1 _5161_ (.B1(_1393_),
    .Y(_1394_),
    .A1(net2094),
    .A2(_1392_));
 sg13g2_inv_1 _5162_ (.Y(_0169_),
    .A(_1394_));
 sg13g2_nand2b_2 _5163_ (.Y(_1395_),
    .B(net1158),
    .A_N(_1012_));
 sg13g2_nor2_1 _5164_ (.A(\led_controller.cpu.i_timer_100hz ),
    .B(net1697),
    .Y(_1396_));
 sg13g2_and2_1 _5165_ (.A(\led_controller.cpu.i_timer_100hz ),
    .B(net1697),
    .X(_1397_));
 sg13g2_nor3_1 _5166_ (.A(_1395_),
    .B(net1698),
    .C(_1397_),
    .Y(_0170_));
 sg13g2_xnor2_1 _5167_ (.Y(_1398_),
    .A(net1961),
    .B(_1397_));
 sg13g2_nor2_1 _5168_ (.A(_1395_),
    .B(net1962),
    .Y(_0171_));
 sg13g2_a21oi_1 _5169_ (.A1(\led_controller.timer_10hz.counter[1] ),
    .A2(_1397_),
    .Y(_1399_),
    .B1(net1558));
 sg13g2_nand3_1 _5170_ (.B(net1961),
    .C(_1397_),
    .A(net1558),
    .Y(_1400_));
 sg13g2_inv_1 _5171_ (.Y(_1401_),
    .A(_1400_));
 sg13g2_nor3_1 _5172_ (.A(_1395_),
    .B(net1559),
    .C(_1401_),
    .Y(_0172_));
 sg13g2_xor2_1 _5173_ (.B(_1400_),
    .A(net1982),
    .X(_1402_));
 sg13g2_nor2_1 _5174_ (.A(_1395_),
    .B(_1402_),
    .Y(_0173_));
 sg13g2_nor2_1 _5175_ (.A(net1111),
    .B(uio_oe[0]),
    .Y(_0174_));
 sg13g2_nand2_1 _5176_ (.Y(_1403_),
    .A(net2159),
    .B(_1181_));
 sg13g2_inv_1 _5177_ (.Y(_1404_),
    .A(_1403_));
 sg13g2_nor4_1 _5178_ (.A(net2307),
    .B(net2200),
    .C(net1770),
    .D(net2159),
    .Y(_1405_));
 sg13g2_nor2_1 _5179_ (.A(net2104),
    .B(net2328),
    .Y(_1406_));
 sg13g2_nand4_1 _5180_ (.B(net2063),
    .C(_1405_),
    .A(net2169),
    .Y(_1407_),
    .D(_1406_));
 sg13g2_nor2_1 _5181_ (.A(net2119),
    .B(net2023),
    .Y(_1408_));
 sg13g2_nor4_1 _5182_ (.A(net2242),
    .B(net1964),
    .C(net1895),
    .D(net2177),
    .Y(_1409_));
 sg13g2_nand4_1 _5183_ (.B(net1455),
    .C(_1408_),
    .A(net1595),
    .Y(_1410_),
    .D(_1409_));
 sg13g2_nor4_1 _5184_ (.A(net2072),
    .B(net1811),
    .C(net2222),
    .D(net2174),
    .Y(_1411_));
 sg13g2_nand2_1 _5185_ (.Y(_1412_),
    .A(net1933),
    .B(net2197));
 sg13g2_nor3_1 _5186_ (.A(net1546),
    .B(net1306),
    .C(_1412_),
    .Y(_1413_));
 sg13g2_nor4_1 _5187_ (.A(net2275),
    .B(\led_controller.timer_100hz.counter[20] ),
    .C(net1900),
    .D(net2182),
    .Y(_1414_));
 sg13g2_nor4_1 _5188_ (.A(net2324),
    .B(net2234),
    .C(net2258),
    .D(net1958),
    .Y(_1415_));
 sg13g2_nand4_1 _5189_ (.B(_1413_),
    .C(_1414_),
    .A(_1411_),
    .Y(_1416_),
    .D(_1415_));
 sg13g2_nor3_1 _5190_ (.A(_1407_),
    .B(_1410_),
    .C(_1416_),
    .Y(_1417_));
 sg13g2_nand2b_1 _5191_ (.Y(_1418_),
    .B(net1158),
    .A_N(_1417_));
 sg13g2_inv_1 _5192_ (.Y(_1419_),
    .A(net914));
 sg13g2_o21ai_1 _5193_ (.B1(net873),
    .Y(_1420_),
    .A1(net2159),
    .A2(_1181_));
 sg13g2_nor2_1 _5194_ (.A(_1404_),
    .B(net2160),
    .Y(_0175_));
 sg13g2_nor2_1 _5195_ (.A(net1770),
    .B(_1404_),
    .Y(_1421_));
 sg13g2_and3_2 _5196_ (.X(_1422_),
    .A(net1770),
    .B(net2159),
    .C(_1181_));
 sg13g2_nor3_1 _5197_ (.A(net914),
    .B(net1771),
    .C(_1422_),
    .Y(_0176_));
 sg13g2_a21oi_1 _5198_ (.A1(net2200),
    .A2(_1422_),
    .Y(_1423_),
    .B1(net914));
 sg13g2_o21ai_1 _5199_ (.B1(_1423_),
    .Y(_1424_),
    .A1(net2200),
    .A2(_1422_));
 sg13g2_inv_1 _5200_ (.Y(_0177_),
    .A(_1424_));
 sg13g2_a21o_1 _5201_ (.A2(_1422_),
    .A1(net2200),
    .B1(net2307),
    .X(_1425_));
 sg13g2_nand3_1 _5202_ (.B(net2200),
    .C(_1422_),
    .A(net2307),
    .Y(_1426_));
 sg13g2_and3_1 _5203_ (.X(_0178_),
    .A(net872),
    .B(_1425_),
    .C(_1426_));
 sg13g2_nor2_1 _5204_ (.A(_0880_),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_a21oi_1 _5205_ (.A1(_0880_),
    .A2(_1426_),
    .Y(_1428_),
    .B1(net914));
 sg13g2_nor2b_1 _5206_ (.A(_1427_),
    .B_N(_1428_),
    .Y(_0179_));
 sg13g2_nor3_1 _5207_ (.A(_0879_),
    .B(_0880_),
    .C(_1426_),
    .Y(_1429_));
 sg13g2_o21ai_1 _5208_ (.B1(net872),
    .Y(_1430_),
    .A1(net2063),
    .A2(_1427_));
 sg13g2_nor2_1 _5209_ (.A(_1429_),
    .B(net2064),
    .Y(_0180_));
 sg13g2_nor4_1 _5210_ (.A(_0878_),
    .B(_0879_),
    .C(_0880_),
    .D(_1426_),
    .Y(_1431_));
 sg13g2_o21ai_1 _5211_ (.B1(net872),
    .Y(_1432_),
    .A1(net2104),
    .A2(_1429_));
 sg13g2_nor2_1 _5212_ (.A(_1431_),
    .B(net2105),
    .Y(_0181_));
 sg13g2_and2_1 _5213_ (.A(net2169),
    .B(_1431_),
    .X(_1433_));
 sg13g2_o21ai_1 _5214_ (.B1(net872),
    .Y(_1434_),
    .A1(net2169),
    .A2(_1431_));
 sg13g2_nor2_1 _5215_ (.A(_1433_),
    .B(net2170),
    .Y(_0182_));
 sg13g2_and3_2 _5216_ (.X(_1435_),
    .A(net2023),
    .B(net2386),
    .C(_1431_));
 sg13g2_o21ai_1 _5217_ (.B1(net872),
    .Y(_1436_),
    .A1(net2023),
    .A2(_1433_));
 sg13g2_nor2_1 _5218_ (.A(_1435_),
    .B(net2024),
    .Y(_0183_));
 sg13g2_o21ai_1 _5219_ (.B1(net872),
    .Y(_1437_),
    .A1(net1455),
    .A2(_1435_));
 sg13g2_a21oi_1 _5220_ (.A1(net1455),
    .A2(_1435_),
    .Y(_0184_),
    .B1(_1437_));
 sg13g2_a21oi_1 _5221_ (.A1(net1455),
    .A2(_1435_),
    .Y(_1438_),
    .B1(net1595));
 sg13g2_and3_1 _5222_ (.X(_1439_),
    .A(net1595),
    .B(net1455),
    .C(_1435_));
 sg13g2_nor3_1 _5223_ (.A(net914),
    .B(net1596),
    .C(_1439_),
    .Y(_0185_));
 sg13g2_and4_1 _5224_ (.A(net2119),
    .B(net1595),
    .C(net1455),
    .D(_1435_),
    .X(_1440_));
 sg13g2_o21ai_1 _5225_ (.B1(net872),
    .Y(_1441_),
    .A1(net2119),
    .A2(_1439_));
 sg13g2_nor2_1 _5226_ (.A(_1440_),
    .B(_1441_),
    .Y(_0186_));
 sg13g2_and2_1 _5227_ (.A(net2177),
    .B(_1440_),
    .X(_1442_));
 sg13g2_o21ai_1 _5228_ (.B1(net872),
    .Y(_1443_),
    .A1(net2177),
    .A2(_1440_));
 sg13g2_nor2_1 _5229_ (.A(_1442_),
    .B(_1443_),
    .Y(_0187_));
 sg13g2_nor2_1 _5230_ (.A(net1895),
    .B(_1442_),
    .Y(_1444_));
 sg13g2_and4_1 _5231_ (.A(net1895),
    .B(net2384),
    .C(\led_controller.timer_100hz.counter[11] ),
    .D(_1439_),
    .X(_1445_));
 sg13g2_nor3_1 _5232_ (.A(net914),
    .B(net1896),
    .C(_1445_),
    .Y(_0188_));
 sg13g2_nor2_1 _5233_ (.A(net1964),
    .B(_1445_),
    .Y(_1446_));
 sg13g2_and2_1 _5234_ (.A(net1964),
    .B(net2385),
    .X(_1447_));
 sg13g2_nor3_1 _5235_ (.A(net913),
    .B(net1965),
    .C(_1447_),
    .Y(_0189_));
 sg13g2_and4_1 _5236_ (.A(net2197),
    .B(net1964),
    .C(net1895),
    .D(_1442_),
    .X(_1448_));
 sg13g2_o21ai_1 _5237_ (.B1(net871),
    .Y(_1449_),
    .A1(net2197),
    .A2(_1447_));
 sg13g2_nor2_1 _5238_ (.A(_1448_),
    .B(net2198),
    .Y(_0190_));
 sg13g2_nor2_1 _5239_ (.A(net1933),
    .B(_1448_),
    .Y(_1450_));
 sg13g2_and3_1 _5240_ (.X(_1451_),
    .A(net1933),
    .B(net2197),
    .C(_1447_));
 sg13g2_nor3_1 _5241_ (.A(net913),
    .B(net1934),
    .C(_1451_),
    .Y(_0191_));
 sg13g2_and3_1 _5242_ (.X(_1452_),
    .A(net2242),
    .B(net1933),
    .C(_1448_));
 sg13g2_o21ai_1 _5243_ (.B1(net871),
    .Y(_1453_),
    .A1(net2242),
    .A2(_1451_));
 sg13g2_nor2_1 _5244_ (.A(_1452_),
    .B(_1453_),
    .Y(_0192_));
 sg13g2_and2_1 _5245_ (.A(net2182),
    .B(_1452_),
    .X(_1454_));
 sg13g2_o21ai_1 _5246_ (.B1(net873),
    .Y(_1455_),
    .A1(net2182),
    .A2(_1452_));
 sg13g2_nor2_1 _5247_ (.A(_1454_),
    .B(net2183),
    .Y(_0193_));
 sg13g2_nor2_1 _5248_ (.A(net1900),
    .B(_1454_),
    .Y(_1456_));
 sg13g2_and4_1 _5249_ (.A(net1900),
    .B(net2182),
    .C(net2242),
    .D(_1451_),
    .X(_1457_));
 sg13g2_nor3_1 _5250_ (.A(net914),
    .B(net1901),
    .C(_1457_),
    .Y(_0194_));
 sg13g2_or2_1 _5251_ (.X(_1458_),
    .B(_1457_),
    .A(net2346));
 sg13g2_nand2_1 _5252_ (.Y(_1459_),
    .A(net2346),
    .B(_1457_));
 sg13g2_and3_1 _5253_ (.X(_0195_),
    .A(net871),
    .B(_1458_),
    .C(_1459_));
 sg13g2_and4_1 _5254_ (.A(\led_controller.timer_100hz.counter[21] ),
    .B(\led_controller.timer_100hz.counter[20] ),
    .C(net1900),
    .D(_1454_),
    .X(_1460_));
 sg13g2_xnor2_1 _5255_ (.Y(_1461_),
    .A(net2275),
    .B(_1459_));
 sg13g2_nand2_1 _5256_ (.Y(_1462_),
    .A(net871),
    .B(net2276));
 sg13g2_inv_1 _5257_ (.Y(_0196_),
    .A(_1462_));
 sg13g2_nor2_1 _5258_ (.A(net1958),
    .B(_1460_),
    .Y(_1463_));
 sg13g2_and4_1 _5259_ (.A(net1958),
    .B(net2275),
    .C(net2347),
    .D(_1457_),
    .X(_1464_));
 sg13g2_nor3_1 _5260_ (.A(net913),
    .B(net1959),
    .C(_1464_),
    .Y(_0197_));
 sg13g2_and3_1 _5261_ (.X(_1465_),
    .A(net2258),
    .B(net1958),
    .C(_1460_));
 sg13g2_o21ai_1 _5262_ (.B1(net871),
    .Y(_1466_),
    .A1(net2258),
    .A2(_1464_));
 sg13g2_nor2_1 _5263_ (.A(_1465_),
    .B(net2259),
    .Y(_0198_));
 sg13g2_nand3_1 _5264_ (.B(net2258),
    .C(_1464_),
    .A(net2234),
    .Y(_1467_));
 sg13g2_o21ai_1 _5265_ (.B1(_1467_),
    .Y(_1468_),
    .A1(net2234),
    .A2(_1465_));
 sg13g2_nor2_1 _5266_ (.A(net913),
    .B(net2235),
    .Y(_0199_));
 sg13g2_and2_1 _5267_ (.A(_0877_),
    .B(_1467_),
    .X(_1469_));
 sg13g2_nor2_1 _5268_ (.A(_0877_),
    .B(_1467_),
    .Y(_1470_));
 sg13g2_nor3_1 _5269_ (.A(net913),
    .B(_1469_),
    .C(_1470_),
    .Y(_0200_));
 sg13g2_and4_1 _5270_ (.A(net2174),
    .B(\led_controller.timer_100hz.counter[25] ),
    .C(\led_controller.timer_100hz.counter[24] ),
    .D(_1465_),
    .X(_1471_));
 sg13g2_o21ai_1 _5271_ (.B1(net871),
    .Y(_1472_),
    .A1(net2174),
    .A2(_1470_));
 sg13g2_nor2_1 _5272_ (.A(_1471_),
    .B(net2175),
    .Y(_0201_));
 sg13g2_nand3_1 _5273_ (.B(net2174),
    .C(_1470_),
    .A(net2222),
    .Y(_1473_));
 sg13g2_o21ai_1 _5274_ (.B1(_1473_),
    .Y(_1474_),
    .A1(net2222),
    .A2(_1471_));
 sg13g2_nor2_1 _5275_ (.A(net913),
    .B(net2223),
    .Y(_0202_));
 sg13g2_nor2b_1 _5276_ (.A(net1811),
    .B_N(_1473_),
    .Y(_1475_));
 sg13g2_and3_1 _5277_ (.X(_1476_),
    .A(net1811),
    .B(\led_controller.timer_100hz.counter[27] ),
    .C(_1471_));
 sg13g2_nor3_1 _5278_ (.A(net913),
    .B(net1812),
    .C(_1476_),
    .Y(_0203_));
 sg13g2_and4_1 _5279_ (.A(net2072),
    .B(net1811),
    .C(\led_controller.timer_100hz.counter[27] ),
    .D(_1471_),
    .X(_1477_));
 sg13g2_o21ai_1 _5280_ (.B1(net871),
    .Y(_1478_),
    .A1(net2072),
    .A2(_1476_));
 sg13g2_nor2_1 _5281_ (.A(_1477_),
    .B(net2073),
    .Y(_0204_));
 sg13g2_o21ai_1 _5282_ (.B1(net871),
    .Y(_1479_),
    .A1(net1306),
    .A2(_1477_));
 sg13g2_a21oi_1 _5283_ (.A1(net1306),
    .A2(_1477_),
    .Y(_0205_),
    .B1(_1479_));
 sg13g2_a21oi_1 _5284_ (.A1(net1306),
    .A2(_1477_),
    .Y(_1480_),
    .B1(net1546));
 sg13g2_and3_1 _5285_ (.X(_1481_),
    .A(net1546),
    .B(net1306),
    .C(_1477_));
 sg13g2_nor3_1 _5286_ (.A(net913),
    .B(net1547),
    .C(_1481_),
    .Y(_0206_));
 sg13g2_and2_1 _5287_ (.A(net1158),
    .B(net2329),
    .X(_0207_));
 sg13g2_nand2_2 _5288_ (.Y(_1482_),
    .A(_1050_),
    .B(_1205_));
 sg13g2_a21oi_2 _5289_ (.B1(net1032),
    .Y(_1483_),
    .A2(_1205_),
    .A1(_1050_));
 sg13g2_nand2_1 _5290_ (.Y(_1484_),
    .A(net1350),
    .B(_1483_));
 sg13g2_o21ai_1 _5291_ (.B1(_1484_),
    .Y(_0208_),
    .A1(net936),
    .A2(_1482_));
 sg13g2_nand2_1 _5292_ (.Y(_1485_),
    .A(net1276),
    .B(_1483_));
 sg13g2_o21ai_1 _5293_ (.B1(_1485_),
    .Y(_0209_),
    .A1(net931),
    .A2(_1482_));
 sg13g2_nand2_1 _5294_ (.Y(_1486_),
    .A(net1363),
    .B(_1483_));
 sg13g2_o21ai_1 _5295_ (.B1(_1486_),
    .Y(_0210_),
    .A1(net930),
    .A2(_1482_));
 sg13g2_nand2_1 _5296_ (.Y(_1487_),
    .A(net1248),
    .B(_1483_));
 sg13g2_o21ai_1 _5297_ (.B1(_1487_),
    .Y(_0211_),
    .A1(net928),
    .A2(_1482_));
 sg13g2_nand2_1 _5298_ (.Y(_1488_),
    .A(net1230),
    .B(_1483_));
 sg13g2_o21ai_1 _5299_ (.B1(_1488_),
    .Y(_0212_),
    .A1(net924),
    .A2(_1482_));
 sg13g2_nand2_1 _5300_ (.Y(_1489_),
    .A(net772),
    .B(_1483_));
 sg13g2_o21ai_1 _5301_ (.B1(_1489_),
    .Y(_0213_),
    .A1(net923),
    .A2(_1482_));
 sg13g2_nand2_1 _5302_ (.Y(_1490_),
    .A(net792),
    .B(_1483_));
 sg13g2_o21ai_1 _5303_ (.B1(_1490_),
    .Y(_0214_),
    .A1(net920),
    .A2(_1482_));
 sg13g2_nand2_1 _5304_ (.Y(_1491_),
    .A(net1309),
    .B(_1483_));
 sg13g2_o21ai_1 _5305_ (.B1(_1491_),
    .Y(_0215_),
    .A1(net916),
    .A2(_1482_));
 sg13g2_nand2_1 _5306_ (.Y(_1492_),
    .A(net1191),
    .B(_0964_));
 sg13g2_a21oi_1 _5307_ (.A1(net1191),
    .A2(_0964_),
    .Y(_1493_),
    .B1(net1408));
 sg13g2_nor3_1 _5308_ (.A(net2109),
    .B(net2188),
    .C(\led_controller.rgbw.high_cycles[0] ),
    .Y(_1494_));
 sg13g2_nor2b_1 _5309_ (.A(_1492_),
    .B_N(_1494_),
    .Y(_1495_));
 sg13g2_nor2b_2 _5310_ (.A(net1191),
    .B_N(\led_controller.rgbw.state[1] ),
    .Y(_1496_));
 sg13g2_nand2_1 _5311_ (.Y(_1497_),
    .A(_0883_),
    .B(\led_controller.rgbw.state[1] ));
 sg13g2_nor4_1 _5312_ (.A(net1111),
    .B(net1409),
    .C(_1495_),
    .D(_1496_),
    .Y(_0216_));
 sg13g2_nor2_1 _5313_ (.A(net1098),
    .B(_0964_),
    .Y(_1498_));
 sg13g2_o21ai_1 _5314_ (.B1(net856),
    .Y(_1499_),
    .A1(\led_controller.rgbw.state[1] ),
    .A2(net1098));
 sg13g2_nor2b_1 _5315_ (.A(_1498_),
    .B_N(_1499_),
    .Y(_1500_));
 sg13g2_nand3_1 _5316_ (.B(_0933_),
    .C(_0964_),
    .A(net1191),
    .Y(_1501_));
 sg13g2_and3_2 _5317_ (.X(_1502_),
    .A(net2353),
    .B(_1500_),
    .C(_1501_));
 sg13g2_a21oi_2 _5318_ (.B1(_1502_),
    .Y(_1503_),
    .A2(_0938_),
    .A1(net2373));
 sg13g2_inv_1 _5319_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_o21ai_1 _5320_ (.B1(net1156),
    .Y(_1505_),
    .A1(net1190),
    .A2(_1502_));
 sg13g2_a21oi_1 _5321_ (.A1(net1190),
    .A2(_1504_),
    .Y(_0217_),
    .B1(_1505_));
 sg13g2_and2_1 _5322_ (.A(net1189),
    .B(net1190),
    .X(_1506_));
 sg13g2_or2_1 _5323_ (.X(_1507_),
    .B(net1097),
    .A(_0965_));
 sg13g2_a22oi_1 _5324_ (.Y(_1508_),
    .B1(_1507_),
    .B2(_1502_),
    .A2(_1503_),
    .A1(net1189));
 sg13g2_nor2_1 _5325_ (.A(net1125),
    .B(_1508_),
    .Y(_0218_));
 sg13g2_xor2_1 _5326_ (.B(_0965_),
    .A(net2204),
    .X(_1509_));
 sg13g2_a22oi_1 _5327_ (.Y(_1510_),
    .B1(_1509_),
    .B2(_1502_),
    .A2(_1503_),
    .A1(net2204));
 sg13g2_nor2_1 _5328_ (.A(net1125),
    .B(net2205),
    .Y(_0219_));
 sg13g2_xnor2_1 _5329_ (.Y(_1511_),
    .A(\led_controller.rgbw.pixel_counter[3] ),
    .B(_0966_));
 sg13g2_inv_2 _5330_ (.Y(_1512_),
    .A(net1020));
 sg13g2_a22oi_1 _5331_ (.Y(_1513_),
    .B1(_1512_),
    .B2(_1502_),
    .A2(_1503_),
    .A1(net1978));
 sg13g2_nor2_1 _5332_ (.A(net1114),
    .B(net1979),
    .Y(_0220_));
 sg13g2_xnor2_1 _5333_ (.Y(_1514_),
    .A(\led_controller.rgbw.pixel_counter[4] ),
    .B(_0967_));
 sg13g2_xnor2_1 _5334_ (.Y(_1515_),
    .A(_0876_),
    .B(_0967_));
 sg13g2_a22oi_1 _5335_ (.Y(_1516_),
    .B1(_1515_),
    .B2(_1502_),
    .A2(_1503_),
    .A1(net2213));
 sg13g2_nor2_1 _5336_ (.A(net1114),
    .B(net2214),
    .Y(_0221_));
 sg13g2_a21oi_1 _5337_ (.A1(_0876_),
    .A2(_0967_),
    .Y(_1517_),
    .B1(_0875_));
 sg13g2_nor2_1 _5338_ (.A(_0968_),
    .B(_1517_),
    .Y(_1518_));
 sg13g2_a221oi_1 _5339_ (.B2(_1502_),
    .C1(net1115),
    .B1(_1518_),
    .A1(_0875_),
    .Y(_0222_),
    .A2(_1503_));
 sg13g2_nand2_1 _5340_ (.Y(_1519_),
    .A(net1165),
    .B(net1163));
 sg13g2_and3_2 _5341_ (.X(_1520_),
    .A(net1165),
    .B(net1187),
    .C(net1163));
 sg13g2_nor2_2 _5342_ (.A(net2228),
    .B(net1187),
    .Y(_1521_));
 sg13g2_nor3_1 _5343_ (.A(net1130),
    .B(net1096),
    .C(_1521_),
    .Y(_0223_));
 sg13g2_nand2_1 _5344_ (.Y(_1522_),
    .A(\led_controller.effect_chase_led_color[1] ),
    .B(_0934_));
 sg13g2_o21ai_1 _5345_ (.B1(_1522_),
    .Y(_1523_),
    .A1(_0871_),
    .A2(_0934_));
 sg13g2_nand2_1 _5346_ (.Y(_1524_),
    .A(\led_controller.effect_chase_led_color[0] ),
    .B(_0934_));
 sg13g2_o21ai_1 _5347_ (.B1(_1524_),
    .Y(_1525_),
    .A1(_0872_),
    .A2(_0934_));
 sg13g2_nor2b_2 _5348_ (.A(_1523_),
    .B_N(_1525_),
    .Y(_1526_));
 sg13g2_a21oi_1 _5349_ (.A1(\led_controller.colors[32] ),
    .A2(net912),
    .Y(_1527_),
    .B1(net996));
 sg13g2_nor2_1 _5350_ (.A(_1523_),
    .B(_1525_),
    .Y(_1528_));
 sg13g2_nor2b_1 _5351_ (.A(_1525_),
    .B_N(_1523_),
    .Y(_1529_));
 sg13g2_a22oi_1 _5352_ (.Y(_1530_),
    .B1(net900),
    .B2(\led_controller.colors[0] ),
    .A2(net906),
    .A1(\led_controller.colors[64] ));
 sg13g2_nand2_1 _5353_ (.Y(_1531_),
    .A(_1527_),
    .B(_1530_));
 sg13g2_a21oi_1 _5354_ (.A1(_0793_),
    .A2(net997),
    .Y(_1532_),
    .B1(net862));
 sg13g2_a22oi_1 _5355_ (.Y(_1533_),
    .B1(_1531_),
    .B2(_1532_),
    .A2(net862),
    .A1(net1669));
 sg13g2_nor2_1 _5356_ (.A(net1129),
    .B(net1670),
    .Y(_0224_));
 sg13g2_a21oi_1 _5357_ (.A1(\led_controller.colors[33] ),
    .A2(net911),
    .Y(_1534_),
    .B1(net995));
 sg13g2_a22oi_1 _5358_ (.Y(_1535_),
    .B1(net899),
    .B2(\led_controller.colors[1] ),
    .A2(net905),
    .A1(\led_controller.colors[65] ));
 sg13g2_nand2_1 _5359_ (.Y(_1536_),
    .A(_1534_),
    .B(_1535_));
 sg13g2_a21oi_1 _5360_ (.A1(_0792_),
    .A2(net999),
    .Y(_1537_),
    .B1(net862));
 sg13g2_a22oi_1 _5361_ (.Y(_1538_),
    .B1(_1536_),
    .B2(_1537_),
    .A2(net862),
    .A1(net1649));
 sg13g2_nor2_1 _5362_ (.A(net1128),
    .B(net1650),
    .Y(_0225_));
 sg13g2_a21oi_1 _5363_ (.A1(\led_controller.colors[34] ),
    .A2(net910),
    .Y(_1539_),
    .B1(net993));
 sg13g2_a22oi_1 _5364_ (.Y(_1540_),
    .B1(net898),
    .B2(\led_controller.colors[2] ),
    .A2(net904),
    .A1(net1693));
 sg13g2_nand2_1 _5365_ (.Y(_1541_),
    .A(_1539_),
    .B(_1540_));
 sg13g2_a21oi_1 _5366_ (.A1(_0791_),
    .A2(net994),
    .Y(_1542_),
    .B1(net858));
 sg13g2_a22oi_1 _5367_ (.Y(_1543_),
    .B1(_1541_),
    .B2(_1542_),
    .A2(net858),
    .A1(net1912));
 sg13g2_nor2_1 _5368_ (.A(net1121),
    .B(net1913),
    .Y(_0226_));
 sg13g2_a21oi_1 _5369_ (.A1(\led_controller.colors[35] ),
    .A2(net910),
    .Y(_1544_),
    .B1(net995));
 sg13g2_a22oi_1 _5370_ (.Y(_1545_),
    .B1(net898),
    .B2(\led_controller.colors[3] ),
    .A2(net904),
    .A1(net1885));
 sg13g2_nand2_1 _5371_ (.Y(_1546_),
    .A(_1544_),
    .B(_1545_));
 sg13g2_a21oi_1 _5372_ (.A1(_0790_),
    .A2(net994),
    .Y(_1547_),
    .B1(net858));
 sg13g2_a22oi_1 _5373_ (.Y(_1548_),
    .B1(_1546_),
    .B2(_1547_),
    .A2(net858),
    .A1(net1991));
 sg13g2_nor2_1 _5374_ (.A(net1121),
    .B(net1992),
    .Y(_0227_));
 sg13g2_a21oi_1 _5375_ (.A1(\led_controller.colors[36] ),
    .A2(net912),
    .Y(_1549_),
    .B1(net993));
 sg13g2_a22oi_1 _5376_ (.Y(_1550_),
    .B1(net899),
    .B2(\led_controller.colors[4] ),
    .A2(net905),
    .A1(\led_controller.colors[68] ));
 sg13g2_nand2_1 _5377_ (.Y(_1551_),
    .A(_1549_),
    .B(_1550_));
 sg13g2_a21oi_1 _5378_ (.A1(_0789_),
    .A2(net997),
    .Y(_1552_),
    .B1(net864));
 sg13g2_a22oi_1 _5379_ (.Y(_1553_),
    .B1(_1551_),
    .B2(_1552_),
    .A2(net860),
    .A1(net1791));
 sg13g2_nor2_1 _5380_ (.A(net1125),
    .B(net1792),
    .Y(_0228_));
 sg13g2_a21oi_1 _5381_ (.A1(\led_controller.colors[37] ),
    .A2(_1526_),
    .Y(_1554_),
    .B1(net993));
 sg13g2_a22oi_1 _5382_ (.Y(_1555_),
    .B1(net901),
    .B2(\led_controller.colors[5] ),
    .A2(net907),
    .A1(\led_controller.colors[69] ));
 sg13g2_nand2_1 _5383_ (.Y(_1556_),
    .A(_1554_),
    .B(_1555_));
 sg13g2_a21oi_1 _5384_ (.A1(_0788_),
    .A2(net998),
    .Y(_1557_),
    .B1(net864));
 sg13g2_a22oi_1 _5385_ (.Y(_1558_),
    .B1(_1556_),
    .B2(_1557_),
    .A2(net856),
    .A1(net1686));
 sg13g2_nor2_1 _5386_ (.A(net1114),
    .B(net1687),
    .Y(_0229_));
 sg13g2_a21oi_1 _5387_ (.A1(\led_controller.colors[38] ),
    .A2(net908),
    .Y(_1559_),
    .B1(net991));
 sg13g2_a22oi_1 _5388_ (.Y(_1560_),
    .B1(net896),
    .B2(\led_controller.colors[6] ),
    .A2(net902),
    .A1(\led_controller.colors[70] ));
 sg13g2_nand2_1 _5389_ (.Y(_1561_),
    .A(_1559_),
    .B(_1560_));
 sg13g2_a21oi_1 _5390_ (.A1(_0787_),
    .A2(net998),
    .Y(_1562_),
    .B1(net864));
 sg13g2_a22oi_1 _5391_ (.Y(_1563_),
    .B1(_1561_),
    .B2(_1562_),
    .A2(net860),
    .A1(net1663));
 sg13g2_nor2_1 _5392_ (.A(net1125),
    .B(net1664),
    .Y(_0230_));
 sg13g2_a21oi_1 _5393_ (.A1(\led_controller.colors[39] ),
    .A2(net908),
    .Y(_1564_),
    .B1(net991));
 sg13g2_a22oi_1 _5394_ (.Y(_1565_),
    .B1(net897),
    .B2(\led_controller.colors[7] ),
    .A2(net903),
    .A1(\led_controller.colors[71] ));
 sg13g2_nand2_1 _5395_ (.Y(_1566_),
    .A(_1564_),
    .B(_1565_));
 sg13g2_a21oi_1 _5396_ (.A1(_0786_),
    .A2(net996),
    .Y(_1567_),
    .B1(net861));
 sg13g2_a22oi_1 _5397_ (.Y(_1568_),
    .B1(_1566_),
    .B2(_1567_),
    .A2(net856),
    .A1(net1659));
 sg13g2_nor2_1 _5398_ (.A(net1114),
    .B(net1660),
    .Y(_0231_));
 sg13g2_a21oi_1 _5399_ (.A1(\led_controller.colors[40] ),
    .A2(net912),
    .Y(_1569_),
    .B1(net996));
 sg13g2_a22oi_1 _5400_ (.Y(_1570_),
    .B1(net900),
    .B2(\led_controller.colors[8] ),
    .A2(net906),
    .A1(\led_controller.colors[72] ));
 sg13g2_nand2_1 _5401_ (.Y(_1571_),
    .A(_1569_),
    .B(_1570_));
 sg13g2_a21oi_1 _5402_ (.A1(_0785_),
    .A2(net999),
    .Y(_1572_),
    .B1(net862));
 sg13g2_a22oi_1 _5403_ (.Y(_1573_),
    .B1(_1571_),
    .B2(_1572_),
    .A2(net862),
    .A1(net1641));
 sg13g2_nor2_1 _5404_ (.A(net1128),
    .B(net1642),
    .Y(_0232_));
 sg13g2_a21oi_1 _5405_ (.A1(net1858),
    .A2(net910),
    .Y(_1574_),
    .B1(net995));
 sg13g2_a22oi_1 _5406_ (.Y(_1575_),
    .B1(net898),
    .B2(\led_controller.colors[9] ),
    .A2(net904),
    .A1(\led_controller.colors[73] ));
 sg13g2_nand2_1 _5407_ (.Y(_1576_),
    .A(_1574_),
    .B(_1575_));
 sg13g2_a21oi_1 _5408_ (.A1(_0784_),
    .A2(net994),
    .Y(_1577_),
    .B1(net858));
 sg13g2_a22oi_1 _5409_ (.Y(_1578_),
    .B1(_1576_),
    .B2(_1577_),
    .A2(net858),
    .A1(net2004));
 sg13g2_nor2_1 _5410_ (.A(net1121),
    .B(net2005),
    .Y(_0233_));
 sg13g2_a21oi_1 _5411_ (.A1(\led_controller.colors[42] ),
    .A2(net910),
    .Y(_1579_),
    .B1(net993));
 sg13g2_a22oi_1 _5412_ (.Y(_1580_),
    .B1(net898),
    .B2(\led_controller.colors[10] ),
    .A2(net904),
    .A1(\led_controller.colors[74] ));
 sg13g2_nand2_1 _5413_ (.Y(_1581_),
    .A(_1579_),
    .B(_1580_));
 sg13g2_a21oi_1 _5414_ (.A1(_0783_),
    .A2(net999),
    .Y(_1582_),
    .B1(net858));
 sg13g2_a22oi_1 _5415_ (.Y(_1583_),
    .B1(_1581_),
    .B2(_1582_),
    .A2(net859),
    .A1(net1716));
 sg13g2_nor2_1 _5416_ (.A(net1128),
    .B(net1717),
    .Y(_0234_));
 sg13g2_a21oi_1 _5417_ (.A1(\led_controller.colors[43] ),
    .A2(net910),
    .Y(_1584_),
    .B1(net995));
 sg13g2_a22oi_1 _5418_ (.Y(_1585_),
    .B1(net898),
    .B2(\led_controller.colors[11] ),
    .A2(net904),
    .A1(\led_controller.colors[75] ));
 sg13g2_nand2_1 _5419_ (.Y(_1586_),
    .A(_1584_),
    .B(_1585_));
 sg13g2_a21oi_1 _5420_ (.A1(_0782_),
    .A2(net999),
    .Y(_1587_),
    .B1(net859));
 sg13g2_a22oi_1 _5421_ (.Y(_1588_),
    .B1(_1586_),
    .B2(_1587_),
    .A2(net859),
    .A1(net1760));
 sg13g2_nor2_1 _5422_ (.A(net1128),
    .B(net1761),
    .Y(_0235_));
 sg13g2_a21oi_1 _5423_ (.A1(\led_controller.colors[44] ),
    .A2(net909),
    .Y(_1589_),
    .B1(net993));
 sg13g2_a22oi_1 _5424_ (.Y(_1590_),
    .B1(net897),
    .B2(\led_controller.colors[12] ),
    .A2(net903),
    .A1(\led_controller.colors[76] ));
 sg13g2_nand2_1 _5425_ (.Y(_1591_),
    .A(_1589_),
    .B(_1590_));
 sg13g2_a21oi_1 _5426_ (.A1(_0781_),
    .A2(net992),
    .Y(_1592_),
    .B1(net866));
 sg13g2_a22oi_1 _5427_ (.Y(_1593_),
    .B1(_1591_),
    .B2(_1592_),
    .A2(net857),
    .A1(net1721));
 sg13g2_nor2_1 _5428_ (.A(net1125),
    .B(net1722),
    .Y(_0236_));
 sg13g2_a21oi_1 _5429_ (.A1(\led_controller.colors[45] ),
    .A2(net908),
    .Y(_1594_),
    .B1(net993));
 sg13g2_a22oi_1 _5430_ (.Y(_1595_),
    .B1(net896),
    .B2(\led_controller.colors[13] ),
    .A2(net902),
    .A1(\led_controller.colors[77] ));
 sg13g2_nand2_1 _5431_ (.Y(_1596_),
    .A(_1594_),
    .B(_1595_));
 sg13g2_a21oi_1 _5432_ (.A1(_0780_),
    .A2(net998),
    .Y(_1597_),
    .B1(net865));
 sg13g2_a22oi_1 _5433_ (.Y(_1598_),
    .B1(_1596_),
    .B2(_1597_),
    .A2(net857),
    .A1(net1730));
 sg13g2_nor2_1 _5434_ (.A(net1115),
    .B(net1731),
    .Y(_0237_));
 sg13g2_a21oi_1 _5435_ (.A1(net1679),
    .A2(net909),
    .Y(_1599_),
    .B1(net991));
 sg13g2_a22oi_1 _5436_ (.Y(_1600_),
    .B1(net897),
    .B2(\led_controller.colors[14] ),
    .A2(net903),
    .A1(\led_controller.colors[78] ));
 sg13g2_nand2_1 _5437_ (.Y(_1601_),
    .A(_1599_),
    .B(_1600_));
 sg13g2_a21oi_1 _5438_ (.A1(_0779_),
    .A2(net992),
    .Y(_1602_),
    .B1(net860));
 sg13g2_a22oi_1 _5439_ (.Y(_1603_),
    .B1(_1601_),
    .B2(_1602_),
    .A2(net860),
    .A1(net1711));
 sg13g2_nor2_1 _5440_ (.A(net1125),
    .B(net1712),
    .Y(_0238_));
 sg13g2_a21oi_1 _5441_ (.A1(\led_controller.colors[47] ),
    .A2(net908),
    .Y(_1604_),
    .B1(net991));
 sg13g2_a22oi_1 _5442_ (.Y(_1605_),
    .B1(net896),
    .B2(\led_controller.colors[15] ),
    .A2(net902),
    .A1(\led_controller.colors[79] ));
 sg13g2_nand2_1 _5443_ (.Y(_1606_),
    .A(_1604_),
    .B(_1605_));
 sg13g2_a21oi_2 _5444_ (.B1(net863),
    .Y(_1607_),
    .A2(net997),
    .A1(_0778_));
 sg13g2_a22oi_1 _5445_ (.Y(_1608_),
    .B1(_1606_),
    .B2(_1607_),
    .A2(net856),
    .A1(net1779));
 sg13g2_nor2_1 _5446_ (.A(net1114),
    .B(net1780),
    .Y(_0239_));
 sg13g2_a21oi_1 _5447_ (.A1(\led_controller.colors[48] ),
    .A2(net912),
    .Y(_1609_),
    .B1(net996));
 sg13g2_a22oi_1 _5448_ (.Y(_1610_),
    .B1(net899),
    .B2(\led_controller.colors[16] ),
    .A2(net905),
    .A1(\led_controller.colors[80] ));
 sg13g2_nand2_1 _5449_ (.Y(_1611_),
    .A(_1609_),
    .B(_1610_));
 sg13g2_a21oi_1 _5450_ (.A1(_0777_),
    .A2(net998),
    .Y(_1612_),
    .B1(net864));
 sg13g2_a22oi_1 _5451_ (.Y(_1613_),
    .B1(_1611_),
    .B2(_1612_),
    .A2(net863),
    .A1(net1637));
 sg13g2_nor2_1 _5452_ (.A(net1129),
    .B(net1638),
    .Y(_0240_));
 sg13g2_a21oi_1 _5453_ (.A1(\led_controller.colors[49] ),
    .A2(net910),
    .Y(_1614_),
    .B1(net995));
 sg13g2_a22oi_1 _5454_ (.Y(_1615_),
    .B1(net898),
    .B2(\led_controller.colors[17] ),
    .A2(net904),
    .A1(\led_controller.colors[81] ));
 sg13g2_nand2_1 _5455_ (.Y(_1616_),
    .A(_1614_),
    .B(_1615_));
 sg13g2_a21oi_1 _5456_ (.A1(_0776_),
    .A2(net999),
    .Y(_1617_),
    .B1(net862));
 sg13g2_a22oi_1 _5457_ (.Y(_1618_),
    .B1(_1616_),
    .B2(_1617_),
    .A2(net863),
    .A1(net1647));
 sg13g2_nor2_1 _5458_ (.A(net1129),
    .B(net1648),
    .Y(_0241_));
 sg13g2_a21oi_1 _5459_ (.A1(\led_controller.colors[50] ),
    .A2(net910),
    .Y(_1619_),
    .B1(net994));
 sg13g2_a22oi_1 _5460_ (.Y(_1620_),
    .B1(net900),
    .B2(\led_controller.colors[18] ),
    .A2(net906),
    .A1(\led_controller.colors[82] ));
 sg13g2_nand2_1 _5461_ (.Y(_1621_),
    .A(_1619_),
    .B(_1620_));
 sg13g2_a21oi_1 _5462_ (.A1(_0775_),
    .A2(net999),
    .Y(_1622_),
    .B1(net862));
 sg13g2_a22oi_1 _5463_ (.Y(_1623_),
    .B1(_1621_),
    .B2(_1622_),
    .A2(net859),
    .A1(net1667));
 sg13g2_nor2_1 _5464_ (.A(net1128),
    .B(net1668),
    .Y(_0242_));
 sg13g2_a21oi_1 _5465_ (.A1(\led_controller.colors[51] ),
    .A2(net911),
    .Y(_1624_),
    .B1(net994));
 sg13g2_a22oi_1 _5466_ (.Y(_1625_),
    .B1(net899),
    .B2(\led_controller.colors[19] ),
    .A2(net905),
    .A1(\led_controller.colors[83] ));
 sg13g2_nand2_1 _5467_ (.Y(_1626_),
    .A(_1624_),
    .B(_1625_));
 sg13g2_a21oi_1 _5468_ (.A1(_0774_),
    .A2(net999),
    .Y(_1627_),
    .B1(net858));
 sg13g2_a22oi_1 _5469_ (.Y(_1628_),
    .B1(_1626_),
    .B2(_1627_),
    .A2(net859),
    .A1(net1740));
 sg13g2_nor2_1 _5470_ (.A(net1128),
    .B(net1741),
    .Y(_0243_));
 sg13g2_a21oi_1 _5471_ (.A1(\led_controller.colors[52] ),
    .A2(net912),
    .Y(_1629_),
    .B1(net992));
 sg13g2_a22oi_1 _5472_ (.Y(_1630_),
    .B1(net899),
    .B2(\led_controller.colors[20] ),
    .A2(net905),
    .A1(\led_controller.colors[84] ));
 sg13g2_nand2_1 _5473_ (.Y(_1631_),
    .A(_1629_),
    .B(_1630_));
 sg13g2_a21oi_1 _5474_ (.A1(_0773_),
    .A2(net996),
    .Y(_1632_),
    .B1(net861));
 sg13g2_a22oi_1 _5475_ (.Y(_1633_),
    .B1(_1631_),
    .B2(_1632_),
    .A2(net861),
    .A1(net1677));
 sg13g2_nor2_1 _5476_ (.A(net1126),
    .B(net1678),
    .Y(_0244_));
 sg13g2_a21oi_1 _5477_ (.A1(\led_controller.colors[53] ),
    .A2(net908),
    .Y(_1634_),
    .B1(net991));
 sg13g2_a22oi_1 _5478_ (.Y(_1635_),
    .B1(net896),
    .B2(\led_controller.colors[21] ),
    .A2(net902),
    .A1(\led_controller.colors[85] ));
 sg13g2_nand2_1 _5479_ (.Y(_1636_),
    .A(_1634_),
    .B(_1635_));
 sg13g2_a21oi_1 _5480_ (.A1(_0772_),
    .A2(net996),
    .Y(_1637_),
    .B1(net861));
 sg13g2_a22oi_1 _5481_ (.Y(_1638_),
    .B1(_1636_),
    .B2(_1637_),
    .A2(net856),
    .A1(net1681));
 sg13g2_nor2_1 _5482_ (.A(net1115),
    .B(net1682),
    .Y(_0245_));
 sg13g2_a21oi_1 _5483_ (.A1(\led_controller.colors[54] ),
    .A2(net909),
    .Y(_1639_),
    .B1(net991));
 sg13g2_a22oi_1 _5484_ (.Y(_1640_),
    .B1(net897),
    .B2(\led_controller.colors[22] ),
    .A2(net903),
    .A1(\led_controller.colors[86] ));
 sg13g2_nand2_1 _5485_ (.Y(_1641_),
    .A(_1639_),
    .B(_1640_));
 sg13g2_a21oi_1 _5486_ (.A1(_0771_),
    .A2(net996),
    .Y(_1642_),
    .B1(net860));
 sg13g2_a22oi_1 _5487_ (.Y(_1643_),
    .B1(_1641_),
    .B2(_1642_),
    .A2(net861),
    .A1(net1781));
 sg13g2_nor2_1 _5488_ (.A(net1126),
    .B(net1782),
    .Y(_0246_));
 sg13g2_a21oi_1 _5489_ (.A1(\led_controller.colors[55] ),
    .A2(net908),
    .Y(_1644_),
    .B1(net991));
 sg13g2_a22oi_1 _5490_ (.Y(_1645_),
    .B1(net896),
    .B2(\led_controller.colors[23] ),
    .A2(net902),
    .A1(\led_controller.colors[87] ));
 sg13g2_nand2_1 _5491_ (.Y(_1646_),
    .A(_1644_),
    .B(_1645_));
 sg13g2_a21oi_1 _5492_ (.A1(_0770_),
    .A2(net1000),
    .Y(_1647_),
    .B1(net865));
 sg13g2_a22oi_1 _5493_ (.Y(_1648_),
    .B1(_1646_),
    .B2(_1647_),
    .A2(net856),
    .A1(net1673));
 sg13g2_nor2_1 _5494_ (.A(net1114),
    .B(net1674),
    .Y(_0247_));
 sg13g2_a21oi_1 _5495_ (.A1(\led_controller.colors[56] ),
    .A2(net912),
    .Y(_1649_),
    .B1(net1000));
 sg13g2_a22oi_1 _5496_ (.Y(_1650_),
    .B1(net899),
    .B2(\led_controller.colors[24] ),
    .A2(net905),
    .A1(\led_controller.colors[88] ));
 sg13g2_nand2_1 _5497_ (.Y(_1651_),
    .A(_1649_),
    .B(_1650_));
 sg13g2_a21oi_1 _5498_ (.A1(_0769_),
    .A2(net997),
    .Y(_1652_),
    .B1(net864));
 sg13g2_a22oi_1 _5499_ (.Y(_1653_),
    .B1(_1651_),
    .B2(_1652_),
    .A2(net864),
    .A1(net1661));
 sg13g2_nor2_1 _5500_ (.A(net1129),
    .B(net1662),
    .Y(_0248_));
 sg13g2_a21oi_1 _5501_ (.A1(\led_controller.colors[57] ),
    .A2(net911),
    .Y(_1654_),
    .B1(net1001));
 sg13g2_a22oi_1 _5502_ (.Y(_1655_),
    .B1(net898),
    .B2(\led_controller.colors[25] ),
    .A2(net904),
    .A1(\led_controller.colors[89] ));
 sg13g2_nand2_1 _5503_ (.Y(_1656_),
    .A(_1654_),
    .B(_1655_));
 sg13g2_a21oi_1 _5504_ (.A1(_0768_),
    .A2(net997),
    .Y(_1657_),
    .B1(net865));
 sg13g2_a22oi_1 _5505_ (.Y(_1658_),
    .B1(_1656_),
    .B2(_1657_),
    .A2(net864),
    .A1(net1700));
 sg13g2_nor2_1 _5506_ (.A(net1129),
    .B(net1701),
    .Y(_0249_));
 sg13g2_a21oi_1 _5507_ (.A1(\led_controller.colors[58] ),
    .A2(net910),
    .Y(_1659_),
    .B1(net995));
 sg13g2_a22oi_1 _5508_ (.Y(_1660_),
    .B1(net898),
    .B2(\led_controller.colors[26] ),
    .A2(net904),
    .A1(\led_controller.colors[90] ));
 sg13g2_nand2_1 _5509_ (.Y(_1661_),
    .A(_1659_),
    .B(_1660_));
 sg13g2_a21oi_1 _5510_ (.A1(_0767_),
    .A2(net997),
    .Y(_1662_),
    .B1(net864));
 sg13g2_a22oi_1 _5511_ (.Y(_1663_),
    .B1(_1661_),
    .B2(_1662_),
    .A2(net861),
    .A1(net1639));
 sg13g2_nor2_1 _5512_ (.A(net1126),
    .B(net1640),
    .Y(_0250_));
 sg13g2_a21oi_1 _5513_ (.A1(\led_controller.colors[59] ),
    .A2(net911),
    .Y(_1664_),
    .B1(net995));
 sg13g2_a22oi_1 _5514_ (.Y(_1665_),
    .B1(net899),
    .B2(\led_controller.colors[27] ),
    .A2(net905),
    .A1(net2011));
 sg13g2_nand2_1 _5515_ (.Y(_1666_),
    .A(_1664_),
    .B(_1665_));
 sg13g2_a21oi_1 _5516_ (.A1(_0766_),
    .A2(net997),
    .Y(_1667_),
    .B1(net863));
 sg13g2_a22oi_1 _5517_ (.Y(_1668_),
    .B1(_1666_),
    .B2(_1667_),
    .A2(net863),
    .A1(net2026));
 sg13g2_nor2_1 _5518_ (.A(net1126),
    .B(net2027),
    .Y(_0251_));
 sg13g2_a21oi_1 _5519_ (.A1(\led_controller.colors[60] ),
    .A2(net909),
    .Y(_1669_),
    .B1(net992));
 sg13g2_a22oi_1 _5520_ (.Y(_1670_),
    .B1(net900),
    .B2(\led_controller.colors[28] ),
    .A2(net906),
    .A1(\led_controller.colors[92] ));
 sg13g2_nand2_1 _5521_ (.Y(_1671_),
    .A(_1669_),
    .B(_1670_));
 sg13g2_a21oi_1 _5522_ (.A1(_0765_),
    .A2(net992),
    .Y(_1672_),
    .B1(net860));
 sg13g2_a22oi_1 _5523_ (.Y(_1673_),
    .B1(_1671_),
    .B2(_1672_),
    .A2(net860),
    .A1(net1754));
 sg13g2_nor2_1 _5524_ (.A(net1125),
    .B(net1755),
    .Y(_0252_));
 sg13g2_a21oi_1 _5525_ (.A1(\led_controller.colors[61] ),
    .A2(net908),
    .Y(_1674_),
    .B1(net992));
 sg13g2_a22oi_1 _5526_ (.Y(_1675_),
    .B1(net896),
    .B2(\led_controller.colors[29] ),
    .A2(net902),
    .A1(\led_controller.colors[93] ));
 sg13g2_nand2_1 _5527_ (.Y(_1676_),
    .A(_1674_),
    .B(_1675_));
 sg13g2_a21oi_1 _5528_ (.A1(_0764_),
    .A2(net997),
    .Y(_1677_),
    .B1(net865));
 sg13g2_a22oi_1 _5529_ (.Y(_1678_),
    .B1(_1676_),
    .B2(_1677_),
    .A2(net857),
    .A1(net1726));
 sg13g2_nor2_1 _5530_ (.A(net1115),
    .B(net1727),
    .Y(_0253_));
 sg13g2_a21oi_1 _5531_ (.A1(\led_controller.colors[62] ),
    .A2(net908),
    .Y(_1679_),
    .B1(net991));
 sg13g2_a22oi_1 _5532_ (.Y(_1680_),
    .B1(net896),
    .B2(\led_controller.colors[30] ),
    .A2(net902),
    .A1(\led_controller.colors[94] ));
 sg13g2_nand2_1 _5533_ (.Y(_1681_),
    .A(_1679_),
    .B(_1680_));
 sg13g2_a21oi_1 _5534_ (.A1(_0763_),
    .A2(net1000),
    .Y(_1682_),
    .B1(net860));
 sg13g2_a22oi_1 _5535_ (.Y(_1683_),
    .B1(_1681_),
    .B2(_1682_),
    .A2(net857),
    .A1(net1671));
 sg13g2_nor2_1 _5536_ (.A(net1125),
    .B(net1672),
    .Y(_0254_));
 sg13g2_a21oi_1 _5537_ (.A1(\led_controller.colors[63] ),
    .A2(net909),
    .Y(_1684_),
    .B1(net992));
 sg13g2_a22oi_1 _5538_ (.Y(_1685_),
    .B1(net896),
    .B2(\led_controller.colors[31] ),
    .A2(net902),
    .A1(\led_controller.colors[95] ));
 sg13g2_nand2_1 _5539_ (.Y(_1686_),
    .A(_1684_),
    .B(_1685_));
 sg13g2_a21oi_1 _5540_ (.A1(_0762_),
    .A2(net996),
    .Y(_1687_),
    .B1(net865));
 sg13g2_a22oi_1 _5541_ (.Y(_1688_),
    .B1(_1686_),
    .B2(_1687_),
    .A2(net856),
    .A1(net1702));
 sg13g2_nor2_1 _5542_ (.A(net1114),
    .B(net1703),
    .Y(_0255_));
 sg13g2_o21ai_1 _5543_ (.B1(_1500_),
    .Y(_1689_),
    .A1(_1494_),
    .A2(_1501_));
 sg13g2_inv_2 _5544_ (.Y(_1690_),
    .A(net822));
 sg13g2_nor2_1 _5545_ (.A(_0932_),
    .B(_1496_),
    .Y(_1691_));
 sg13g2_nand2_1 _5546_ (.Y(_1692_),
    .A(_0933_),
    .B(_1497_));
 sg13g2_nor2_1 _5547_ (.A(net822),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_nand2_1 _5548_ (.Y(_1694_),
    .A(\led_controller.rgbw.color[5] ),
    .B(net1020));
 sg13g2_a21oi_1 _5549_ (.A1(\led_controller.rgbw.color[13] ),
    .A2(_1512_),
    .Y(_1695_),
    .B1(net1190));
 sg13g2_nand2_1 _5550_ (.Y(_1696_),
    .A(\led_controller.rgbw.color[12] ),
    .B(_1512_));
 sg13g2_a21oi_1 _5551_ (.A1(\led_controller.rgbw.color[4] ),
    .A2(net1020),
    .Y(_1697_),
    .B1(net1189));
 sg13g2_a221oi_1 _5552_ (.B2(_1697_),
    .C1(_1515_),
    .B1(_1696_),
    .A1(_1694_),
    .Y(_1698_),
    .A2(_1695_));
 sg13g2_nand2_1 _5553_ (.Y(_1699_),
    .A(\led_controller.rgbw.color[28] ),
    .B(_1512_));
 sg13g2_a21oi_1 _5554_ (.A1(\led_controller.rgbw.color[20] ),
    .A2(net1020),
    .Y(_1700_),
    .B1(net1189));
 sg13g2_nand2_1 _5555_ (.Y(_1701_),
    .A(\led_controller.rgbw.color[21] ),
    .B(net1020));
 sg13g2_a21oi_1 _5556_ (.A1(\led_controller.rgbw.color[29] ),
    .A2(_1512_),
    .Y(_1702_),
    .B1(net1190));
 sg13g2_a221oi_1 _5557_ (.B2(_1702_),
    .C1(_1514_),
    .B1(_1701_),
    .A1(_1699_),
    .Y(_1703_),
    .A2(_1700_));
 sg13g2_nor3_1 _5558_ (.A(_1507_),
    .B(_1698_),
    .C(_1703_),
    .Y(_1704_));
 sg13g2_mux4_1 _5559_ (.S0(net1020),
    .A0(\led_controller.rgbw.color[30] ),
    .A1(\led_controller.rgbw.color[22] ),
    .A2(\led_controller.rgbw.color[14] ),
    .A3(\led_controller.rgbw.color[6] ),
    .S1(_1514_),
    .X(_1705_));
 sg13g2_nand2b_1 _5560_ (.Y(_1706_),
    .B(net1097),
    .A_N(_1705_));
 sg13g2_mux4_1 _5561_ (.S0(net1020),
    .A0(\led_controller.rgbw.color[31] ),
    .A1(\led_controller.rgbw.color[23] ),
    .A2(\led_controller.rgbw.color[15] ),
    .A3(\led_controller.rgbw.color[7] ),
    .S1(_1514_),
    .X(_1707_));
 sg13g2_o21ai_1 _5562_ (.B1(_1706_),
    .Y(_1708_),
    .A1(\led_controller.rgbw.pixel_counter[2] ),
    .A2(_1707_));
 sg13g2_o21ai_1 _5563_ (.B1(_1509_),
    .Y(_1709_),
    .A1(_1704_),
    .A2(_1708_));
 sg13g2_a22oi_1 _5564_ (.Y(_1710_),
    .B1(net1190),
    .B2(\led_controller.rgbw.color[24] ),
    .A2(net1189),
    .A1(\led_controller.rgbw.color[25] ));
 sg13g2_or2_1 _5565_ (.X(_1711_),
    .B(_1710_),
    .A(net1097));
 sg13g2_a22oi_1 _5566_ (.Y(_1712_),
    .B1(net1097),
    .B2(\led_controller.rgbw.color[26] ),
    .A2(\led_controller.rgbw.pixel_counter[2] ),
    .A1(\led_controller.rgbw.color[27] ));
 sg13g2_a22oi_1 _5567_ (.Y(_1713_),
    .B1(\led_controller.rgbw.pixel_counter[0] ),
    .B2(\led_controller.rgbw.color[16] ),
    .A2(net1189),
    .A1(\led_controller.rgbw.color[17] ));
 sg13g2_a22oi_1 _5568_ (.Y(_1714_),
    .B1(net1097),
    .B2(\led_controller.rgbw.color[18] ),
    .A2(_0965_),
    .A1(\led_controller.rgbw.color[19] ));
 sg13g2_o21ai_1 _5569_ (.B1(_1714_),
    .Y(_1715_),
    .A1(net1097),
    .A2(_1713_));
 sg13g2_a21oi_1 _5570_ (.A1(_1711_),
    .A2(_1712_),
    .Y(_1716_),
    .B1(net1020));
 sg13g2_a21oi_1 _5571_ (.A1(_1511_),
    .A2(_1715_),
    .Y(_1717_),
    .B1(_1716_));
 sg13g2_a22oi_1 _5572_ (.Y(_1718_),
    .B1(\led_controller.rgbw.pixel_counter[0] ),
    .B2(\led_controller.rgbw.color[8] ),
    .A2(\led_controller.rgbw.pixel_counter[1] ),
    .A1(\led_controller.rgbw.color[9] ));
 sg13g2_a22oi_1 _5573_ (.Y(_1719_),
    .B1(net1097),
    .B2(\led_controller.rgbw.color[10] ),
    .A2(_0965_),
    .A1(\led_controller.rgbw.color[11] ));
 sg13g2_o21ai_1 _5574_ (.B1(_1719_),
    .Y(_1720_),
    .A1(net1097),
    .A2(_1718_));
 sg13g2_a22oi_1 _5575_ (.Y(_1721_),
    .B1(\led_controller.rgbw.pixel_counter[0] ),
    .B2(\led_controller.rgbw.color[0] ),
    .A2(\led_controller.rgbw.pixel_counter[1] ),
    .A1(\led_controller.rgbw.color[1] ));
 sg13g2_a22oi_1 _5576_ (.Y(_1722_),
    .B1(_1506_),
    .B2(\led_controller.rgbw.color[2] ),
    .A2(_0965_),
    .A1(\led_controller.rgbw.color[3] ));
 sg13g2_o21ai_1 _5577_ (.B1(_1722_),
    .Y(_1723_),
    .A1(_1506_),
    .A2(_1721_));
 sg13g2_mux2_1 _5578_ (.A0(_1720_),
    .A1(_1723_),
    .S(_1511_),
    .X(_1724_));
 sg13g2_a21oi_1 _5579_ (.A1(_1514_),
    .A2(_1724_),
    .Y(_1725_),
    .B1(_1509_));
 sg13g2_o21ai_1 _5580_ (.B1(_1725_),
    .Y(_1726_),
    .A1(_1514_),
    .A2(_1717_));
 sg13g2_nand3_1 _5581_ (.B(_1709_),
    .C(_1726_),
    .A(_1518_),
    .Y(_1727_));
 sg13g2_or2_1 _5582_ (.X(_1728_),
    .B(_1727_),
    .A(_0933_));
 sg13g2_or2_1 _5583_ (.X(_1729_),
    .B(_1728_),
    .A(_0883_));
 sg13g2_o21ai_1 _5584_ (.B1(_1729_),
    .Y(_1730_),
    .A1(net2172),
    .A2(_1692_));
 sg13g2_nor2_1 _5585_ (.A(net822),
    .B(_1730_),
    .Y(_1731_));
 sg13g2_o21ai_1 _5586_ (.B1(net1153),
    .Y(_1732_),
    .A1(net2172),
    .A2(_1690_));
 sg13g2_nor2_1 _5587_ (.A(_1731_),
    .B(_1732_),
    .Y(_0256_));
 sg13g2_a21o_1 _5588_ (.A2(_1691_),
    .A1(\led_controller.rgbw.low_cycles[0] ),
    .B1(net822),
    .X(_1733_));
 sg13g2_a22oi_1 _5589_ (.Y(_1734_),
    .B1(_1733_),
    .B2(net1704),
    .A2(_1693_),
    .A1(_0924_));
 sg13g2_nor2_1 _5590_ (.A(net1111),
    .B(net1705),
    .Y(_0257_));
 sg13g2_nor2b_1 _5591_ (.A(_0924_),
    .B_N(net2112),
    .Y(_1735_));
 sg13g2_a221oi_1 _5592_ (.B2(_1497_),
    .C1(net823),
    .B1(_1735_),
    .A1(_0925_),
    .Y(_1736_),
    .A2(_1691_));
 sg13g2_o21ai_1 _5593_ (.B1(net1153),
    .Y(_1737_),
    .A1(net2112),
    .A2(_1690_));
 sg13g2_a21oi_1 _5594_ (.A1(_1729_),
    .A2(_1736_),
    .Y(_0258_),
    .B1(_1737_));
 sg13g2_nor2_1 _5595_ (.A(_0933_),
    .B(_0968_),
    .Y(_1738_));
 sg13g2_and2_1 _5596_ (.A(_1727_),
    .B(_1738_),
    .X(_1739_));
 sg13g2_nand2b_1 _5597_ (.Y(_1740_),
    .B(net2028),
    .A_N(_0925_));
 sg13g2_o21ai_1 _5598_ (.B1(_1740_),
    .Y(_1741_),
    .A1(_0926_),
    .A2(_0932_));
 sg13g2_a221oi_1 _5599_ (.B2(_1497_),
    .C1(net823),
    .B1(_1741_),
    .A1(\led_controller.rgbw.state[2] ),
    .Y(_1742_),
    .A2(_1739_));
 sg13g2_o21ai_1 _5600_ (.B1(net1153),
    .Y(_1743_),
    .A1(net2028),
    .A2(_1690_));
 sg13g2_nor2_1 _5601_ (.A(_1742_),
    .B(_1743_),
    .Y(_0259_));
 sg13g2_nor2_1 _5602_ (.A(_0927_),
    .B(_0932_),
    .Y(_1744_));
 sg13g2_a21oi_1 _5603_ (.A1(net1646),
    .A2(_0926_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_nor2_1 _5604_ (.A(_1496_),
    .B(_1745_),
    .Y(_1746_));
 sg13g2_o21ai_1 _5605_ (.B1(net1153),
    .Y(_1747_),
    .A1(net822),
    .A2(_1746_));
 sg13g2_a21oi_1 _5606_ (.A1(_0874_),
    .A2(net822),
    .Y(_0260_),
    .B1(_1747_));
 sg13g2_a21oi_1 _5607_ (.A1(_1690_),
    .A2(_1744_),
    .Y(_1748_),
    .B1(net2164));
 sg13g2_a21oi_1 _5608_ (.A1(net2164),
    .A2(_0928_),
    .Y(_1749_),
    .B1(_1496_));
 sg13g2_nor2_1 _5609_ (.A(net822),
    .B(_1749_),
    .Y(_1750_));
 sg13g2_o21ai_1 _5610_ (.B1(net1153),
    .Y(_0261_),
    .A1(_1748_),
    .A2(_1750_));
 sg13g2_o21ai_1 _5611_ (.B1(net2096),
    .Y(_1751_),
    .A1(\led_controller.rgbw.low_cycles[5] ),
    .A2(_0927_));
 sg13g2_nand2b_1 _5612_ (.Y(_1752_),
    .B(_1751_),
    .A_N(_0929_));
 sg13g2_a22oi_1 _5613_ (.Y(_1753_),
    .B1(_1693_),
    .B2(_1752_),
    .A2(net823),
    .A1(net2096));
 sg13g2_nor2_1 _5614_ (.A(net1111),
    .B(net2097),
    .Y(_0262_));
 sg13g2_xor2_1 _5615_ (.B(_0929_),
    .A(net2092),
    .X(_1754_));
 sg13g2_a22oi_1 _5616_ (.Y(_1755_),
    .B1(_1693_),
    .B2(_1754_),
    .A2(net823),
    .A1(net2092));
 sg13g2_nor2_1 _5617_ (.A(net1111),
    .B(net2093),
    .Y(_0263_));
 sg13g2_and2_1 _5618_ (.A(net2099),
    .B(_0930_),
    .X(_1756_));
 sg13g2_a21oi_1 _5619_ (.A1(net1890),
    .A2(_0931_),
    .Y(_1757_),
    .B1(_1756_));
 sg13g2_nor3_1 _5620_ (.A(_1496_),
    .B(net823),
    .C(_1757_),
    .Y(_1758_));
 sg13g2_a21oi_1 _5621_ (.A1(net2099),
    .A2(net822),
    .Y(_1759_),
    .B1(_1758_));
 sg13g2_nand2_1 _5622_ (.Y(_0264_),
    .A(net1153),
    .B(_1759_));
 sg13g2_o21ai_1 _5623_ (.B1(_1690_),
    .Y(_1760_),
    .A1(_0931_),
    .A2(_1496_));
 sg13g2_a21o_1 _5624_ (.A2(_1760_),
    .A1(net1890),
    .B1(net1117),
    .X(_0265_));
 sg13g2_a21oi_2 _5625_ (.B1(_1492_),
    .Y(_1761_),
    .A2(_1494_),
    .A1(_0933_));
 sg13g2_o21ai_1 _5626_ (.B1(_1761_),
    .Y(_1762_),
    .A1(net2268),
    .A2(_0932_));
 sg13g2_nor2_1 _5627_ (.A(_1739_),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_o21ai_1 _5628_ (.B1(net1152),
    .Y(_1764_),
    .A1(net2268),
    .A2(_1761_));
 sg13g2_nor2_1 _5629_ (.A(_1763_),
    .B(_1764_),
    .Y(_0266_));
 sg13g2_xnor2_1 _5630_ (.Y(_1765_),
    .A(net2188),
    .B(\led_controller.rgbw.high_cycles[0] ));
 sg13g2_a21oi_1 _5631_ (.A1(_0933_),
    .A2(_1765_),
    .Y(_1766_),
    .B1(_1738_));
 sg13g2_o21ai_1 _5632_ (.B1(net1152),
    .Y(_1767_),
    .A1(net2188),
    .A2(_1761_));
 sg13g2_a21oi_1 _5633_ (.A1(_1761_),
    .A2(_1766_),
    .Y(_0267_),
    .B1(_1767_));
 sg13g2_o21ai_1 _5634_ (.B1(net2109),
    .Y(_1768_),
    .A1(\led_controller.rgbw.high_cycles[1] ),
    .A2(\led_controller.rgbw.high_cycles[0] ));
 sg13g2_o21ai_1 _5635_ (.B1(_1761_),
    .Y(_1769_),
    .A1(_0932_),
    .A2(_1768_));
 sg13g2_inv_1 _5636_ (.Y(_1770_),
    .A(_1769_));
 sg13g2_o21ai_1 _5637_ (.B1(net1152),
    .Y(_1771_),
    .A1(net2109),
    .A2(_1761_));
 sg13g2_a21oi_1 _5638_ (.A1(_1728_),
    .A2(_1770_),
    .Y(_0268_),
    .B1(_1771_));
 sg13g2_and2_1 _5639_ (.A(net1176),
    .B(_1009_),
    .X(_1772_));
 sg13g2_and2_1 _5640_ (.A(_0798_),
    .B(_1772_),
    .X(_1773_));
 sg13g2_nand2_2 _5641_ (.Y(_1774_),
    .A(_0798_),
    .B(_1772_));
 sg13g2_and2_1 _5642_ (.A(net2310),
    .B(net967),
    .X(_1775_));
 sg13g2_nor2_2 _5643_ (.A(net1176),
    .B(_1010_),
    .Y(_1776_));
 sg13g2_nor3_1 _5644_ (.A(net2310),
    .B(net967),
    .C(_1776_),
    .Y(_1777_));
 sg13g2_nor3_1 _5645_ (.A(net1040),
    .B(_1775_),
    .C(_1777_),
    .Y(_0269_));
 sg13g2_nor3_2 _5646_ (.A(net1176),
    .B(net1040),
    .C(_1010_),
    .Y(_1778_));
 sg13g2_nand2_1 _5647_ (.Y(_1779_),
    .A(net1522),
    .B(_1778_));
 sg13g2_and2_1 _5648_ (.A(\led_controller.flash.master.sck ),
    .B(_1772_),
    .X(_1780_));
 sg13g2_nor2_1 _5649_ (.A(_1776_),
    .B(_1780_),
    .Y(_1781_));
 sg13g2_nor4_1 _5650_ (.A(_0805_),
    .B(\led_controller.flash.master.bit_counter[2] ),
    .C(\led_controller.flash.master.bit_counter[1] ),
    .D(\led_controller.flash.master.bit_counter[0] ),
    .Y(_1782_));
 sg13g2_nand2_1 _5651_ (.Y(_1783_),
    .A(_1772_),
    .B(_1782_));
 sg13g2_o21ai_1 _5652_ (.B1(_1772_),
    .Y(_1784_),
    .A1(net1333),
    .A2(_1782_));
 sg13g2_nor2b_2 _5653_ (.A(_1776_),
    .B_N(_1784_),
    .Y(_1785_));
 sg13g2_nand2_1 _5654_ (.Y(_1786_),
    .A(_1781_),
    .B(_1783_));
 sg13g2_a221oi_1 _5655_ (.B2(\led_controller.flash.master.tx_data[0] ),
    .C1(net895),
    .B1(_1780_),
    .A1(\led_controller.flash.master.i_tx_data[1] ),
    .Y(_1787_),
    .A2(net967));
 sg13g2_o21ai_1 _5656_ (.B1(net1054),
    .Y(_1788_),
    .A1(\led_controller.flash.master.tx_data[1] ),
    .A2(_1786_));
 sg13g2_o21ai_1 _5657_ (.B1(net1523),
    .Y(_0270_),
    .A1(_1787_),
    .A2(_1788_));
 sg13g2_a22oi_1 _5658_ (.Y(_1789_),
    .B1(_1780_),
    .B2(\led_controller.flash.master.tx_data[1] ),
    .A2(net967),
    .A1(net1610));
 sg13g2_or2_1 _5659_ (.X(_1790_),
    .B(_1789_),
    .A(_1785_));
 sg13g2_a22oi_1 _5660_ (.Y(_1791_),
    .B1(_1785_),
    .B2(net1945),
    .A2(_1776_),
    .A1(\led_controller.flash.master.i_tx_data[1] ));
 sg13g2_a21oi_1 _5661_ (.A1(_1790_),
    .A2(net1946),
    .Y(_0271_),
    .B1(net1040));
 sg13g2_nand2_1 _5662_ (.Y(_1792_),
    .A(net1610),
    .B(_1778_));
 sg13g2_a221oi_1 _5663_ (.B2(\led_controller.flash.master.tx_data[2] ),
    .C1(_1785_),
    .B1(_1780_),
    .A1(\led_controller.flash.master.i_tx_data[3] ),
    .Y(_1793_),
    .A2(net967));
 sg13g2_o21ai_1 _5664_ (.B1(net1055),
    .Y(_1794_),
    .A1(\led_controller.flash.master.tx_data[3] ),
    .A2(_1786_));
 sg13g2_o21ai_1 _5665_ (.B1(_1792_),
    .Y(_0272_),
    .A1(_1793_),
    .A2(_1794_));
 sg13g2_a22oi_1 _5666_ (.Y(_1795_),
    .B1(_1780_),
    .B2(\led_controller.flash.master.tx_data[3] ),
    .A2(net967),
    .A1(\led_controller.flash.master.i_tx_data[4] ));
 sg13g2_or2_1 _5667_ (.X(_1796_),
    .B(_1795_),
    .A(net895));
 sg13g2_a22oi_1 _5668_ (.Y(_1797_),
    .B1(net895),
    .B2(net1892),
    .A2(_1776_),
    .A1(\led_controller.flash.master.i_tx_data[3] ));
 sg13g2_a21oi_1 _5669_ (.A1(_1796_),
    .A2(net1893),
    .Y(_0273_),
    .B1(net1040));
 sg13g2_a22oi_1 _5670_ (.Y(_1798_),
    .B1(_1780_),
    .B2(net1892),
    .A2(net967),
    .A1(net1584));
 sg13g2_or2_1 _5671_ (.X(_1799_),
    .B(_1798_),
    .A(net895));
 sg13g2_a22oi_1 _5672_ (.Y(_1800_),
    .B1(net895),
    .B2(net1980),
    .A2(_1776_),
    .A1(\led_controller.flash.master.i_tx_data[4] ));
 sg13g2_a21oi_1 _5673_ (.A1(_1799_),
    .A2(net1981),
    .Y(_0274_),
    .B1(net1040));
 sg13g2_nand2_1 _5674_ (.Y(_1801_),
    .A(net1584),
    .B(_1778_));
 sg13g2_a221oi_1 _5675_ (.B2(\led_controller.flash.master.tx_data[5] ),
    .C1(net895),
    .B1(_1780_),
    .A1(\led_controller.flash.master.i_tx_data[6] ),
    .Y(_1802_),
    .A2(net967));
 sg13g2_o21ai_1 _5676_ (.B1(net1055),
    .Y(_1803_),
    .A1(\led_controller.flash.master.tx_data[6] ),
    .A2(_1786_));
 sg13g2_o21ai_1 _5677_ (.B1(net1585),
    .Y(_0275_),
    .A1(_1802_),
    .A2(_1803_));
 sg13g2_a22oi_1 _5678_ (.Y(_1804_),
    .B1(_1780_),
    .B2(\led_controller.flash.master.tx_data[6] ),
    .A2(net968),
    .A1(\led_controller.flash.master.i_tx_data[7] ));
 sg13g2_or2_1 _5679_ (.X(_1805_),
    .B(_1804_),
    .A(net895));
 sg13g2_a22oi_1 _5680_ (.Y(_1806_),
    .B1(net895),
    .B2(net1938),
    .A2(_1776_),
    .A1(\led_controller.flash.master.i_tx_data[6] ));
 sg13g2_a21oi_1 _5681_ (.A1(_1805_),
    .A2(net1939),
    .Y(_0276_),
    .B1(net1040));
 sg13g2_o21ai_1 _5682_ (.B1(net1098),
    .Y(_1807_),
    .A1(\led_controller.cpu.led_write_pending ),
    .A2(net2066));
 sg13g2_nor2_1 _5683_ (.A(net1035),
    .B(net2067),
    .Y(_0277_));
 sg13g2_nand2_2 _5684_ (.Y(_1808_),
    .A(\led_controller.cpu.led_write_pending ),
    .B(net1098));
 sg13g2_o21ai_1 _5685_ (.B1(net1059),
    .Y(_1809_),
    .A1(\led_controller.cpu.led_write_color[0] ),
    .A2(_1808_));
 sg13g2_a21oi_1 _5686_ (.A1(_0872_),
    .A2(_1808_),
    .Y(_0278_),
    .B1(_1809_));
 sg13g2_o21ai_1 _5687_ (.B1(net1060),
    .Y(_1810_),
    .A1(\led_controller.cpu.led_write_color[1] ),
    .A2(_1808_));
 sg13g2_a21oi_1 _5688_ (.A1(_0871_),
    .A2(_1808_),
    .Y(_0279_),
    .B1(_1810_));
 sg13g2_nor2_1 _5689_ (.A(_0870_),
    .B(\led_controller.cpu.o_led_strb ),
    .Y(_1811_));
 sg13g2_a221oi_1 _5690_ (.B2(net1098),
    .C1(net1035),
    .B1(_1811_),
    .A1(_0870_),
    .Y(_0280_),
    .A2(_1808_));
 sg13g2_a22oi_1 _5691_ (.Y(_1812_),
    .B1(_1087_),
    .B2(\led_controller.cpu.led_write_strb ),
    .A2(_0917_),
    .A1(net2138));
 sg13g2_nor2_1 _5692_ (.A(net1034),
    .B(net2139),
    .Y(_0281_));
 sg13g2_and2_1 _5693_ (.A(\led_controller.cpu.current_instruction[12] ),
    .B(_1061_),
    .X(_1813_));
 sg13g2_nor2_2 _5694_ (.A(\led_controller.cpu.current_instruction[9] ),
    .B(\led_controller.cpu.current_instruction[8] ),
    .Y(_1814_));
 sg13g2_nor2_2 _5695_ (.A(\led_controller.cpu.current_instruction[11] ),
    .B(\led_controller.cpu.current_instruction[10] ),
    .Y(_1815_));
 sg13g2_and3_2 _5696_ (.X(_1816_),
    .A(_1813_),
    .B(_1814_),
    .C(_1815_));
 sg13g2_and2_1 _5697_ (.A(_1098_),
    .B(_1816_),
    .X(_1817_));
 sg13g2_nor2b_1 _5698_ (.A(_1817_),
    .B_N(net2369),
    .Y(_1818_));
 sg13g2_nor2_1 _5699_ (.A(_0844_),
    .B(_0845_),
    .Y(_1819_));
 sg13g2_o21ai_1 _5700_ (.B1(\led_controller.cpu.current_instruction[11] ),
    .Y(_1820_),
    .A1(\led_controller.cpu.current_instruction[10] ),
    .A2(\led_controller.cpu.current_instruction[9] ));
 sg13g2_nor2_2 _5701_ (.A(_1063_),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_nand2b_1 _5702_ (.Y(_1822_),
    .B(_1062_),
    .A_N(_1820_));
 sg13g2_nand2_1 _5703_ (.Y(_1823_),
    .A(\led_controller.cpu.current_instruction[0] ),
    .B(net981));
 sg13g2_mux4_1 _5704_ (.S0(net1207),
    .A0(\led_controller.cpu.scratch_memory[0][0] ),
    .A1(\led_controller.cpu.scratch_memory[1][0] ),
    .A2(\led_controller.cpu.scratch_memory[2][0] ),
    .A3(\led_controller.cpu.scratch_memory[3][0] ),
    .S1(net1198),
    .X(_1824_));
 sg13g2_and2_1 _5705_ (.A(net1099),
    .B(_1824_),
    .X(_1825_));
 sg13g2_nand2b_1 _5706_ (.Y(_1826_),
    .B(\led_controller.cpu.scratch_memory[4][0] ),
    .A_N(net1212));
 sg13g2_a21oi_1 _5707_ (.A1(net1215),
    .A2(\led_controller.cpu.scratch_memory[5][0] ),
    .Y(_1827_),
    .B1(net1201));
 sg13g2_nor2b_1 _5708_ (.A(net1215),
    .B_N(\led_controller.cpu.scratch_memory[6][0] ),
    .Y(_1828_));
 sg13g2_a21oi_1 _5709_ (.A1(net1215),
    .A2(\led_controller.cpu.scratch_memory[7][0] ),
    .Y(_1829_),
    .B1(_1828_));
 sg13g2_a221oi_1 _5710_ (.B2(net1201),
    .C1(net1101),
    .B1(_1829_),
    .A1(_1826_),
    .Y(_1830_),
    .A2(_1827_));
 sg13g2_or3_1 _5711_ (.A(net1195),
    .B(_1825_),
    .C(_1830_),
    .X(_1831_));
 sg13g2_mux4_1 _5712_ (.S0(net1213),
    .A0(\led_controller.cpu.scratch_memory[8][0] ),
    .A1(\led_controller.cpu.scratch_memory[9][0] ),
    .A2(\led_controller.cpu.scratch_memory[10][0] ),
    .A3(\led_controller.cpu.scratch_memory[11][0] ),
    .S1(net1204),
    .X(_1832_));
 sg13g2_nand2b_1 _5713_ (.Y(_1833_),
    .B(\led_controller.cpu.scratch_memory[12][0] ),
    .A_N(net1217));
 sg13g2_a21oi_1 _5714_ (.A1(net1217),
    .A2(\led_controller.cpu.scratch_memory[13][0] ),
    .Y(_1834_),
    .B1(net1203));
 sg13g2_nand2b_1 _5715_ (.Y(_1835_),
    .B(\led_controller.cpu.scratch_memory[14][0] ),
    .A_N(net1218));
 sg13g2_nand2_1 _5716_ (.Y(_1836_),
    .A(net1218),
    .B(\led_controller.cpu.scratch_memory[15][0] ));
 sg13g2_nand3_1 _5717_ (.B(_1835_),
    .C(_1836_),
    .A(net1203),
    .Y(_1837_));
 sg13g2_a21oi_1 _5718_ (.A1(_1833_),
    .A2(_1834_),
    .Y(_1838_),
    .B1(net1100));
 sg13g2_a221oi_1 _5719_ (.B2(_1838_),
    .C1(_0895_),
    .B1(_1837_),
    .A1(net1100),
    .Y(_1839_),
    .A2(_1832_));
 sg13g2_nor2_1 _5720_ (.A(_1060_),
    .B(_1839_),
    .Y(_1840_));
 sg13g2_and4_1 _5721_ (.A(_0850_),
    .B(_0851_),
    .C(_1054_),
    .D(_1057_),
    .X(_1841_));
 sg13g2_and2_1 _5722_ (.A(_1052_),
    .B(_1841_),
    .X(_1842_));
 sg13g2_nand2_1 _5723_ (.Y(_1843_),
    .A(_1052_),
    .B(_1841_));
 sg13g2_and2_1 _5724_ (.A(_1124_),
    .B(_1841_),
    .X(_1844_));
 sg13g2_a221oi_1 _5725_ (.B2(\led_controller.cpu.i_num_colors[0] ),
    .C1(_1842_),
    .B1(_1844_),
    .A1(_1831_),
    .Y(_1845_),
    .A2(_1840_));
 sg13g2_o21ai_1 _5726_ (.B1(_1821_),
    .Y(_1846_),
    .A1(\led_controller.cpu.i_num_leds[0] ),
    .A2(_1843_));
 sg13g2_nor2_1 _5727_ (.A(_1845_),
    .B(_1846_),
    .Y(_1847_));
 sg13g2_a21oi_2 _5728_ (.B1(_1847_),
    .Y(_1848_),
    .A2(net981),
    .A1(\led_controller.cpu.current_instruction[0] ));
 sg13g2_o21ai_1 _5729_ (.B1(_1823_),
    .Y(_1849_),
    .A1(_1845_),
    .A2(_1846_));
 sg13g2_nor2_2 _5730_ (.A(_0846_),
    .B(\led_controller.cpu.current_instruction[8] ),
    .Y(_1850_));
 sg13g2_a21oi_1 _5731_ (.A1(_1815_),
    .A2(_1850_),
    .Y(_1851_),
    .B1(\led_controller.cpu.status_negative ));
 sg13g2_nor2_2 _5732_ (.A(\led_controller.cpu.current_instruction[9] ),
    .B(_0847_),
    .Y(_1852_));
 sg13g2_nand2_1 _5733_ (.Y(_1853_),
    .A(_1815_),
    .B(_1852_));
 sg13g2_a21oi_1 _5734_ (.A1(\led_controller.cpu.status_negative ),
    .A2(_1853_),
    .Y(_1854_),
    .B1(_1851_));
 sg13g2_nor2_2 _5735_ (.A(_0844_),
    .B(\led_controller.cpu.current_instruction[10] ),
    .Y(_1855_));
 sg13g2_a21oi_1 _5736_ (.A1(_1814_),
    .A2(_1855_),
    .Y(_1856_),
    .B1(_0858_));
 sg13g2_nor2_2 _5737_ (.A(_0846_),
    .B(_0847_),
    .Y(_1857_));
 sg13g2_nor2_2 _5738_ (.A(\led_controller.cpu.current_instruction[11] ),
    .B(_0845_),
    .Y(_1858_));
 sg13g2_a21oi_1 _5739_ (.A1(_1857_),
    .A2(_1858_),
    .Y(_1859_),
    .B1(\led_controller.cpu.status_zero ));
 sg13g2_nor3_1 _5740_ (.A(_1063_),
    .B(_1856_),
    .C(_1859_),
    .Y(_1860_));
 sg13g2_a21oi_2 _5741_ (.B1(_1860_),
    .Y(_1861_),
    .A2(_1854_),
    .A1(_1813_));
 sg13g2_a21o_2 _5742_ (.A2(_1854_),
    .A1(_1813_),
    .B1(_1860_),
    .X(_1862_));
 sg13g2_nor2_1 _5743_ (.A(_1816_),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_nor3_1 _5744_ (.A(net875),
    .B(_1848_),
    .C(_1863_),
    .Y(_1864_));
 sg13g2_o21ai_1 _5745_ (.B1(net1045),
    .Y(_1865_),
    .A1(_1818_),
    .A2(_1864_));
 sg13g2_a21oi_1 _5746_ (.A1(_1818_),
    .A2(_1864_),
    .Y(_0282_),
    .B1(_1865_));
 sg13g2_nand2_1 _5747_ (.Y(_1866_),
    .A(\led_controller.cpu.current_instruction[1] ),
    .B(net981));
 sg13g2_mux4_1 _5748_ (.S0(net1207),
    .A0(\led_controller.cpu.scratch_memory[0][1] ),
    .A1(\led_controller.cpu.scratch_memory[1][1] ),
    .A2(\led_controller.cpu.scratch_memory[2][1] ),
    .A3(\led_controller.cpu.scratch_memory[3][1] ),
    .S1(net1197),
    .X(_1867_));
 sg13g2_nand2b_1 _5749_ (.Y(_1868_),
    .B(\led_controller.cpu.scratch_memory[4][1] ),
    .A_N(net1208));
 sg13g2_a21oi_1 _5750_ (.A1(net1209),
    .A2(\led_controller.cpu.scratch_memory[5][1] ),
    .Y(_1869_),
    .B1(net1199));
 sg13g2_nand2b_1 _5751_ (.Y(_1870_),
    .B(\led_controller.cpu.scratch_memory[6][1] ),
    .A_N(net1209));
 sg13g2_nand2_1 _5752_ (.Y(_1871_),
    .A(net1209),
    .B(\led_controller.cpu.scratch_memory[7][1] ));
 sg13g2_nand3_1 _5753_ (.B(_1870_),
    .C(_1871_),
    .A(net1199),
    .Y(_1872_));
 sg13g2_a21oi_1 _5754_ (.A1(_1868_),
    .A2(_1869_),
    .Y(_1873_),
    .B1(net1099));
 sg13g2_a221oi_1 _5755_ (.B2(_1873_),
    .C1(net1195),
    .B1(_1872_),
    .A1(net1099),
    .Y(_1874_),
    .A2(_1867_));
 sg13g2_mux4_1 _5756_ (.S0(net1210),
    .A0(\led_controller.cpu.scratch_memory[8][1] ),
    .A1(\led_controller.cpu.scratch_memory[9][1] ),
    .A2(\led_controller.cpu.scratch_memory[10][1] ),
    .A3(\led_controller.cpu.scratch_memory[11][1] ),
    .S1(net1200),
    .X(_1875_));
 sg13g2_nand2_1 _5757_ (.Y(_1876_),
    .A(net1102),
    .B(_1875_));
 sg13g2_nand2b_1 _5758_ (.Y(_1877_),
    .B(\led_controller.cpu.scratch_memory[12][1] ),
    .A_N(net1219));
 sg13g2_a21oi_1 _5759_ (.A1(net1219),
    .A2(\led_controller.cpu.scratch_memory[13][1] ),
    .Y(_1878_),
    .B1(net1203));
 sg13g2_nor2b_1 _5760_ (.A(net1220),
    .B_N(\led_controller.cpu.scratch_memory[14][1] ),
    .Y(_1879_));
 sg13g2_a21oi_1 _5761_ (.A1(net1220),
    .A2(\led_controller.cpu.scratch_memory[15][1] ),
    .Y(_1880_),
    .B1(_1879_));
 sg13g2_a221oi_1 _5762_ (.B2(net1203),
    .C1(net1100),
    .B1(_1880_),
    .A1(_1877_),
    .Y(_1881_),
    .A2(_1878_));
 sg13g2_nand3b_1 _5763_ (.B(net1195),
    .C(_1876_),
    .Y(_1882_),
    .A_N(_1881_));
 sg13g2_nor2_1 _5764_ (.A(_1060_),
    .B(_1874_),
    .Y(_1883_));
 sg13g2_a221oi_1 _5765_ (.B2(_1883_),
    .C1(_1842_),
    .B1(_1882_),
    .A1(\led_controller.cpu.i_num_colors[1] ),
    .Y(_1884_),
    .A2(_1844_));
 sg13g2_o21ai_1 _5766_ (.B1(_1821_),
    .Y(_1885_),
    .A1(\led_controller.cpu.i_num_leds[1] ),
    .A2(_1843_));
 sg13g2_o21ai_1 _5767_ (.B1(_1866_),
    .Y(_1886_),
    .A1(_1884_),
    .A2(_1885_));
 sg13g2_inv_2 _5768_ (.Y(_1887_),
    .A(_1886_));
 sg13g2_a22oi_1 _5769_ (.Y(_1888_),
    .B1(_1817_),
    .B2(_1886_),
    .A2(net875),
    .A1(net1186));
 sg13g2_nand2_1 _5770_ (.Y(_1889_),
    .A(\led_controller.cpu.pc[0] ),
    .B(_1849_));
 sg13g2_nand2b_1 _5771_ (.Y(_1890_),
    .B(_1886_),
    .A_N(net1186));
 sg13g2_xor2_1 _5772_ (.B(_1886_),
    .A(net1186),
    .X(_1891_));
 sg13g2_xnor2_1 _5773_ (.Y(_1892_),
    .A(_1889_),
    .B(_1891_));
 sg13g2_nand2_1 _5774_ (.Y(_1893_),
    .A(_1862_),
    .B(_1892_));
 sg13g2_nand2_1 _5775_ (.Y(_1894_),
    .A(net1186),
    .B(net894));
 sg13g2_nand2b_2 _5776_ (.Y(_1895_),
    .B(_1098_),
    .A_N(_1816_));
 sg13g2_nor2_2 _5777_ (.A(net875),
    .B(_1816_),
    .Y(_1896_));
 sg13g2_nand3_1 _5778_ (.B(_1894_),
    .C(_1896_),
    .A(_1893_),
    .Y(_1897_));
 sg13g2_a21oi_1 _5779_ (.A1(_1888_),
    .A2(_1897_),
    .Y(_0283_),
    .B1(net1027));
 sg13g2_nand2b_1 _5780_ (.Y(_1898_),
    .B(\led_controller.cpu.scratch_memory[8][2] ),
    .A_N(net1213));
 sg13g2_a21oi_1 _5781_ (.A1(net1214),
    .A2(\led_controller.cpu.scratch_memory[9][2] ),
    .Y(_1899_),
    .B1(net1204));
 sg13g2_nor2b_1 _5782_ (.A(net1213),
    .B_N(\led_controller.cpu.scratch_memory[10][2] ),
    .Y(_1900_));
 sg13g2_a21oi_1 _5783_ (.A1(net1213),
    .A2(\led_controller.cpu.scratch_memory[11][2] ),
    .Y(_1901_),
    .B1(_1900_));
 sg13g2_a221oi_1 _5784_ (.B2(net1204),
    .C1(net1196),
    .B1(_1901_),
    .A1(_1898_),
    .Y(_1902_),
    .A2(_1899_));
 sg13g2_nand2b_1 _5785_ (.Y(_1903_),
    .B(\led_controller.cpu.scratch_memory[12][2] ),
    .A_N(net1219));
 sg13g2_a21oi_1 _5786_ (.A1(net1215),
    .A2(\led_controller.cpu.scratch_memory[13][2] ),
    .Y(_1904_),
    .B1(net1202));
 sg13g2_nor2b_1 _5787_ (.A(net1219),
    .B_N(\led_controller.cpu.scratch_memory[14][2] ),
    .Y(_1905_));
 sg13g2_a21oi_1 _5788_ (.A1(net1219),
    .A2(\led_controller.cpu.scratch_memory[15][2] ),
    .Y(_1906_),
    .B1(_1905_));
 sg13g2_a221oi_1 _5789_ (.B2(net1203),
    .C1(net1100),
    .B1(_1906_),
    .A1(_1903_),
    .Y(_1907_),
    .A2(_1904_));
 sg13g2_nor3_1 _5790_ (.A(_0895_),
    .B(_1902_),
    .C(_1907_),
    .Y(_1908_));
 sg13g2_mux4_1 _5791_ (.S0(net1207),
    .A0(\led_controller.cpu.scratch_memory[0][2] ),
    .A1(\led_controller.cpu.scratch_memory[1][2] ),
    .A2(\led_controller.cpu.scratch_memory[2][2] ),
    .A3(\led_controller.cpu.scratch_memory[3][2] ),
    .S1(net1197),
    .X(_1909_));
 sg13g2_a21oi_1 _5792_ (.A1(net1208),
    .A2(\led_controller.cpu.scratch_memory[5][2] ),
    .Y(_1910_),
    .B1(net1199));
 sg13g2_o21ai_1 _5793_ (.B1(_1910_),
    .Y(_1911_),
    .A1(net1209),
    .A2(_0896_));
 sg13g2_nor2b_1 _5794_ (.A(net1216),
    .B_N(\led_controller.cpu.scratch_memory[6][2] ),
    .Y(_1912_));
 sg13g2_a21oi_1 _5795_ (.A1(net1216),
    .A2(\led_controller.cpu.scratch_memory[7][2] ),
    .Y(_1913_),
    .B1(_1912_));
 sg13g2_a21oi_1 _5796_ (.A1(net1200),
    .A2(_1913_),
    .Y(_1914_),
    .B1(net1099));
 sg13g2_a221oi_1 _5797_ (.B2(_1914_),
    .C1(net1195),
    .B1(_1911_),
    .A1(net1099),
    .Y(_1915_),
    .A2(_1909_));
 sg13g2_or3_1 _5798_ (.A(_1060_),
    .B(_1908_),
    .C(_1915_),
    .X(_1916_));
 sg13g2_a21oi_1 _5799_ (.A1(\led_controller.cpu.i_num_leds[2] ),
    .A2(_1842_),
    .Y(_1917_),
    .B1(net981));
 sg13g2_a22oi_1 _5800_ (.Y(_1918_),
    .B1(_1916_),
    .B2(_1917_),
    .A2(net981),
    .A1(_0853_));
 sg13g2_a22oi_1 _5801_ (.Y(_1919_),
    .B1(_1817_),
    .B2(net870),
    .A2(_1095_),
    .A1(net2351));
 sg13g2_xnor2_1 _5802_ (.Y(_1920_),
    .A(\led_controller.cpu.pc[2] ),
    .B(net1186));
 sg13g2_inv_1 _5803_ (.Y(_1921_),
    .A(_1920_));
 sg13g2_and2_1 _5804_ (.A(net870),
    .B(_1921_),
    .X(_1922_));
 sg13g2_nand2b_1 _5805_ (.Y(_1923_),
    .B(_1920_),
    .A_N(net870));
 sg13g2_nor2b_1 _5806_ (.A(_1922_),
    .B_N(_1923_),
    .Y(_1924_));
 sg13g2_o21ai_1 _5807_ (.B1(_1890_),
    .Y(_1925_),
    .A1(_1889_),
    .A2(_1891_));
 sg13g2_xnor2_1 _5808_ (.Y(_1926_),
    .A(_1924_),
    .B(_1925_));
 sg13g2_a21oi_1 _5809_ (.A1(_1862_),
    .A2(_1926_),
    .Y(_1927_),
    .B1(net846));
 sg13g2_o21ai_1 _5810_ (.B1(_1927_),
    .Y(_1928_),
    .A1(_1862_),
    .A2(_1921_));
 sg13g2_a21oi_1 _5811_ (.A1(_1919_),
    .A2(_1928_),
    .Y(_0284_),
    .B1(net1028));
 sg13g2_nand2b_1 _5812_ (.Y(_1929_),
    .B(\led_controller.cpu.scratch_memory[0][3] ),
    .A_N(net1208));
 sg13g2_a21oi_1 _5813_ (.A1(net1208),
    .A2(\led_controller.cpu.scratch_memory[1][3] ),
    .Y(_1930_),
    .B1(net1197));
 sg13g2_nor2b_1 _5814_ (.A(net1206),
    .B_N(\led_controller.cpu.scratch_memory[2][3] ),
    .Y(_1931_));
 sg13g2_a21oi_1 _5815_ (.A1(net1206),
    .A2(\led_controller.cpu.scratch_memory[3][3] ),
    .Y(_1932_),
    .B1(_1931_));
 sg13g2_a221oi_1 _5816_ (.B2(net1197),
    .C1(net1196),
    .B1(_1932_),
    .A1(_1929_),
    .Y(_1933_),
    .A2(_1930_));
 sg13g2_nand2b_1 _5817_ (.Y(_1934_),
    .B(\led_controller.cpu.scratch_memory[4][3] ),
    .A_N(net1211));
 sg13g2_a21oi_1 _5818_ (.A1(net1211),
    .A2(\led_controller.cpu.scratch_memory[5][3] ),
    .Y(_1935_),
    .B1(net1199));
 sg13g2_nor2b_1 _5819_ (.A(net1211),
    .B_N(\led_controller.cpu.scratch_memory[6][3] ),
    .Y(_1936_));
 sg13g2_a21oi_1 _5820_ (.A1(net1211),
    .A2(\led_controller.cpu.scratch_memory[7][3] ),
    .Y(_1937_),
    .B1(_1936_));
 sg13g2_a221oi_1 _5821_ (.B2(net1199),
    .C1(net1099),
    .B1(_1937_),
    .A1(_1934_),
    .Y(_1938_),
    .A2(_1935_));
 sg13g2_nor3_1 _5822_ (.A(net1195),
    .B(_1933_),
    .C(_1938_),
    .Y(_1939_));
 sg13g2_nand2b_1 _5823_ (.Y(_1940_),
    .B(\led_controller.cpu.scratch_memory[8][3] ),
    .A_N(net1213));
 sg13g2_a21oi_1 _5824_ (.A1(net1214),
    .A2(\led_controller.cpu.scratch_memory[9][3] ),
    .Y(_1941_),
    .B1(net1204));
 sg13g2_nor2b_1 _5825_ (.A(net1213),
    .B_N(\led_controller.cpu.scratch_memory[10][3] ),
    .Y(_1942_));
 sg13g2_a21oi_1 _5826_ (.A1(net1213),
    .A2(\led_controller.cpu.scratch_memory[11][3] ),
    .Y(_1943_),
    .B1(_1942_));
 sg13g2_a221oi_1 _5827_ (.B2(net1204),
    .C1(net1196),
    .B1(_1943_),
    .A1(_1940_),
    .Y(_1944_),
    .A2(_1941_));
 sg13g2_nand2b_1 _5828_ (.Y(_1945_),
    .B(\led_controller.cpu.scratch_memory[12][3] ),
    .A_N(net1217));
 sg13g2_a21oi_1 _5829_ (.A1(net1217),
    .A2(\led_controller.cpu.scratch_memory[13][3] ),
    .Y(_1946_),
    .B1(net1201));
 sg13g2_nor2b_1 _5830_ (.A(net1217),
    .B_N(\led_controller.cpu.scratch_memory[14][3] ),
    .Y(_1947_));
 sg13g2_a21oi_1 _5831_ (.A1(net1217),
    .A2(\led_controller.cpu.scratch_memory[15][3] ),
    .Y(_1948_),
    .B1(_1947_));
 sg13g2_a221oi_1 _5832_ (.B2(net1204),
    .C1(net1100),
    .B1(_1948_),
    .A1(_1945_),
    .Y(_1949_),
    .A2(_1946_));
 sg13g2_nor3_1 _5833_ (.A(_0895_),
    .B(_1944_),
    .C(_1949_),
    .Y(_1950_));
 sg13g2_or3_1 _5834_ (.A(_1060_),
    .B(_1939_),
    .C(_1950_),
    .X(_1951_));
 sg13g2_a21oi_1 _5835_ (.A1(\led_controller.cpu.i_num_leds[3] ),
    .A2(_1842_),
    .Y(_1952_),
    .B1(net981));
 sg13g2_a22oi_1 _5836_ (.Y(_1953_),
    .B1(_1951_),
    .B2(_1952_),
    .A2(net982),
    .A1(_0852_));
 sg13g2_nand2_1 _5837_ (.Y(_1954_),
    .A(_1817_),
    .B(net868));
 sg13g2_nand3_1 _5838_ (.B(\led_controller.cpu.pc[2] ),
    .C(net1186),
    .A(\led_controller.cpu.pc[3] ),
    .Y(_1955_));
 sg13g2_a21o_1 _5839_ (.A2(net1186),
    .A1(\led_controller.cpu.pc[2] ),
    .B1(\led_controller.cpu.pc[3] ),
    .X(_1956_));
 sg13g2_nand2_2 _5840_ (.Y(_1957_),
    .A(_1955_),
    .B(_1956_));
 sg13g2_inv_1 _5841_ (.Y(_1958_),
    .A(_1957_));
 sg13g2_nand2b_1 _5842_ (.Y(_1959_),
    .B(_1957_),
    .A_N(net868));
 sg13g2_inv_1 _5843_ (.Y(_1960_),
    .A(_1959_));
 sg13g2_a21oi_1 _5844_ (.A1(_1923_),
    .A2(_1925_),
    .Y(_1961_),
    .B1(_1922_));
 sg13g2_a221oi_1 _5845_ (.B2(_1958_),
    .C1(_1922_),
    .B1(net868),
    .A1(_1924_),
    .Y(_1962_),
    .A2(_1925_));
 sg13g2_xnor2_1 _5846_ (.Y(_1963_),
    .A(net868),
    .B(_1957_));
 sg13g2_a21oi_1 _5847_ (.A1(net894),
    .A2(_1957_),
    .Y(_1964_),
    .B1(net846));
 sg13g2_xnor2_1 _5848_ (.Y(_1965_),
    .A(_1961_),
    .B(_1963_));
 sg13g2_nand2b_1 _5849_ (.Y(_1966_),
    .B(_1862_),
    .A_N(_1965_));
 sg13g2_a22oi_1 _5850_ (.Y(_1967_),
    .B1(_1964_),
    .B2(_1966_),
    .A2(net876),
    .A1(net2352));
 sg13g2_a21oi_1 _5851_ (.A1(_1954_),
    .A2(_1967_),
    .Y(_0285_),
    .B1(net1026));
 sg13g2_nand2b_1 _5852_ (.Y(_1968_),
    .B(\led_controller.cpu.scratch_memory[0][4] ),
    .A_N(net1208));
 sg13g2_a21oi_1 _5853_ (.A1(net1208),
    .A2(\led_controller.cpu.scratch_memory[1][4] ),
    .Y(_1969_),
    .B1(net1197));
 sg13g2_nor2b_1 _5854_ (.A(net1206),
    .B_N(\led_controller.cpu.scratch_memory[2][4] ),
    .Y(_1970_));
 sg13g2_a21oi_1 _5855_ (.A1(net1206),
    .A2(\led_controller.cpu.scratch_memory[3][4] ),
    .Y(_1971_),
    .B1(_1970_));
 sg13g2_a221oi_1 _5856_ (.B2(net1198),
    .C1(net1196),
    .B1(_1971_),
    .A1(_1968_),
    .Y(_1972_),
    .A2(_1969_));
 sg13g2_nand2b_1 _5857_ (.Y(_1973_),
    .B(\led_controller.cpu.scratch_memory[4][4] ),
    .A_N(net1212));
 sg13g2_a21oi_1 _5858_ (.A1(net1212),
    .A2(\led_controller.cpu.scratch_memory[5][4] ),
    .Y(_1974_),
    .B1(net1201));
 sg13g2_nor2b_1 _5859_ (.A(net1216),
    .B_N(\led_controller.cpu.scratch_memory[6][4] ),
    .Y(_1975_));
 sg13g2_a21oi_1 _5860_ (.A1(net1216),
    .A2(\led_controller.cpu.scratch_memory[7][4] ),
    .Y(_1976_),
    .B1(_1975_));
 sg13g2_a221oi_1 _5861_ (.B2(net1201),
    .C1(net1101),
    .B1(_1976_),
    .A1(_1973_),
    .Y(_1977_),
    .A2(_1974_));
 sg13g2_nor2_1 _5862_ (.A(_1972_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_mux4_1 _5863_ (.S0(net1210),
    .A0(\led_controller.cpu.scratch_memory[8][4] ),
    .A1(\led_controller.cpu.scratch_memory[9][4] ),
    .A2(\led_controller.cpu.scratch_memory[10][4] ),
    .A3(\led_controller.cpu.scratch_memory[11][4] ),
    .S1(net1200),
    .X(_1979_));
 sg13g2_nand2_1 _5864_ (.Y(_1980_),
    .A(net1102),
    .B(_1979_));
 sg13g2_a21oi_1 _5865_ (.A1(net1215),
    .A2(\led_controller.cpu.scratch_memory[13][4] ),
    .Y(_1981_),
    .B1(net1202));
 sg13g2_o21ai_1 _5866_ (.B1(_1981_),
    .Y(_1982_),
    .A1(net1219),
    .A2(_0897_));
 sg13g2_nor2b_1 _5867_ (.A(net1220),
    .B_N(\led_controller.cpu.scratch_memory[14][4] ),
    .Y(_1983_));
 sg13g2_a21oi_1 _5868_ (.A1(net1220),
    .A2(\led_controller.cpu.scratch_memory[15][4] ),
    .Y(_1984_),
    .B1(_1983_));
 sg13g2_a21oi_1 _5869_ (.A1(net1203),
    .A2(_1984_),
    .Y(_1985_),
    .B1(net1100));
 sg13g2_a21oi_1 _5870_ (.A1(_1982_),
    .A2(_1985_),
    .Y(_1986_),
    .B1(_0895_));
 sg13g2_a22oi_1 _5871_ (.Y(_1987_),
    .B1(_1980_),
    .B2(_1986_),
    .A2(_1978_),
    .A1(_0895_));
 sg13g2_a221oi_1 _5872_ (.B2(_1059_),
    .C1(net981),
    .B1(_1987_),
    .A1(\led_controller.cpu.i_num_leds[4] ),
    .Y(_1988_),
    .A2(_1842_));
 sg13g2_a21oi_2 _5873_ (.B1(_1988_),
    .Y(_1989_),
    .A2(net982),
    .A1(_0851_));
 sg13g2_a22oi_1 _5874_ (.Y(_1990_),
    .B1(_1817_),
    .B2(net845),
    .A2(_1095_),
    .A1(net2322));
 sg13g2_nor2_2 _5875_ (.A(_0869_),
    .B(_1955_),
    .Y(_1991_));
 sg13g2_xnor2_1 _5876_ (.Y(_1992_),
    .A(_0869_),
    .B(_1955_));
 sg13g2_inv_1 _5877_ (.Y(_1993_),
    .A(_1992_));
 sg13g2_nand2_1 _5878_ (.Y(_1994_),
    .A(net845),
    .B(_1993_));
 sg13g2_xnor2_1 _5879_ (.Y(_1995_),
    .A(net845),
    .B(_1993_));
 sg13g2_o21ai_1 _5880_ (.B1(_1995_),
    .Y(_1996_),
    .A1(_1960_),
    .A2(_1962_));
 sg13g2_or3_1 _5881_ (.A(_1960_),
    .B(_1962_),
    .C(_1995_),
    .X(_1997_));
 sg13g2_a21oi_1 _5882_ (.A1(_1996_),
    .A2(_1997_),
    .Y(_1998_),
    .B1(net894));
 sg13g2_nor2_1 _5883_ (.A(_1862_),
    .B(_1993_),
    .Y(_1999_));
 sg13g2_or3_1 _5884_ (.A(_1895_),
    .B(_1998_),
    .C(_1999_),
    .X(_2000_));
 sg13g2_a21oi_1 _5885_ (.A1(_1990_),
    .A2(_2000_),
    .Y(_0286_),
    .B1(net1026));
 sg13g2_nand2b_1 _5886_ (.Y(_2001_),
    .B(\led_controller.cpu.scratch_memory[0][5] ),
    .A_N(net1207));
 sg13g2_a21oi_1 _5887_ (.A1(net1208),
    .A2(\led_controller.cpu.scratch_memory[1][5] ),
    .Y(_2002_),
    .B1(net1197));
 sg13g2_nor2b_1 _5888_ (.A(net1206),
    .B_N(\led_controller.cpu.scratch_memory[2][5] ),
    .Y(_2003_));
 sg13g2_a21oi_1 _5889_ (.A1(net1206),
    .A2(\led_controller.cpu.scratch_memory[3][5] ),
    .Y(_2004_),
    .B1(_2003_));
 sg13g2_a221oi_1 _5890_ (.B2(net1197),
    .C1(net1196),
    .B1(_2004_),
    .A1(_2001_),
    .Y(_2005_),
    .A2(_2002_));
 sg13g2_nand2b_1 _5891_ (.Y(_2006_),
    .B(\led_controller.cpu.scratch_memory[4][5] ),
    .A_N(net1212));
 sg13g2_a21oi_1 _5892_ (.A1(net1212),
    .A2(\led_controller.cpu.scratch_memory[5][5] ),
    .Y(_2007_),
    .B1(net1201));
 sg13g2_nor2b_1 _5893_ (.A(net1215),
    .B_N(\led_controller.cpu.scratch_memory[6][5] ),
    .Y(_2008_));
 sg13g2_a21oi_1 _5894_ (.A1(net1215),
    .A2(\led_controller.cpu.scratch_memory[7][5] ),
    .Y(_2009_),
    .B1(_2008_));
 sg13g2_a221oi_1 _5895_ (.B2(net1201),
    .C1(net1101),
    .B1(_2009_),
    .A1(_2006_),
    .Y(_2010_),
    .A2(_2007_));
 sg13g2_nor2_1 _5896_ (.A(_2005_),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_mux4_1 _5897_ (.S0(net1213),
    .A0(\led_controller.cpu.scratch_memory[8][5] ),
    .A1(\led_controller.cpu.scratch_memory[9][5] ),
    .A2(\led_controller.cpu.scratch_memory[10][5] ),
    .A3(\led_controller.cpu.scratch_memory[11][5] ),
    .S1(net1200),
    .X(_2012_));
 sg13g2_nand2_1 _5898_ (.Y(_2013_),
    .A(net1102),
    .B(_2012_));
 sg13g2_a21oi_1 _5899_ (.A1(net1215),
    .A2(\led_controller.cpu.scratch_memory[13][5] ),
    .Y(_2014_),
    .B1(net1202));
 sg13g2_o21ai_1 _5900_ (.B1(_2014_),
    .Y(_2015_),
    .A1(net1217),
    .A2(_0898_));
 sg13g2_nor2b_1 _5901_ (.A(net1218),
    .B_N(\led_controller.cpu.scratch_memory[14][5] ),
    .Y(_2016_));
 sg13g2_a21oi_1 _5902_ (.A1(net1217),
    .A2(\led_controller.cpu.scratch_memory[15][5] ),
    .Y(_2017_),
    .B1(_2016_));
 sg13g2_a21oi_1 _5903_ (.A1(net1203),
    .A2(_2017_),
    .Y(_2018_),
    .B1(net1100));
 sg13g2_a21oi_1 _5904_ (.A1(_2015_),
    .A2(_2018_),
    .Y(_2019_),
    .B1(_0895_));
 sg13g2_a22oi_1 _5905_ (.Y(_2020_),
    .B1(_2013_),
    .B2(_2019_),
    .A2(_2011_),
    .A1(_0895_));
 sg13g2_a22oi_1 _5906_ (.Y(_2021_),
    .B1(_2020_),
    .B2(_1059_),
    .A2(_1842_),
    .A1(\led_controller.cpu.i_num_leds[5] ));
 sg13g2_mux2_1 _5907_ (.A0(_0850_),
    .A1(_2021_),
    .S(_1821_),
    .X(_2022_));
 sg13g2_inv_2 _5908_ (.Y(_2023_),
    .A(net844));
 sg13g2_a22oi_1 _5909_ (.Y(_2024_),
    .B1(_1817_),
    .B2(_2023_),
    .A2(_1095_),
    .A1(net2358));
 sg13g2_nand2_1 _5910_ (.Y(_2025_),
    .A(_1994_),
    .B(_1997_));
 sg13g2_xnor2_1 _5911_ (.Y(_2026_),
    .A(\led_controller.cpu.pc[5] ),
    .B(_1991_));
 sg13g2_nand2_1 _5912_ (.Y(_2027_),
    .A(net844),
    .B(_2026_));
 sg13g2_or2_1 _5913_ (.X(_2028_),
    .B(_2026_),
    .A(net844));
 sg13g2_nand2_1 _5914_ (.Y(_2029_),
    .A(_2027_),
    .B(_2028_));
 sg13g2_xnor2_1 _5915_ (.Y(_2030_),
    .A(_2025_),
    .B(_2029_));
 sg13g2_a21oi_1 _5916_ (.A1(net894),
    .A2(_2026_),
    .Y(_2031_),
    .B1(_1895_));
 sg13g2_o21ai_1 _5917_ (.B1(_2031_),
    .Y(_2032_),
    .A1(net894),
    .A2(_2030_));
 sg13g2_a21oi_1 _5918_ (.A1(net2359),
    .A2(_2032_),
    .Y(_0287_),
    .B1(net1024));
 sg13g2_nand2b_1 _5919_ (.Y(_2033_),
    .B(\led_controller.cpu.scratch_memory[0][6] ),
    .A_N(net1207));
 sg13g2_a21oi_1 _5920_ (.A1(net1208),
    .A2(\led_controller.cpu.scratch_memory[1][6] ),
    .Y(_2034_),
    .B1(net1198));
 sg13g2_nor2b_1 _5921_ (.A(net1206),
    .B_N(\led_controller.cpu.scratch_memory[2][6] ),
    .Y(_2035_));
 sg13g2_a21oi_1 _5922_ (.A1(net1206),
    .A2(\led_controller.cpu.scratch_memory[3][6] ),
    .Y(_2036_),
    .B1(_2035_));
 sg13g2_a221oi_1 _5923_ (.B2(net1198),
    .C1(net1196),
    .B1(_2036_),
    .A1(_2033_),
    .Y(_2037_),
    .A2(_2034_));
 sg13g2_nand2b_1 _5924_ (.Y(_2038_),
    .B(\led_controller.cpu.scratch_memory[4][6] ),
    .A_N(net1211));
 sg13g2_a21oi_1 _5925_ (.A1(net1212),
    .A2(\led_controller.cpu.scratch_memory[5][6] ),
    .Y(_2039_),
    .B1(net1201));
 sg13g2_nor2b_1 _5926_ (.A(net1216),
    .B_N(\led_controller.cpu.scratch_memory[6][6] ),
    .Y(_2040_));
 sg13g2_a21oi_1 _5927_ (.A1(net1216),
    .A2(\led_controller.cpu.scratch_memory[7][6] ),
    .Y(_2041_),
    .B1(_2040_));
 sg13g2_a221oi_1 _5928_ (.B2(net1202),
    .C1(net1101),
    .B1(_2041_),
    .A1(_2038_),
    .Y(_2042_),
    .A2(_2039_));
 sg13g2_nor3_1 _5929_ (.A(net1195),
    .B(_2037_),
    .C(_2042_),
    .Y(_2043_));
 sg13g2_mux4_1 _5930_ (.S0(net1214),
    .A0(\led_controller.cpu.scratch_memory[8][6] ),
    .A1(\led_controller.cpu.scratch_memory[9][6] ),
    .A2(\led_controller.cpu.scratch_memory[10][6] ),
    .A3(\led_controller.cpu.scratch_memory[11][6] ),
    .S1(net1204),
    .X(_2044_));
 sg13g2_a21oi_1 _5931_ (.A1(net1219),
    .A2(\led_controller.cpu.scratch_memory[13][6] ),
    .Y(_2045_),
    .B1(net1202));
 sg13g2_o21ai_1 _5932_ (.B1(_2045_),
    .Y(_2046_),
    .A1(net1219),
    .A2(_0899_));
 sg13g2_nor2b_1 _5933_ (.A(net1220),
    .B_N(\led_controller.cpu.scratch_memory[14][6] ),
    .Y(_2047_));
 sg13g2_a21oi_1 _5934_ (.A1(net1220),
    .A2(\led_controller.cpu.scratch_memory[15][6] ),
    .Y(_2048_),
    .B1(_2047_));
 sg13g2_a21oi_1 _5935_ (.A1(net1203),
    .A2(_2048_),
    .Y(_2049_),
    .B1(net1100));
 sg13g2_a221oi_1 _5936_ (.B2(_2049_),
    .C1(_0895_),
    .B1(_2046_),
    .A1(net1101),
    .Y(_2050_),
    .A2(_2044_));
 sg13g2_nor3_1 _5937_ (.A(_1060_),
    .B(_2043_),
    .C(_2050_),
    .Y(_2051_));
 sg13g2_a21oi_1 _5938_ (.A1(\led_controller.cpu.i_num_leds[6] ),
    .A2(_1842_),
    .Y(_2052_),
    .B1(_2051_));
 sg13g2_nand2_1 _5939_ (.Y(_2053_),
    .A(net1443),
    .B(net982));
 sg13g2_o21ai_1 _5940_ (.B1(_2053_),
    .Y(_2054_),
    .A1(net982),
    .A2(_2052_));
 sg13g2_inv_1 _5941_ (.Y(_2055_),
    .A(net843));
 sg13g2_a22oi_1 _5942_ (.Y(_2056_),
    .B1(_1817_),
    .B2(net843),
    .A2(_1095_),
    .A1(net2348));
 sg13g2_nand3_1 _5943_ (.B(\led_controller.cpu.pc[5] ),
    .C(_1991_),
    .A(\led_controller.cpu.pc[6] ),
    .Y(_2057_));
 sg13g2_a21o_1 _5944_ (.A2(_1991_),
    .A1(\led_controller.cpu.pc[5] ),
    .B1(\led_controller.cpu.pc[6] ),
    .X(_2058_));
 sg13g2_nand2_1 _5945_ (.Y(_2059_),
    .A(_2057_),
    .B(_2058_));
 sg13g2_nand3_1 _5946_ (.B(_2057_),
    .C(_2058_),
    .A(net843),
    .Y(_2060_));
 sg13g2_xnor2_1 _5947_ (.Y(_2061_),
    .A(net843),
    .B(_2059_));
 sg13g2_nand3_1 _5948_ (.B(_1997_),
    .C(_2028_),
    .A(_1994_),
    .Y(_2062_));
 sg13g2_a21o_1 _5949_ (.A2(_2062_),
    .A1(_2027_),
    .B1(_2061_),
    .X(_2063_));
 sg13g2_nand3_1 _5950_ (.B(_2061_),
    .C(_2062_),
    .A(_2027_),
    .Y(_2064_));
 sg13g2_a21oi_1 _5951_ (.A1(_2063_),
    .A2(_2064_),
    .Y(_2065_),
    .B1(net894));
 sg13g2_a21oi_1 _5952_ (.A1(_1861_),
    .A2(_2059_),
    .Y(_2066_),
    .B1(_2065_));
 sg13g2_nand2_1 _5953_ (.Y(_2067_),
    .A(_1896_),
    .B(_2066_));
 sg13g2_a21oi_1 _5954_ (.A1(net2349),
    .A2(_2067_),
    .Y(_0288_),
    .B1(net1024));
 sg13g2_mux2_1 _5955_ (.A0(\led_controller.cpu.scratch_memory[12][7] ),
    .A1(\led_controller.cpu.scratch_memory[13][7] ),
    .S(net1211),
    .X(_2068_));
 sg13g2_o21ai_1 _5956_ (.B1(net1205),
    .Y(_2069_),
    .A1(net1218),
    .A2(_0901_));
 sg13g2_a21oi_1 _5957_ (.A1(net1218),
    .A2(\led_controller.cpu.scratch_memory[15][7] ),
    .Y(_2070_),
    .B1(_2069_));
 sg13g2_o21ai_1 _5958_ (.B1(_0002_),
    .Y(_2071_),
    .A1(net1204),
    .A2(_2068_));
 sg13g2_nand2b_1 _5959_ (.Y(_2072_),
    .B(\led_controller.cpu.scratch_memory[8][7] ),
    .A_N(net1210));
 sg13g2_a21oi_1 _5960_ (.A1(net1210),
    .A2(\led_controller.cpu.scratch_memory[9][7] ),
    .Y(_2073_),
    .B1(net1200));
 sg13g2_nor2b_1 _5961_ (.A(net1210),
    .B_N(\led_controller.cpu.scratch_memory[10][7] ),
    .Y(_2074_));
 sg13g2_a21oi_1 _5962_ (.A1(net1210),
    .A2(\led_controller.cpu.scratch_memory[11][7] ),
    .Y(_2075_),
    .B1(_2074_));
 sg13g2_a221oi_1 _5963_ (.B2(net1200),
    .C1(net1196),
    .B1(_2075_),
    .A1(_2072_),
    .Y(_2076_),
    .A2(_2073_));
 sg13g2_o21ai_1 _5964_ (.B1(_0003_),
    .Y(_2077_),
    .A1(_2070_),
    .A2(_2071_));
 sg13g2_mux4_1 _5965_ (.S0(net1207),
    .A0(\led_controller.cpu.scratch_memory[0][7] ),
    .A1(\led_controller.cpu.scratch_memory[1][7] ),
    .A2(\led_controller.cpu.scratch_memory[2][7] ),
    .A3(\led_controller.cpu.scratch_memory[3][7] ),
    .S1(net1197),
    .X(_2078_));
 sg13g2_a21oi_1 _5966_ (.A1(net1209),
    .A2(\led_controller.cpu.scratch_memory[5][7] ),
    .Y(_2079_),
    .B1(net1199));
 sg13g2_o21ai_1 _5967_ (.B1(_2079_),
    .Y(_2080_),
    .A1(net1209),
    .A2(_0900_));
 sg13g2_nor2b_1 _5968_ (.A(net1211),
    .B_N(\led_controller.cpu.scratch_memory[6][7] ),
    .Y(_2081_));
 sg13g2_a21oi_1 _5969_ (.A1(net1211),
    .A2(\led_controller.cpu.scratch_memory[7][7] ),
    .Y(_2082_),
    .B1(_2081_));
 sg13g2_a21oi_1 _5970_ (.A1(net1200),
    .A2(_2082_),
    .Y(_2083_),
    .B1(net1099));
 sg13g2_a221oi_1 _5971_ (.B2(_2083_),
    .C1(net1195),
    .B1(_2080_),
    .A1(net1099),
    .Y(_2084_),
    .A2(_2078_));
 sg13g2_o21ai_1 _5972_ (.B1(_1059_),
    .Y(_2085_),
    .A1(_2076_),
    .A2(_2077_));
 sg13g2_a21oi_1 _5973_ (.A1(\led_controller.cpu.i_num_leds[7] ),
    .A2(_1842_),
    .Y(_2086_),
    .B1(net981));
 sg13g2_o21ai_1 _5974_ (.B1(_2086_),
    .Y(_2087_),
    .A1(_2084_),
    .A2(_2085_));
 sg13g2_o21ai_1 _5975_ (.B1(_2087_),
    .Y(_2088_),
    .A1(\led_controller.cpu.current_instruction[7] ),
    .A2(_1821_));
 sg13g2_inv_1 _5976_ (.Y(_2089_),
    .A(net841));
 sg13g2_a22oi_1 _5977_ (.Y(_2090_),
    .B1(_1817_),
    .B2(_2089_),
    .A2(_1095_),
    .A1(net2363));
 sg13g2_nand4_1 _5978_ (.B(\led_controller.cpu.pc[6] ),
    .C(\led_controller.cpu.pc[5] ),
    .A(\led_controller.cpu.pc[7] ),
    .Y(_2091_),
    .D(_1991_));
 sg13g2_xor2_1 _5979_ (.B(_2057_),
    .A(\led_controller.cpu.pc[7] ),
    .X(_2092_));
 sg13g2_nand2_2 _5980_ (.Y(_2093_),
    .A(net840),
    .B(_2092_));
 sg13g2_or2_1 _5981_ (.X(_2094_),
    .B(_2092_),
    .A(net840));
 sg13g2_nand3_1 _5982_ (.B(_2064_),
    .C(_2094_),
    .A(_2060_),
    .Y(_2095_));
 sg13g2_nor2b_1 _5983_ (.A(_2095_),
    .B_N(_2093_),
    .Y(_2096_));
 sg13g2_a22oi_1 _5984_ (.Y(_2097_),
    .B1(_2093_),
    .B2(_2094_),
    .A2(_2064_),
    .A1(_2060_));
 sg13g2_or2_1 _5985_ (.X(_2098_),
    .B(_2097_),
    .A(net892));
 sg13g2_a21oi_1 _5986_ (.A1(net892),
    .A2(_2092_),
    .Y(_2099_),
    .B1(net846));
 sg13g2_o21ai_1 _5987_ (.B1(_2099_),
    .Y(_2100_),
    .A1(_2096_),
    .A2(_2098_));
 sg13g2_a21oi_1 _5988_ (.A1(_2090_),
    .A2(_2100_),
    .Y(_0289_),
    .B1(net1023));
 sg13g2_nand2_1 _5989_ (.Y(_2101_),
    .A(net1907),
    .B(net874));
 sg13g2_nor2_1 _5990_ (.A(_0867_),
    .B(_2091_),
    .Y(_2102_));
 sg13g2_xnor2_1 _5991_ (.Y(_2103_),
    .A(_0867_),
    .B(_2091_));
 sg13g2_xor2_1 _5992_ (.B(_2103_),
    .A(net839),
    .X(_2104_));
 sg13g2_nand3_1 _5993_ (.B(_2095_),
    .C(_2104_),
    .A(_2093_),
    .Y(_2105_));
 sg13g2_a21o_1 _5994_ (.A2(_2095_),
    .A1(_2093_),
    .B1(_2104_),
    .X(_2106_));
 sg13g2_a21o_1 _5995_ (.A2(_2106_),
    .A1(_2105_),
    .B1(net892),
    .X(_2107_));
 sg13g2_nand2_1 _5996_ (.Y(_2108_),
    .A(net892),
    .B(_2103_));
 sg13g2_nand3_1 _5997_ (.B(_2107_),
    .C(_2108_),
    .A(_1896_),
    .Y(_2109_));
 sg13g2_a21oi_1 _5998_ (.A1(_2101_),
    .A2(_2109_),
    .Y(_0290_),
    .B1(net1026));
 sg13g2_nand2_1 _5999_ (.Y(_2110_),
    .A(net2286),
    .B(net874));
 sg13g2_o21ai_1 _6000_ (.B1(_2105_),
    .Y(_2111_),
    .A1(net839),
    .A2(_2103_));
 sg13g2_xnor2_1 _6001_ (.Y(_2112_),
    .A(\led_controller.cpu.pc[9] ),
    .B(_2102_));
 sg13g2_xor2_1 _6002_ (.B(_2112_),
    .A(net839),
    .X(_2113_));
 sg13g2_xor2_1 _6003_ (.B(_2113_),
    .A(_2111_),
    .X(_2114_));
 sg13g2_a21oi_1 _6004_ (.A1(net892),
    .A2(_2112_),
    .Y(_2115_),
    .B1(net846));
 sg13g2_o21ai_1 _6005_ (.B1(_2115_),
    .Y(_2116_),
    .A1(net892),
    .A2(_2114_));
 sg13g2_a21oi_1 _6006_ (.A1(_2110_),
    .A2(_2116_),
    .Y(_0291_),
    .B1(net1024));
 sg13g2_nand3_1 _6007_ (.B(\led_controller.cpu.pc[9] ),
    .C(_2102_),
    .A(\led_controller.cpu.pc[10] ),
    .Y(_2117_));
 sg13g2_a21o_1 _6008_ (.A2(_2102_),
    .A1(\led_controller.cpu.pc[9] ),
    .B1(\led_controller.cpu.pc[10] ),
    .X(_2118_));
 sg13g2_nand2_1 _6009_ (.Y(_2119_),
    .A(_2117_),
    .B(_2118_));
 sg13g2_or2_1 _6010_ (.X(_2120_),
    .B(_2119_),
    .A(net839));
 sg13g2_xnor2_1 _6011_ (.Y(_2121_),
    .A(net839),
    .B(_2119_));
 sg13g2_a21o_1 _6012_ (.A2(_2112_),
    .A1(_2103_),
    .B1(net839),
    .X(_2122_));
 sg13g2_nand4_1 _6013_ (.B(_2095_),
    .C(_2104_),
    .A(_2093_),
    .Y(_2123_),
    .D(_2113_));
 sg13g2_and2_1 _6014_ (.A(_2122_),
    .B(_2123_),
    .X(_2124_));
 sg13g2_xnor2_1 _6015_ (.Y(_2125_),
    .A(_2121_),
    .B(_2124_));
 sg13g2_nand2_1 _6016_ (.Y(_2126_),
    .A(net892),
    .B(_2119_));
 sg13g2_nand2_1 _6017_ (.Y(_2127_),
    .A(_1896_),
    .B(_2126_));
 sg13g2_a21oi_1 _6018_ (.A1(_1862_),
    .A2(_2125_),
    .Y(_2128_),
    .B1(_2127_));
 sg13g2_a21oi_1 _6019_ (.A1(net2203),
    .A2(net874),
    .Y(_2129_),
    .B1(_2128_));
 sg13g2_nor2_1 _6020_ (.A(net1026),
    .B(_2129_),
    .Y(_0292_));
 sg13g2_nand2_1 _6021_ (.Y(_2130_),
    .A(net2056),
    .B(net874));
 sg13g2_nor2_1 _6022_ (.A(_0866_),
    .B(_2117_),
    .Y(_2131_));
 sg13g2_xnor2_1 _6023_ (.Y(_2132_),
    .A(_0866_),
    .B(_2117_));
 sg13g2_xor2_1 _6024_ (.B(_2132_),
    .A(net839),
    .X(_2133_));
 sg13g2_o21ai_1 _6025_ (.B1(_2120_),
    .Y(_2134_),
    .A1(_2121_),
    .A2(_2124_));
 sg13g2_xor2_1 _6026_ (.B(_2134_),
    .A(_2133_),
    .X(_2135_));
 sg13g2_a21oi_1 _6027_ (.A1(net892),
    .A2(_2132_),
    .Y(_2136_),
    .B1(net846));
 sg13g2_o21ai_1 _6028_ (.B1(_2136_),
    .Y(_2137_),
    .A1(net893),
    .A2(_2135_));
 sg13g2_a21oi_1 _6029_ (.A1(_2130_),
    .A2(_2137_),
    .Y(_0293_),
    .B1(net1026));
 sg13g2_nand2_1 _6030_ (.Y(_2138_),
    .A(net2248),
    .B(net874));
 sg13g2_and2_1 _6031_ (.A(\led_controller.cpu.pc[12] ),
    .B(_2131_),
    .X(_2139_));
 sg13g2_xnor2_1 _6032_ (.Y(_2140_),
    .A(\led_controller.cpu.pc[12] ),
    .B(_2131_));
 sg13g2_nor2_1 _6033_ (.A(net840),
    .B(_2140_),
    .Y(_2141_));
 sg13g2_nand2_1 _6034_ (.Y(_2142_),
    .A(net840),
    .B(_2140_));
 sg13g2_nand2b_1 _6035_ (.Y(_2143_),
    .B(_2142_),
    .A_N(_2141_));
 sg13g2_nand2b_1 _6036_ (.Y(_2144_),
    .B(_2133_),
    .A_N(_2121_));
 sg13g2_o21ai_1 _6037_ (.B1(_2122_),
    .Y(_2145_),
    .A1(net839),
    .A2(_2132_));
 sg13g2_nor2b_1 _6038_ (.A(_2145_),
    .B_N(_2120_),
    .Y(_2146_));
 sg13g2_o21ai_1 _6039_ (.B1(_2146_),
    .Y(_2147_),
    .A1(_2123_),
    .A2(_2144_));
 sg13g2_xnor2_1 _6040_ (.Y(_2148_),
    .A(_2143_),
    .B(_2147_));
 sg13g2_nor2_1 _6041_ (.A(net893),
    .B(_2148_),
    .Y(_2149_));
 sg13g2_a21oi_1 _6042_ (.A1(net893),
    .A2(_2140_),
    .Y(_2150_),
    .B1(_2149_));
 sg13g2_nand2_1 _6043_ (.Y(_2151_),
    .A(_1896_),
    .B(_2150_));
 sg13g2_a21oi_1 _6044_ (.A1(_2138_),
    .A2(_2151_),
    .Y(_0294_),
    .B1(net1023));
 sg13g2_nand2_1 _6045_ (.Y(_2152_),
    .A(net2246),
    .B(net875));
 sg13g2_a21oi_1 _6046_ (.A1(_2142_),
    .A2(_2147_),
    .Y(_2153_),
    .B1(_2141_));
 sg13g2_xnor2_1 _6047_ (.Y(_2154_),
    .A(\led_controller.cpu.pc[13] ),
    .B(_2139_));
 sg13g2_nand2_1 _6048_ (.Y(_2155_),
    .A(net842),
    .B(_2154_));
 sg13g2_or2_1 _6049_ (.X(_2156_),
    .B(_2154_),
    .A(net840));
 sg13g2_nand2_1 _6050_ (.Y(_2157_),
    .A(_2155_),
    .B(_2156_));
 sg13g2_xor2_1 _6051_ (.B(_2157_),
    .A(_2153_),
    .X(_2158_));
 sg13g2_a21oi_1 _6052_ (.A1(net893),
    .A2(_2154_),
    .Y(_2159_),
    .B1(net846));
 sg13g2_o21ai_1 _6053_ (.B1(_2159_),
    .Y(_2160_),
    .A1(net893),
    .A2(_2158_));
 sg13g2_a21oi_1 _6054_ (.A1(_2152_),
    .A2(_2160_),
    .Y(_0295_),
    .B1(net1026));
 sg13g2_nand3_1 _6055_ (.B(\led_controller.cpu.pc[13] ),
    .C(_2139_),
    .A(\led_controller.cpu.pc[14] ),
    .Y(_2161_));
 sg13g2_a21o_1 _6056_ (.A2(_2139_),
    .A1(\led_controller.cpu.pc[13] ),
    .B1(\led_controller.cpu.pc[14] ),
    .X(_2162_));
 sg13g2_nand2_1 _6057_ (.Y(_2163_),
    .A(_2161_),
    .B(_2162_));
 sg13g2_xor2_1 _6058_ (.B(_2163_),
    .A(net841),
    .X(_2164_));
 sg13g2_nand2_1 _6059_ (.Y(_2165_),
    .A(_2153_),
    .B(_2156_));
 sg13g2_a21oi_1 _6060_ (.A1(_2155_),
    .A2(_2165_),
    .Y(_2166_),
    .B1(_2164_));
 sg13g2_nand3_1 _6061_ (.B(_2164_),
    .C(_2165_),
    .A(_2155_),
    .Y(_2167_));
 sg13g2_nand2b_1 _6062_ (.Y(_2168_),
    .B(_2167_),
    .A_N(_2166_));
 sg13g2_nand2_1 _6063_ (.Y(_2169_),
    .A(net893),
    .B(_2163_));
 sg13g2_a21oi_1 _6064_ (.A1(_1862_),
    .A2(_2168_),
    .Y(_2170_),
    .B1(net846));
 sg13g2_a22oi_1 _6065_ (.Y(_2171_),
    .B1(_2169_),
    .B2(_2170_),
    .A2(net875),
    .A1(net2289));
 sg13g2_nor2_1 _6066_ (.A(net1026),
    .B(_2171_),
    .Y(_0296_));
 sg13g2_nand2_1 _6067_ (.Y(_2172_),
    .A(net2060),
    .B(net875));
 sg13g2_o21ai_1 _6068_ (.B1(_2167_),
    .Y(_2173_),
    .A1(net840),
    .A2(_2163_));
 sg13g2_xor2_1 _6069_ (.B(_2161_),
    .A(\led_controller.cpu.pc[15] ),
    .X(_2174_));
 sg13g2_xnor2_1 _6070_ (.Y(_2175_),
    .A(net840),
    .B(_2174_));
 sg13g2_xnor2_1 _6071_ (.Y(_2176_),
    .A(_2173_),
    .B(_2175_));
 sg13g2_a21oi_1 _6072_ (.A1(net893),
    .A2(_2174_),
    .Y(_2177_),
    .B1(net846));
 sg13g2_o21ai_1 _6073_ (.B1(_2177_),
    .Y(_2178_),
    .A1(net893),
    .A2(_2176_));
 sg13g2_a21oi_1 _6074_ (.A1(_2172_),
    .A2(_2178_),
    .Y(_0297_),
    .B1(net1026));
 sg13g2_nand3_1 _6075_ (.B(_1814_),
    .C(_1858_),
    .A(_1813_),
    .Y(_2179_));
 sg13g2_nand3_1 _6076_ (.B(_1850_),
    .C(_1858_),
    .A(_1062_),
    .Y(_2180_));
 sg13g2_and2_1 _6077_ (.A(net979),
    .B(net975),
    .X(_2181_));
 sg13g2_nand2_1 _6078_ (.Y(_2182_),
    .A(net978),
    .B(net975));
 sg13g2_a22oi_1 _6079_ (.Y(_2183_),
    .B1(_1855_),
    .B2(_1850_),
    .A2(_1852_),
    .A1(_1815_));
 sg13g2_o21ai_1 _6080_ (.B1(_2181_),
    .Y(_2184_),
    .A1(_1063_),
    .A2(_2183_));
 sg13g2_nand2_1 _6081_ (.Y(_2185_),
    .A(_1094_),
    .B(_2184_));
 sg13g2_nor2b_2 _6082_ (.A(net875),
    .B_N(_2184_),
    .Y(_2186_));
 sg13g2_o21ai_1 _6083_ (.B1(net1046),
    .Y(_2187_),
    .A1(net2231),
    .A2(net838));
 sg13g2_nor2_1 _6084_ (.A(net2231),
    .B(_2181_),
    .Y(_2188_));
 sg13g2_a21oi_1 _6085_ (.A1(_1849_),
    .A2(_2181_),
    .Y(_2189_),
    .B1(_2188_));
 sg13g2_a21oi_1 _6086_ (.A1(net838),
    .A2(_2189_),
    .Y(_0298_),
    .B1(_2187_));
 sg13g2_nor2b_1 _6087_ (.A(_1886_),
    .B_N(net977),
    .Y(_2190_));
 sg13g2_xor2_1 _6088_ (.B(net1185),
    .A(net1184),
    .X(_2191_));
 sg13g2_o21ai_1 _6089_ (.B1(net980),
    .Y(_2192_),
    .A1(net977),
    .A2(_2191_));
 sg13g2_nor2_1 _6090_ (.A(_2190_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_nor2_1 _6091_ (.A(net1184),
    .B(net837),
    .Y(_2194_));
 sg13g2_o21ai_1 _6092_ (.B1(net837),
    .Y(_2195_),
    .A1(net980),
    .A2(_2191_));
 sg13g2_nor2_1 _6093_ (.A(_2193_),
    .B(_2195_),
    .Y(_2196_));
 sg13g2_nor3_1 _6094_ (.A(net1025),
    .B(_2194_),
    .C(_2196_),
    .Y(_0299_));
 sg13g2_and3_2 _6095_ (.X(_2197_),
    .A(net1183),
    .B(net1184),
    .C(net1185));
 sg13g2_a21oi_1 _6096_ (.A1(net1184),
    .A2(net1185),
    .Y(_2198_),
    .B1(net1183));
 sg13g2_o21ai_1 _6097_ (.B1(net978),
    .Y(_2199_),
    .A1(_2197_),
    .A2(_2198_));
 sg13g2_a22oi_1 _6098_ (.Y(_2200_),
    .B1(_2182_),
    .B2(_2199_),
    .A2(net975),
    .A1(net870));
 sg13g2_o21ai_1 _6099_ (.B1(net1183),
    .Y(_2201_),
    .A1(\led_controller.cpu.register_x[1] ),
    .A2(net1185));
 sg13g2_inv_1 _6100_ (.Y(_2202_),
    .A(_2201_));
 sg13g2_nor3_2 _6101_ (.A(net1183),
    .B(net1184),
    .C(net1185),
    .Y(_2203_));
 sg13g2_nor3_1 _6102_ (.A(net978),
    .B(_2202_),
    .C(_2203_),
    .Y(_2204_));
 sg13g2_o21ai_1 _6103_ (.B1(net837),
    .Y(_2205_),
    .A1(_2200_),
    .A2(_2204_));
 sg13g2_o21ai_1 _6104_ (.B1(_2205_),
    .Y(_2206_),
    .A1(net1183),
    .A2(net837));
 sg13g2_nor2_1 _6105_ (.A(net1025),
    .B(_2206_),
    .Y(_0300_));
 sg13g2_xnor2_1 _6106_ (.Y(_2207_),
    .A(\led_controller.cpu.register_x[3] ),
    .B(_2197_));
 sg13g2_nand2_1 _6107_ (.Y(_2208_),
    .A(net978),
    .B(_2207_));
 sg13g2_a22oi_1 _6108_ (.Y(_2209_),
    .B1(_2182_),
    .B2(_2208_),
    .A2(net975),
    .A1(net869));
 sg13g2_xnor2_1 _6109_ (.Y(_2210_),
    .A(_0864_),
    .B(_2203_));
 sg13g2_nor2_1 _6110_ (.A(net978),
    .B(_2210_),
    .Y(_2211_));
 sg13g2_o21ai_1 _6111_ (.B1(net837),
    .Y(_2212_),
    .A1(_2209_),
    .A2(_2211_));
 sg13g2_o21ai_1 _6112_ (.B1(_2212_),
    .Y(_2213_),
    .A1(net2332),
    .A2(net837));
 sg13g2_nor2_1 _6113_ (.A(net1025),
    .B(_2213_),
    .Y(_0301_));
 sg13g2_nand3_1 _6114_ (.B(\led_controller.cpu.register_x[3] ),
    .C(_2197_),
    .A(net1182),
    .Y(_2214_));
 sg13g2_a21o_1 _6115_ (.A2(_2197_),
    .A1(\led_controller.cpu.register_x[3] ),
    .B1(net1182),
    .X(_2215_));
 sg13g2_nand2_1 _6116_ (.Y(_2216_),
    .A(_2214_),
    .B(_2215_));
 sg13g2_o21ai_1 _6117_ (.B1(net978),
    .Y(_2217_),
    .A1(net975),
    .A2(_2216_));
 sg13g2_a21oi_1 _6118_ (.A1(net845),
    .A2(net976),
    .Y(_2218_),
    .B1(_2217_));
 sg13g2_and3_1 _6119_ (.X(_2219_),
    .A(_0863_),
    .B(_0864_),
    .C(_2203_));
 sg13g2_a21oi_1 _6120_ (.A1(_0864_),
    .A2(_2203_),
    .Y(_2220_),
    .B1(_0863_));
 sg13g2_nor3_1 _6121_ (.A(net978),
    .B(_2219_),
    .C(_2220_),
    .Y(_2221_));
 sg13g2_o21ai_1 _6122_ (.B1(net838),
    .Y(_2222_),
    .A1(_2218_),
    .A2(_2221_));
 sg13g2_o21ai_1 _6123_ (.B1(_2222_),
    .Y(_2223_),
    .A1(net1182),
    .A2(net838));
 sg13g2_nor2_1 _6124_ (.A(net1025),
    .B(_2223_),
    .Y(_0302_));
 sg13g2_nand4_1 _6125_ (.B(net1182),
    .C(\led_controller.cpu.register_x[3] ),
    .A(\led_controller.cpu.register_x[5] ),
    .Y(_2224_),
    .D(_2197_));
 sg13g2_xor2_1 _6126_ (.B(_2214_),
    .A(\led_controller.cpu.register_x[5] ),
    .X(_2225_));
 sg13g2_o21ai_1 _6127_ (.B1(net979),
    .Y(_2226_),
    .A1(net976),
    .A2(_2225_));
 sg13g2_a21oi_1 _6128_ (.A1(_2023_),
    .A2(net975),
    .Y(_2227_),
    .B1(_2226_));
 sg13g2_nor2b_1 _6129_ (.A(_2219_),
    .B_N(\led_controller.cpu.register_x[5] ),
    .Y(_2228_));
 sg13g2_nor2b_1 _6130_ (.A(\led_controller.cpu.register_x[5] ),
    .B_N(_2219_),
    .Y(_2229_));
 sg13g2_nor3_1 _6131_ (.A(net978),
    .B(_2228_),
    .C(_2229_),
    .Y(_2230_));
 sg13g2_o21ai_1 _6132_ (.B1(net838),
    .Y(_2231_),
    .A1(_2227_),
    .A2(_2230_));
 sg13g2_o21ai_1 _6133_ (.B1(_2231_),
    .Y(_2232_),
    .A1(net2325),
    .A2(net838));
 sg13g2_nor2_1 _6134_ (.A(net1025),
    .B(_2232_),
    .Y(_0303_));
 sg13g2_nor2_1 _6135_ (.A(_0862_),
    .B(_2224_),
    .Y(_2233_));
 sg13g2_xnor2_1 _6136_ (.Y(_2234_),
    .A(_0862_),
    .B(_2224_));
 sg13g2_o21ai_1 _6137_ (.B1(net979),
    .Y(_2235_),
    .A1(net976),
    .A2(_2234_));
 sg13g2_a21oi_1 _6138_ (.A1(net843),
    .A2(net976),
    .Y(_2236_),
    .B1(_2235_));
 sg13g2_nor2_1 _6139_ (.A(_0862_),
    .B(_2229_),
    .Y(_2237_));
 sg13g2_and2_1 _6140_ (.A(_0862_),
    .B(_2229_),
    .X(_2238_));
 sg13g2_nor3_1 _6141_ (.A(net979),
    .B(_2237_),
    .C(_2238_),
    .Y(_2239_));
 sg13g2_o21ai_1 _6142_ (.B1(net838),
    .Y(_2240_),
    .A1(_2236_),
    .A2(_2239_));
 sg13g2_o21ai_1 _6143_ (.B1(_2240_),
    .Y(_2241_),
    .A1(net2256),
    .A2(net837));
 sg13g2_nor2_1 _6144_ (.A(net1030),
    .B(_2241_),
    .Y(_0304_));
 sg13g2_o21ai_1 _6145_ (.B1(net1046),
    .Y(_2242_),
    .A1(net2337),
    .A2(net837));
 sg13g2_xnor2_1 _6146_ (.Y(_2243_),
    .A(\led_controller.cpu.register_x[7] ),
    .B(_2233_));
 sg13g2_inv_1 _6147_ (.Y(_2244_),
    .A(_2243_));
 sg13g2_o21ai_1 _6148_ (.B1(net979),
    .Y(_2245_),
    .A1(net975),
    .A2(_2244_));
 sg13g2_a21oi_1 _6149_ (.A1(net842),
    .A2(net975),
    .Y(_2246_),
    .B1(_2245_));
 sg13g2_xnor2_1 _6150_ (.Y(_2247_),
    .A(net2337),
    .B(_2238_));
 sg13g2_nor2_1 _6151_ (.A(net979),
    .B(_2247_),
    .Y(_2248_));
 sg13g2_nor3_1 _6152_ (.A(_2185_),
    .B(_2246_),
    .C(_2248_),
    .Y(_2249_));
 sg13g2_nor2_1 _6153_ (.A(_2242_),
    .B(_2249_),
    .Y(_0305_));
 sg13g2_and3_1 _6154_ (.X(_2250_),
    .A(_1813_),
    .B(_1815_),
    .C(_1857_));
 sg13g2_nand3_1 _6155_ (.B(_1815_),
    .C(_1857_),
    .A(_1813_),
    .Y(_2251_));
 sg13g2_and3_2 _6156_ (.X(_2252_),
    .A(_1062_),
    .B(_1852_),
    .C(_1858_));
 sg13g2_nand3_1 _6157_ (.B(_1852_),
    .C(_1858_),
    .A(_1062_),
    .Y(_2253_));
 sg13g2_nor2_1 _6158_ (.A(net974),
    .B(net972),
    .Y(_2254_));
 sg13g2_a22oi_1 _6159_ (.Y(_2255_),
    .B1(_1855_),
    .B2(_1857_),
    .A2(_1850_),
    .A1(_1815_));
 sg13g2_o21ai_1 _6160_ (.B1(_2254_),
    .Y(_2256_),
    .A1(_1063_),
    .A2(_2255_));
 sg13g2_nand2_1 _6161_ (.Y(_2257_),
    .A(_1098_),
    .B(_2256_));
 sg13g2_nor2b_2 _6162_ (.A(net874),
    .B_N(_2256_),
    .Y(_2258_));
 sg13g2_nand2b_1 _6163_ (.Y(_2259_),
    .B(_2256_),
    .A_N(net874));
 sg13g2_o21ai_1 _6164_ (.B1(net1045),
    .Y(_2260_),
    .A1(net1181),
    .A2(_2258_));
 sg13g2_and2_1 _6165_ (.A(_1849_),
    .B(_2254_),
    .X(_2261_));
 sg13g2_nor2_1 _6166_ (.A(net1181),
    .B(_2254_),
    .Y(_2262_));
 sg13g2_nor3_1 _6167_ (.A(_2259_),
    .B(_2261_),
    .C(_2262_),
    .Y(_2263_));
 sg13g2_nor2_1 _6168_ (.A(_2260_),
    .B(_2263_),
    .Y(_0306_));
 sg13g2_xor2_1 _6169_ (.B(net1181),
    .A(net1180),
    .X(_2264_));
 sg13g2_nand2_1 _6170_ (.Y(_2265_),
    .A(_1886_),
    .B(_2253_));
 sg13g2_a21oi_1 _6171_ (.A1(_2252_),
    .A2(_2264_),
    .Y(_2266_),
    .B1(net974));
 sg13g2_a221oi_1 _6172_ (.B2(_2266_),
    .C1(_2257_),
    .B1(_2265_),
    .A1(net974),
    .Y(_2267_),
    .A2(_2264_));
 sg13g2_a21oi_1 _6173_ (.A1(net1180),
    .A2(net836),
    .Y(_2268_),
    .B1(_2267_));
 sg13g2_nor2_1 _6174_ (.A(net1023),
    .B(net2357),
    .Y(_0307_));
 sg13g2_nand3_1 _6175_ (.B(net1180),
    .C(net1181),
    .A(\led_controller.cpu.register_y[2] ),
    .Y(_2269_));
 sg13g2_a21o_1 _6176_ (.A2(net1181),
    .A1(net1180),
    .B1(\led_controller.cpu.register_y[2] ),
    .X(_2270_));
 sg13g2_nand2_1 _6177_ (.Y(_2271_),
    .A(_2269_),
    .B(_2270_));
 sg13g2_o21ai_1 _6178_ (.B1(_2251_),
    .Y(_2272_),
    .A1(_2253_),
    .A2(_2271_));
 sg13g2_a21oi_1 _6179_ (.A1(net870),
    .A2(_2253_),
    .Y(_2273_),
    .B1(_2272_));
 sg13g2_nor3_1 _6180_ (.A(\led_controller.cpu.register_y[2] ),
    .B(net1180),
    .C(net1181),
    .Y(_2274_));
 sg13g2_o21ai_1 _6181_ (.B1(\led_controller.cpu.register_y[2] ),
    .Y(_2275_),
    .A1(net1180),
    .A2(net1181));
 sg13g2_nor2b_1 _6182_ (.A(_2274_),
    .B_N(_2275_),
    .Y(_2276_));
 sg13g2_a21oi_1 _6183_ (.A1(net973),
    .A2(_2276_),
    .Y(_2277_),
    .B1(_2273_));
 sg13g2_o21ai_1 _6184_ (.B1(net1045),
    .Y(_2278_),
    .A1(_2257_),
    .A2(_2277_));
 sg13g2_a21oi_1 _6185_ (.A1(_0861_),
    .A2(net836),
    .Y(_0308_),
    .B1(_2278_));
 sg13g2_nor2_2 _6186_ (.A(_0860_),
    .B(_2269_),
    .Y(_2279_));
 sg13g2_xnor2_1 _6187_ (.Y(_2280_),
    .A(_0860_),
    .B(_2269_));
 sg13g2_and2_1 _6188_ (.A(_0860_),
    .B(_2274_),
    .X(_2281_));
 sg13g2_xnor2_1 _6189_ (.Y(_2282_),
    .A(_0860_),
    .B(_2274_));
 sg13g2_a21oi_1 _6190_ (.A1(net972),
    .A2(_2280_),
    .Y(_2283_),
    .B1(net973));
 sg13g2_o21ai_1 _6191_ (.B1(_2283_),
    .Y(_2284_),
    .A1(net868),
    .A2(net972));
 sg13g2_a21oi_1 _6192_ (.A1(net973),
    .A2(_2282_),
    .Y(_2285_),
    .B1(net836));
 sg13g2_a221oi_1 _6193_ (.B2(_2285_),
    .C1(net1023),
    .B1(_2284_),
    .A1(_0860_),
    .Y(_0309_),
    .A2(net836));
 sg13g2_nand2b_1 _6194_ (.Y(_2286_),
    .B(_2253_),
    .A_N(net845));
 sg13g2_xor2_1 _6195_ (.B(_2279_),
    .A(net1179),
    .X(_2287_));
 sg13g2_nor2_1 _6196_ (.A(_2253_),
    .B(_2287_),
    .Y(_2288_));
 sg13g2_nor2_1 _6197_ (.A(net973),
    .B(_2288_),
    .Y(_2289_));
 sg13g2_nand2b_1 _6198_ (.Y(_2290_),
    .B(_2281_),
    .A_N(net1179));
 sg13g2_xor2_1 _6199_ (.B(_2281_),
    .A(net1179),
    .X(_2291_));
 sg13g2_nor2_1 _6200_ (.A(net1179),
    .B(_2258_),
    .Y(_2292_));
 sg13g2_a221oi_1 _6201_ (.B2(net973),
    .C1(_2257_),
    .B1(_2291_),
    .A1(_2286_),
    .Y(_2293_),
    .A2(_2289_));
 sg13g2_nor3_1 _6202_ (.A(net1023),
    .B(_2292_),
    .C(_2293_),
    .Y(_0310_));
 sg13g2_nand3_1 _6203_ (.B(net1179),
    .C(_2279_),
    .A(net1177),
    .Y(_2294_));
 sg13g2_a21o_1 _6204_ (.A2(_2279_),
    .A1(net1179),
    .B1(net1177),
    .X(_2295_));
 sg13g2_and2_1 _6205_ (.A(_2294_),
    .B(_2295_),
    .X(_2296_));
 sg13g2_a21oi_1 _6206_ (.A1(net972),
    .A2(_2296_),
    .Y(_2297_),
    .B1(net973));
 sg13g2_o21ai_1 _6207_ (.B1(_2297_),
    .Y(_2298_),
    .A1(net844),
    .A2(net972));
 sg13g2_nor2_1 _6208_ (.A(net1177),
    .B(_2290_),
    .Y(_2299_));
 sg13g2_a21oi_1 _6209_ (.A1(net1177),
    .A2(_2290_),
    .Y(_2300_),
    .B1(_2251_));
 sg13g2_nand2b_1 _6210_ (.Y(_2301_),
    .B(_2300_),
    .A_N(_2299_));
 sg13g2_nor2_1 _6211_ (.A(net1177),
    .B(_2258_),
    .Y(_2302_));
 sg13g2_a21oi_1 _6212_ (.A1(_2298_),
    .A2(_2301_),
    .Y(_2303_),
    .B1(net836));
 sg13g2_nor3_1 _6213_ (.A(net1023),
    .B(_2302_),
    .C(_2303_),
    .Y(_0311_));
 sg13g2_nand4_1 _6214_ (.B(net1177),
    .C(net1179),
    .A(\led_controller.cpu.register_y[6] ),
    .Y(_2304_),
    .D(_2279_));
 sg13g2_xnor2_1 _6215_ (.Y(_2305_),
    .A(\led_controller.cpu.register_y[6] ),
    .B(_2294_));
 sg13g2_a21o_1 _6216_ (.A2(_2305_),
    .A1(net972),
    .B1(net974),
    .X(_2306_));
 sg13g2_a21oi_1 _6217_ (.A1(net843),
    .A2(_2253_),
    .Y(_2307_),
    .B1(_2306_));
 sg13g2_nor2b_1 _6218_ (.A(_2299_),
    .B_N(\led_controller.cpu.register_y[6] ),
    .Y(_2308_));
 sg13g2_nor3_1 _6219_ (.A(\led_controller.cpu.register_y[6] ),
    .B(net1177),
    .C(_2290_),
    .Y(_2309_));
 sg13g2_nor3_1 _6220_ (.A(_2251_),
    .B(_2308_),
    .C(_2309_),
    .Y(_2310_));
 sg13g2_o21ai_1 _6221_ (.B1(_2258_),
    .Y(_2311_),
    .A1(_2307_),
    .A2(_2310_));
 sg13g2_o21ai_1 _6222_ (.B1(_2311_),
    .Y(_2312_),
    .A1(net2335),
    .A2(_2258_));
 sg13g2_nor2_1 _6223_ (.A(net1023),
    .B(_2312_),
    .Y(_0312_));
 sg13g2_xnor2_1 _6224_ (.Y(_2313_),
    .A(\led_controller.cpu.register_y[7] ),
    .B(_2304_));
 sg13g2_nand2_1 _6225_ (.Y(_2314_),
    .A(net972),
    .B(_2313_));
 sg13g2_o21ai_1 _6226_ (.B1(_2314_),
    .Y(_2315_),
    .A1(net841),
    .A2(net972));
 sg13g2_nand2_1 _6227_ (.Y(_2316_),
    .A(_2251_),
    .B(_2315_));
 sg13g2_xnor2_1 _6228_ (.Y(_2317_),
    .A(_0859_),
    .B(_2309_));
 sg13g2_a21oi_1 _6229_ (.A1(net974),
    .A2(_2317_),
    .Y(_2318_),
    .B1(net836));
 sg13g2_a221oi_1 _6230_ (.B2(_2318_),
    .C1(net1023),
    .B1(_2316_),
    .A1(_0859_),
    .Y(_0313_),
    .A2(net836));
 sg13g2_a22oi_1 _6231_ (.Y(_2319_),
    .B1(_1858_),
    .B2(_1814_),
    .A2(_1852_),
    .A1(_1819_));
 sg13g2_nor2_2 _6232_ (.A(_1063_),
    .B(_2319_),
    .Y(_2320_));
 sg13g2_xnor2_1 _6233_ (.Y(_2321_),
    .A(_0859_),
    .B(net841));
 sg13g2_nand2_1 _6234_ (.Y(_2322_),
    .A(net1178),
    .B(net844));
 sg13g2_xnor2_1 _6235_ (.Y(_2323_),
    .A(net1178),
    .B(net844));
 sg13g2_nor2b_1 _6236_ (.A(\led_controller.cpu.register_y[4] ),
    .B_N(net845),
    .Y(_2324_));
 sg13g2_nor2b_1 _6237_ (.A(net845),
    .B_N(net1179),
    .Y(_2325_));
 sg13g2_nor3_1 _6238_ (.A(_2323_),
    .B(_2324_),
    .C(_2325_),
    .Y(_2326_));
 sg13g2_nand2b_1 _6239_ (.Y(_2327_),
    .B(\led_controller.cpu.register_y[2] ),
    .A_N(net870));
 sg13g2_nand2b_1 _6240_ (.Y(_2328_),
    .B(\led_controller.cpu.register_y[3] ),
    .A_N(net868));
 sg13g2_nand2_1 _6241_ (.Y(_2329_),
    .A(_2327_),
    .B(_2328_));
 sg13g2_nand2b_1 _6242_ (.Y(_2330_),
    .B(net843),
    .A_N(\led_controller.cpu.register_y[6] ));
 sg13g2_nand2_1 _6243_ (.Y(_2331_),
    .A(_0860_),
    .B(net868));
 sg13g2_nand2_1 _6244_ (.Y(_2332_),
    .A(_2328_),
    .B(_2331_));
 sg13g2_a21oi_1 _6245_ (.A1(_0861_),
    .A2(net870),
    .Y(_2333_),
    .B1(_2332_));
 sg13g2_nand4_1 _6246_ (.B(_2327_),
    .C(_2330_),
    .A(_2326_),
    .Y(_2334_),
    .D(_2333_));
 sg13g2_nand2_1 _6247_ (.Y(_2335_),
    .A(\led_controller.cpu.register_y[1] ),
    .B(_1887_));
 sg13g2_nand2b_1 _6248_ (.Y(_2336_),
    .B(_1849_),
    .A_N(\led_controller.cpu.register_y[0] ));
 sg13g2_o21ai_1 _6249_ (.B1(_2336_),
    .Y(_2337_),
    .A1(\led_controller.cpu.register_y[1] ),
    .A2(_1887_));
 sg13g2_a21oi_1 _6250_ (.A1(_2335_),
    .A2(_2337_),
    .Y(_2338_),
    .B1(_2334_));
 sg13g2_nand2_1 _6251_ (.Y(_2339_),
    .A(\led_controller.cpu.register_y[6] ),
    .B(_2055_));
 sg13g2_nand3_1 _6252_ (.B(_2329_),
    .C(_2331_),
    .A(_2326_),
    .Y(_2340_));
 sg13g2_o21ai_1 _6253_ (.B1(_2325_),
    .Y(_2341_),
    .A1(net1177),
    .A2(net844));
 sg13g2_nand4_1 _6254_ (.B(_2339_),
    .C(_2340_),
    .A(_2322_),
    .Y(_2342_),
    .D(_2341_));
 sg13g2_a21oi_1 _6255_ (.A1(_2330_),
    .A2(_2342_),
    .Y(_2343_),
    .B1(_2338_));
 sg13g2_nor2b_1 _6256_ (.A(_2343_),
    .B_N(_2321_),
    .Y(_2344_));
 sg13g2_a21oi_1 _6257_ (.A1(\led_controller.cpu.register_y[7] ),
    .A2(net841),
    .Y(_2345_),
    .B1(_2344_));
 sg13g2_nand2_1 _6258_ (.Y(_2346_),
    .A(\led_controller.cpu.register_y[0] ),
    .B(_1848_));
 sg13g2_nand3_1 _6259_ (.B(_2339_),
    .C(_2346_),
    .A(_2335_),
    .Y(_2347_));
 sg13g2_nor4_1 _6260_ (.A(_2334_),
    .B(_2337_),
    .C(_2345_),
    .D(_2347_),
    .Y(_2348_));
 sg13g2_nor2b_1 _6261_ (.A(_2348_),
    .B_N(_2320_),
    .Y(_2349_));
 sg13g2_xnor2_1 _6262_ (.Y(_2350_),
    .A(_2321_),
    .B(_2343_));
 sg13g2_nand2_1 _6263_ (.Y(_2351_),
    .A(_2320_),
    .B(_2350_));
 sg13g2_a22oi_1 _6264_ (.Y(_2352_),
    .B1(_1857_),
    .B2(_1815_),
    .A2(_1819_),
    .A1(_1814_));
 sg13g2_nor2_2 _6265_ (.A(_1063_),
    .B(_2352_),
    .Y(_2353_));
 sg13g2_or4_1 _6266_ (.A(_1849_),
    .B(net870),
    .C(net868),
    .D(_2286_),
    .X(_2354_));
 sg13g2_nand4_1 _6267_ (.B(_2055_),
    .C(net841),
    .A(net844),
    .Y(_2355_),
    .D(_2190_));
 sg13g2_o21ai_1 _6268_ (.B1(_2251_),
    .Y(_2356_),
    .A1(_2354_),
    .A2(_2355_));
 sg13g2_nor3_1 _6269_ (.A(\led_controller.cpu.register_y[3] ),
    .B(\led_controller.cpu.register_y[2] ),
    .C(net1180),
    .Y(_2357_));
 sg13g2_nand2_1 _6270_ (.Y(_2358_),
    .A(net1181),
    .B(_2357_));
 sg13g2_or4_1 _6271_ (.A(_2287_),
    .B(_2296_),
    .C(_2305_),
    .D(_2358_),
    .X(_2359_));
 sg13g2_o21ai_1 _6272_ (.B1(net973),
    .Y(_2360_),
    .A1(_2313_),
    .A2(_2359_));
 sg13g2_nand3_1 _6273_ (.B(_2356_),
    .C(_2360_),
    .A(net980),
    .Y(_2361_));
 sg13g2_nand2_1 _6274_ (.Y(_2362_),
    .A(_0864_),
    .B(net1185));
 sg13g2_nor4_1 _6275_ (.A(net1182),
    .B(net1183),
    .C(\led_controller.cpu.register_x[1] ),
    .D(_2362_),
    .Y(_2363_));
 sg13g2_nor2_1 _6276_ (.A(net979),
    .B(_2244_),
    .Y(_2364_));
 sg13g2_nand4_1 _6277_ (.B(_2234_),
    .C(_2363_),
    .A(_2225_),
    .Y(_2365_),
    .D(_2364_));
 sg13g2_a21oi_1 _6278_ (.A1(_2361_),
    .A2(_2365_),
    .Y(_2366_),
    .B1(_2353_));
 sg13g2_nor2_1 _6279_ (.A(_2320_),
    .B(_2366_),
    .Y(_2367_));
 sg13g2_nand2_1 _6280_ (.Y(_2368_),
    .A(\led_controller.cpu.register_x[7] ),
    .B(net841));
 sg13g2_nand2_1 _6281_ (.Y(_2369_),
    .A(_0862_),
    .B(net843));
 sg13g2_nand2_1 _6282_ (.Y(_2370_),
    .A(net1184),
    .B(_1887_));
 sg13g2_nand2b_1 _6283_ (.Y(_2371_),
    .B(_1849_),
    .A_N(net1185));
 sg13g2_o21ai_1 _6284_ (.B1(_2371_),
    .Y(_2372_),
    .A1(net1184),
    .A2(_1887_));
 sg13g2_nand2_1 _6285_ (.Y(_2373_),
    .A(\led_controller.cpu.register_x[5] ),
    .B(_2022_));
 sg13g2_or2_1 _6286_ (.X(_2374_),
    .B(_2022_),
    .A(\led_controller.cpu.register_x[5] ));
 sg13g2_nand2b_1 _6287_ (.Y(_2375_),
    .B(net1182),
    .A_N(net845));
 sg13g2_nand3_1 _6288_ (.B(_2374_),
    .C(_2375_),
    .A(_2373_),
    .Y(_2376_));
 sg13g2_a21oi_1 _6289_ (.A1(_0863_),
    .A2(_1989_),
    .Y(_2377_),
    .B1(_2376_));
 sg13g2_nand2b_1 _6290_ (.Y(_2378_),
    .B(\led_controller.cpu.register_x[3] ),
    .A_N(net869));
 sg13g2_nand2_1 _6291_ (.Y(_2379_),
    .A(_0864_),
    .B(net869));
 sg13g2_xnor2_1 _6292_ (.Y(_2380_),
    .A(\led_controller.cpu.register_x[2] ),
    .B(_1918_));
 sg13g2_nand4_1 _6293_ (.B(_2378_),
    .C(_2379_),
    .A(_2377_),
    .Y(_2381_),
    .D(_2380_));
 sg13g2_a21oi_1 _6294_ (.A1(_2370_),
    .A2(_2372_),
    .Y(_2382_),
    .B1(_2381_));
 sg13g2_o21ai_1 _6295_ (.B1(_2378_),
    .Y(_2383_),
    .A1(_0865_),
    .A2(_1918_));
 sg13g2_nand3_1 _6296_ (.B(_2379_),
    .C(_2383_),
    .A(_2377_),
    .Y(_2384_));
 sg13g2_nand2_1 _6297_ (.Y(_2385_),
    .A(\led_controller.cpu.register_x[6] ),
    .B(_2055_));
 sg13g2_nand3b_1 _6298_ (.B(_2374_),
    .C(\led_controller.cpu.register_x[4] ),
    .Y(_2386_),
    .A_N(_1989_));
 sg13g2_nand4_1 _6299_ (.B(_2384_),
    .C(_2385_),
    .A(_2373_),
    .Y(_2387_),
    .D(_2386_));
 sg13g2_o21ai_1 _6300_ (.B1(_2369_),
    .Y(_2388_),
    .A1(_2382_),
    .A2(_2387_));
 sg13g2_o21ai_1 _6301_ (.B1(_2353_),
    .Y(_2389_),
    .A1(\led_controller.cpu.register_x[7] ),
    .A2(net841));
 sg13g2_a21o_1 _6302_ (.A2(_2388_),
    .A1(_2368_),
    .B1(_2389_),
    .X(_2390_));
 sg13g2_or2_1 _6303_ (.X(_2391_),
    .B(_2388_),
    .A(_2368_));
 sg13g2_nand2_1 _6304_ (.Y(_2392_),
    .A(\led_controller.cpu.register_x[0] ),
    .B(_1848_));
 sg13g2_nand4_1 _6305_ (.B(_2370_),
    .C(_2385_),
    .A(_2369_),
    .Y(_2393_),
    .D(_2392_));
 sg13g2_nor3_1 _6306_ (.A(_2372_),
    .B(_2381_),
    .C(_2393_),
    .Y(_2394_));
 sg13g2_nand2_1 _6307_ (.Y(_2395_),
    .A(_2391_),
    .B(_2394_));
 sg13g2_o21ai_1 _6308_ (.B1(_2367_),
    .Y(_2396_),
    .A1(_2390_),
    .A2(_2395_));
 sg13g2_nor3_1 _6309_ (.A(_2184_),
    .B(_2320_),
    .C(_2353_),
    .Y(_2397_));
 sg13g2_o21ai_1 _6310_ (.B1(net836),
    .Y(_2398_),
    .A1(net874),
    .A2(_2397_));
 sg13g2_nand3b_1 _6311_ (.B(_2351_),
    .C(_2396_),
    .Y(_2399_),
    .A_N(_2349_));
 sg13g2_nand2_1 _6312_ (.Y(_2400_),
    .A(_2398_),
    .B(_2399_));
 sg13g2_o21ai_1 _6313_ (.B1(_2400_),
    .Y(_2401_),
    .A1(net2186),
    .A2(_2398_));
 sg13g2_nor2_1 _6314_ (.A(net1024),
    .B(_2401_),
    .Y(_0314_));
 sg13g2_nor2_1 _6315_ (.A(_2391_),
    .B(_2394_),
    .Y(_2402_));
 sg13g2_nand2b_1 _6316_ (.Y(_2403_),
    .B(_2313_),
    .A_N(_2359_));
 sg13g2_nand3_1 _6317_ (.B(_2317_),
    .C(_2403_),
    .A(net973),
    .Y(_2404_));
 sg13g2_o21ai_1 _6318_ (.B1(net977),
    .Y(_2405_),
    .A1(_0859_),
    .A2(_2253_));
 sg13g2_a21o_1 _6319_ (.A2(_2253_),
    .A1(_2089_),
    .B1(_2405_),
    .X(_2406_));
 sg13g2_o21ai_1 _6320_ (.B1(_2406_),
    .Y(_2407_),
    .A1(\led_controller.cpu.register_x[7] ),
    .A2(net977));
 sg13g2_o21ai_1 _6321_ (.B1(_2404_),
    .Y(_2408_),
    .A1(net974),
    .A2(_2407_));
 sg13g2_nand4_1 _6322_ (.B(_2234_),
    .C(_2244_),
    .A(_2225_),
    .Y(_2409_),
    .D(_2363_));
 sg13g2_a221oi_1 _6323_ (.B2(_2248_),
    .C1(_2353_),
    .B1(_2409_),
    .A1(net980),
    .Y(_2410_),
    .A2(_2408_));
 sg13g2_nor2_1 _6324_ (.A(_2320_),
    .B(_2410_),
    .Y(_2411_));
 sg13g2_o21ai_1 _6325_ (.B1(_2411_),
    .Y(_2412_),
    .A1(_2390_),
    .A2(_2402_));
 sg13g2_o21ai_1 _6326_ (.B1(_2349_),
    .Y(_2413_),
    .A1(_2345_),
    .A2(_2350_));
 sg13g2_nand3_1 _6327_ (.B(_2412_),
    .C(_2413_),
    .A(_2398_),
    .Y(_2414_));
 sg13g2_o21ai_1 _6328_ (.B1(_2414_),
    .Y(_2415_),
    .A1(net2196),
    .A2(_2398_));
 sg13g2_nor2_1 _6329_ (.A(net1024),
    .B(_2415_),
    .Y(_0315_));
 sg13g2_and2_1 _6330_ (.A(\led_controller.cpu.i_timer_100hz ),
    .B(_1093_),
    .X(_2416_));
 sg13g2_nor2b_1 _6331_ (.A(net2232),
    .B_N(_2416_),
    .Y(_2417_));
 sg13g2_nand3_1 _6332_ (.B(_1852_),
    .C(_1855_),
    .A(_1062_),
    .Y(_2418_));
 sg13g2_nor2_2 _6333_ (.A(net876),
    .B(_2418_),
    .Y(_2419_));
 sg13g2_nor2_2 _6334_ (.A(_2416_),
    .B(_2419_),
    .Y(_2420_));
 sg13g2_a21oi_1 _6335_ (.A1(net2232),
    .A2(_2420_),
    .Y(_2421_),
    .B1(_2417_));
 sg13g2_nand2_1 _6336_ (.Y(_2422_),
    .A(_1849_),
    .B(_2419_));
 sg13g2_a21oi_1 _6337_ (.A1(_2421_),
    .A2(_2422_),
    .Y(_0316_),
    .B1(net1032));
 sg13g2_xor2_1 _6338_ (.B(_2417_),
    .A(net2288),
    .X(_2423_));
 sg13g2_a21oi_1 _6339_ (.A1(_1886_),
    .A2(_2419_),
    .Y(_2424_),
    .B1(_2423_));
 sg13g2_nor2_1 _6340_ (.A(net1032),
    .B(_2424_),
    .Y(_0317_));
 sg13g2_o21ai_1 _6341_ (.B1(net2142),
    .Y(_2425_),
    .A1(\led_controller.cpu.stall_counter[1] ),
    .A2(\led_controller.cpu.stall_counter[0] ));
 sg13g2_nand2b_1 _6342_ (.Y(_2426_),
    .B(_2425_),
    .A_N(_1089_));
 sg13g2_nand3_1 _6343_ (.B(_1093_),
    .C(_2426_),
    .A(\led_controller.cpu.i_timer_100hz ),
    .Y(_2427_));
 sg13g2_a22oi_1 _6344_ (.Y(_2428_),
    .B1(_2420_),
    .B2(net2142),
    .A2(_2419_),
    .A1(_1918_));
 sg13g2_a21oi_1 _6345_ (.A1(_2427_),
    .A2(_2428_),
    .Y(_0318_),
    .B1(net1032));
 sg13g2_nand2_1 _6346_ (.Y(_2429_),
    .A(_1090_),
    .B(_2416_));
 sg13g2_nand2_1 _6347_ (.Y(_2430_),
    .A(net1626),
    .B(_2420_));
 sg13g2_xor2_1 _6348_ (.B(_1089_),
    .A(net1626),
    .X(_2431_));
 sg13g2_a22oi_1 _6349_ (.Y(_2432_),
    .B1(_2431_),
    .B2(_2416_),
    .A2(_2419_),
    .A1(net869));
 sg13g2_a21oi_1 _6350_ (.A1(_2430_),
    .A2(_2432_),
    .Y(_0319_),
    .B1(net1032));
 sg13g2_xnor2_1 _6351_ (.Y(_2433_),
    .A(net2313),
    .B(_2429_));
 sg13g2_a21oi_1 _6352_ (.A1(_1989_),
    .A2(_2419_),
    .Y(_2434_),
    .B1(_2433_));
 sg13g2_nor2_1 _6353_ (.A(net1032),
    .B(_2434_),
    .Y(_0320_));
 sg13g2_nor3_1 _6354_ (.A(net2342),
    .B(net2313),
    .C(_2429_),
    .Y(_2435_));
 sg13g2_o21ai_1 _6355_ (.B1(net2342),
    .Y(_2436_),
    .A1(net2313),
    .A2(_2429_));
 sg13g2_nand2b_1 _6356_ (.Y(_2437_),
    .B(_2436_),
    .A_N(_2435_));
 sg13g2_a21oi_1 _6357_ (.A1(_2023_),
    .A2(_2419_),
    .Y(_2438_),
    .B1(_2437_));
 sg13g2_nor2_1 _6358_ (.A(net1025),
    .B(_2438_),
    .Y(_0321_));
 sg13g2_xor2_1 _6359_ (.B(_2435_),
    .A(net2211),
    .X(_2439_));
 sg13g2_a21oi_1 _6360_ (.A1(_2054_),
    .A2(_2419_),
    .Y(_2440_),
    .B1(net2212));
 sg13g2_nor2_1 _6361_ (.A(net1032),
    .B(_2440_),
    .Y(_0322_));
 sg13g2_nand3_1 _6362_ (.B(\led_controller.cpu.i_timer_100hz ),
    .C(_1092_),
    .A(net1531),
    .Y(_2441_));
 sg13g2_o21ai_1 _6363_ (.B1(_2441_),
    .Y(_2442_),
    .A1(net842),
    .A2(_2416_));
 sg13g2_o21ai_1 _6364_ (.B1(net1047),
    .Y(_2443_),
    .A1(_2420_),
    .A2(_2442_));
 sg13g2_a21oi_1 _6365_ (.A1(_0857_),
    .A2(_2420_),
    .Y(_0323_),
    .B1(_2443_));
 sg13g2_nand2_1 _6366_ (.Y(_2444_),
    .A(_1050_),
    .B(_1841_));
 sg13g2_nor3_2 _6367_ (.A(_1064_),
    .B(net876),
    .C(_2444_),
    .Y(_2445_));
 sg13g2_nor2_1 _6368_ (.A(net1612),
    .B(_2445_),
    .Y(_2446_));
 sg13g2_and2_1 _6369_ (.A(net936),
    .B(_2445_),
    .X(_2447_));
 sg13g2_nor3_1 _6370_ (.A(net1035),
    .B(_2446_),
    .C(_2447_),
    .Y(_0324_));
 sg13g2_nor2_1 _6371_ (.A(net1591),
    .B(_2445_),
    .Y(_2448_));
 sg13g2_and2_1 _6372_ (.A(net932),
    .B(_2445_),
    .X(_2449_));
 sg13g2_nor3_1 _6373_ (.A(net1035),
    .B(_2448_),
    .C(_2449_),
    .Y(_0325_));
 sg13g2_nor2_1 _6374_ (.A(net1133),
    .B(\led_controller.cpu.bus_hi_valid ),
    .Y(_2450_));
 sg13g2_nand2b_2 _6375_ (.Y(_2451_),
    .B(\led_controller.cpu.i_bus_data_valid ),
    .A_N(\led_controller.cpu.bus_hi_valid ));
 sg13g2_nand2_2 _6376_ (.Y(_2452_),
    .A(net835),
    .B(_2451_));
 sg13g2_nand2_1 _6377_ (.Y(_2453_),
    .A(\led_controller.cpu.fetch_pc[0] ),
    .B(net948));
 sg13g2_a22oi_1 _6378_ (.Y(_2454_),
    .B1(net848),
    .B2(net2369),
    .A2(net948),
    .A1(net1971));
 sg13g2_o21ai_1 _6379_ (.B1(_2454_),
    .Y(_2455_),
    .A1(net2375),
    .A2(_1236_));
 sg13g2_xor2_1 _6380_ (.B(_2455_),
    .A(net828),
    .X(_2456_));
 sg13g2_nor2_1 _6381_ (.A(net1039),
    .B(_2456_),
    .Y(_0326_));
 sg13g2_xor2_1 _6382_ (.B(\led_controller.cpu.o_bus_addr[0] ),
    .A(\led_controller.cpu.o_bus_addr[1] ),
    .X(_2457_));
 sg13g2_o21ai_1 _6383_ (.B1(_1230_),
    .Y(_2458_),
    .A1(net948),
    .A2(_2457_));
 sg13g2_nand3_1 _6384_ (.B(net828),
    .C(_2458_),
    .A(_1228_),
    .Y(_2459_));
 sg13g2_o21ai_1 _6385_ (.B1(_2459_),
    .Y(_2460_),
    .A1(net2287),
    .A2(net828));
 sg13g2_nor2_1 _6386_ (.A(net1039),
    .B(_2460_),
    .Y(_0327_));
 sg13g2_and3_2 _6387_ (.X(_2461_),
    .A(\led_controller.cpu.o_bus_addr[2] ),
    .B(\led_controller.cpu.o_bus_addr[1] ),
    .C(\led_controller.cpu.o_bus_addr[0] ));
 sg13g2_a21oi_1 _6388_ (.A1(\led_controller.cpu.o_bus_addr[1] ),
    .A2(\led_controller.cpu.o_bus_addr[0] ),
    .Y(_2462_),
    .B1(net1728));
 sg13g2_o21ai_1 _6389_ (.B1(net1019),
    .Y(_2463_),
    .A1(_2461_),
    .A2(_2462_));
 sg13g2_a21oi_1 _6390_ (.A1(net830),
    .A2(_2463_),
    .Y(_2464_),
    .B1(_1234_));
 sg13g2_nor2_1 _6391_ (.A(net1728),
    .B(net828),
    .Y(_2465_));
 sg13g2_nor2_1 _6392_ (.A(_2464_),
    .B(_2465_),
    .Y(_0328_));
 sg13g2_nor2_1 _6393_ (.A(net2101),
    .B(_2452_),
    .Y(_2466_));
 sg13g2_xnor2_1 _6394_ (.Y(_2467_),
    .A(net2101),
    .B(_2461_));
 sg13g2_nand2_1 _6395_ (.Y(_2468_),
    .A(net1019),
    .B(_2467_));
 sg13g2_a21oi_1 _6396_ (.A1(net830),
    .A2(_2468_),
    .Y(_2469_),
    .B1(_1242_));
 sg13g2_nor2_1 _6397_ (.A(net2102),
    .B(_2469_),
    .Y(_0329_));
 sg13g2_nor2_1 _6398_ (.A(net1856),
    .B(net828),
    .Y(_2470_));
 sg13g2_and3_1 _6399_ (.X(_2471_),
    .A(\led_controller.cpu.o_bus_addr[4] ),
    .B(\led_controller.cpu.o_bus_addr[3] ),
    .C(_2461_));
 sg13g2_a21oi_1 _6400_ (.A1(\led_controller.cpu.o_bus_addr[3] ),
    .A2(_2461_),
    .Y(_2472_),
    .B1(net1856));
 sg13g2_o21ai_1 _6401_ (.B1(net1017),
    .Y(_2473_),
    .A1(_2471_),
    .A2(_2472_));
 sg13g2_a21oi_1 _6402_ (.A1(net830),
    .A2(_2473_),
    .Y(_2474_),
    .B1(_1246_));
 sg13g2_nor2_1 _6403_ (.A(_2470_),
    .B(_2474_),
    .Y(_0330_));
 sg13g2_nor2_1 _6404_ (.A(net1816),
    .B(_2452_),
    .Y(_2475_));
 sg13g2_and2_1 _6405_ (.A(net1816),
    .B(_2471_),
    .X(_2476_));
 sg13g2_nor2_1 _6406_ (.A(net1816),
    .B(_2471_),
    .Y(_2477_));
 sg13g2_o21ai_1 _6407_ (.B1(net1017),
    .Y(_2478_),
    .A1(_2476_),
    .A2(_2477_));
 sg13g2_a21oi_1 _6408_ (.A1(net829),
    .A2(_2478_),
    .Y(_2479_),
    .B1(_1249_));
 sg13g2_nor2_1 _6409_ (.A(net1817),
    .B(_2479_),
    .Y(_0331_));
 sg13g2_and2_1 _6410_ (.A(\led_controller.cpu.o_bus_addr[6] ),
    .B(_2476_),
    .X(_2480_));
 sg13g2_nand2_1 _6411_ (.Y(_2481_),
    .A(net1019),
    .B(_2480_));
 sg13g2_o21ai_1 _6412_ (.B1(_2481_),
    .Y(_2482_),
    .A1(net2220),
    .A2(_2476_));
 sg13g2_o21ai_1 _6413_ (.B1(_1253_),
    .Y(_2483_),
    .A1(_1236_),
    .A2(_2482_));
 sg13g2_o21ai_1 _6414_ (.B1(_2483_),
    .Y(_2484_),
    .A1(net2220),
    .A2(_2452_));
 sg13g2_nor2_1 _6415_ (.A(net1038),
    .B(net2221),
    .Y(_0332_));
 sg13g2_and2_1 _6416_ (.A(net2388),
    .B(_2480_),
    .X(_2485_));
 sg13g2_nand2_1 _6417_ (.Y(_2486_),
    .A(net1019),
    .B(_2485_));
 sg13g2_o21ai_1 _6418_ (.B1(_2486_),
    .Y(_2487_),
    .A1(net2157),
    .A2(_2480_));
 sg13g2_o21ai_1 _6419_ (.B1(_1257_),
    .Y(_2488_),
    .A1(_1236_),
    .A2(_2487_));
 sg13g2_o21ai_1 _6420_ (.B1(_2488_),
    .Y(_2489_),
    .A1(net2157),
    .A2(net827));
 sg13g2_nor2_1 _6421_ (.A(net1038),
    .B(net2158),
    .Y(_0333_));
 sg13g2_and2_1 _6422_ (.A(net2146),
    .B(_2485_),
    .X(_2490_));
 sg13g2_nand2_1 _6423_ (.Y(_2491_),
    .A(net1017),
    .B(_2490_));
 sg13g2_o21ai_1 _6424_ (.B1(_2491_),
    .Y(_2492_),
    .A1(net2146),
    .A2(_2485_));
 sg13g2_o21ai_1 _6425_ (.B1(_1262_),
    .Y(_2493_),
    .A1(_1236_),
    .A2(_2492_));
 sg13g2_o21ai_1 _6426_ (.B1(_2493_),
    .Y(_2494_),
    .A1(net2146),
    .A2(net827));
 sg13g2_nor2_1 _6427_ (.A(net1038),
    .B(_2494_),
    .Y(_0334_));
 sg13g2_and2_1 _6428_ (.A(\led_controller.cpu.o_bus_addr[9] ),
    .B(_2490_),
    .X(_2495_));
 sg13g2_nand2_1 _6429_ (.Y(_2496_),
    .A(net1017),
    .B(_2495_));
 sg13g2_o21ai_1 _6430_ (.B1(_2496_),
    .Y(_2497_),
    .A1(net2193),
    .A2(_2490_));
 sg13g2_o21ai_1 _6431_ (.B1(_1267_),
    .Y(_2498_),
    .A1(_1236_),
    .A2(_2497_));
 sg13g2_o21ai_1 _6432_ (.B1(_2498_),
    .Y(_2499_),
    .A1(net2193),
    .A2(net828));
 sg13g2_nor2_1 _6433_ (.A(net1038),
    .B(net2194),
    .Y(_0335_));
 sg13g2_o21ai_1 _6434_ (.B1(net828),
    .Y(_2500_),
    .A1(_1271_),
    .A2(_2495_));
 sg13g2_and2_1 _6435_ (.A(net1602),
    .B(_2495_),
    .X(_2501_));
 sg13g2_nand2_1 _6436_ (.Y(_2502_),
    .A(net1017),
    .B(_2501_));
 sg13g2_a22oi_1 _6437_ (.Y(_2503_),
    .B1(_2502_),
    .B2(net829),
    .A2(_1271_),
    .A1(net1052));
 sg13g2_a21oi_1 _6438_ (.A1(_0812_),
    .A2(_2500_),
    .Y(_0336_),
    .B1(_2503_));
 sg13g2_o21ai_1 _6439_ (.B1(net834),
    .Y(_2504_),
    .A1(net2190),
    .A2(_2501_));
 sg13g2_and2_1 _6440_ (.A(net2190),
    .B(_2501_),
    .X(_2505_));
 sg13g2_a21o_1 _6441_ (.A2(_2505_),
    .A1(net1017),
    .B1(_2504_),
    .X(_2506_));
 sg13g2_o21ai_1 _6442_ (.B1(net1052),
    .Y(_2507_),
    .A1(net2190),
    .A2(net827));
 sg13g2_a21oi_1 _6443_ (.A1(_1277_),
    .A2(_2506_),
    .Y(_0337_),
    .B1(_2507_));
 sg13g2_nand2_1 _6444_ (.Y(_2508_),
    .A(net2236),
    .B(_2505_));
 sg13g2_o21ai_1 _6445_ (.B1(net834),
    .Y(_2509_),
    .A1(\led_controller.cpu.o_bus_addr[12] ),
    .A2(_2505_));
 sg13g2_nand2b_1 _6446_ (.Y(_2510_),
    .B(_2508_),
    .A_N(_2509_));
 sg13g2_nand4_1 _6447_ (.B(_1282_),
    .C(net827),
    .A(_1278_),
    .Y(_2511_),
    .D(_2510_));
 sg13g2_o21ai_1 _6448_ (.B1(_2511_),
    .Y(_2512_),
    .A1(net2236),
    .A2(net827));
 sg13g2_nor2_1 _6449_ (.A(net1037),
    .B(net2237),
    .Y(_0338_));
 sg13g2_nand2_1 _6450_ (.Y(_2513_),
    .A(_1285_),
    .B(_2508_));
 sg13g2_a21oi_1 _6451_ (.A1(net827),
    .A2(_2513_),
    .Y(_2514_),
    .B1(net1537));
 sg13g2_and3_2 _6452_ (.X(_2515_),
    .A(net1537),
    .B(\led_controller.cpu.o_bus_addr[12] ),
    .C(_2505_));
 sg13g2_nand2_1 _6453_ (.Y(_2516_),
    .A(net1017),
    .B(_2515_));
 sg13g2_a21oi_1 _6454_ (.A1(net829),
    .A2(_2516_),
    .Y(_2517_),
    .B1(_1286_));
 sg13g2_nor2_1 _6455_ (.A(net1538),
    .B(_2517_),
    .Y(_0339_));
 sg13g2_nand2_1 _6456_ (.Y(_2518_),
    .A(\led_controller.cpu.o_bus_addr[14] ),
    .B(_2515_));
 sg13g2_nand3_1 _6457_ (.B(net1017),
    .C(_2515_),
    .A(net2218),
    .Y(_2519_));
 sg13g2_and2_1 _6458_ (.A(net834),
    .B(_2519_),
    .X(_2520_));
 sg13g2_o21ai_1 _6459_ (.B1(_2520_),
    .Y(_2521_),
    .A1(net2218),
    .A2(_2515_));
 sg13g2_o21ai_1 _6460_ (.B1(net1050),
    .Y(_2522_),
    .A1(net2218),
    .A2(net827));
 sg13g2_a21oi_1 _6461_ (.A1(_1290_),
    .A2(_2521_),
    .Y(_0340_),
    .B1(_2522_));
 sg13g2_nor3_1 _6462_ (.A(net1621),
    .B(_1236_),
    .C(_2518_),
    .Y(_2523_));
 sg13g2_o21ai_1 _6463_ (.B1(net827),
    .Y(_2524_),
    .A1(_1294_),
    .A2(_2523_));
 sg13g2_nand2_1 _6464_ (.Y(_2525_),
    .A(net1621),
    .B(_2520_));
 sg13g2_a21oi_1 _6465_ (.A1(_2524_),
    .A2(net1622),
    .Y(_0341_),
    .B1(net1039));
 sg13g2_and2_1 _6466_ (.A(\led_controller.cpu.i_bus_data_valid ),
    .B(net1617),
    .X(_2526_));
 sg13g2_o21ai_1 _6467_ (.B1(net830),
    .Y(_0342_),
    .A1(_0856_),
    .A2(net1094));
 sg13g2_nand2_1 _6468_ (.Y(_2527_),
    .A(net1573),
    .B(net1095));
 sg13g2_nand2_1 _6469_ (.Y(_2528_),
    .A(\led_controller.cpu.i_bus_data[0] ),
    .B(net1018));
 sg13g2_a21oi_1 _6470_ (.A1(_2527_),
    .A2(_2528_),
    .Y(_0343_),
    .B1(net1029));
 sg13g2_nand2_1 _6471_ (.Y(_2529_),
    .A(net1453),
    .B(net1095));
 sg13g2_nand2_1 _6472_ (.Y(_2530_),
    .A(\led_controller.cpu.i_bus_data[1] ),
    .B(net1018));
 sg13g2_a21oi_1 _6473_ (.A1(_2529_),
    .A2(_2530_),
    .Y(_0344_),
    .B1(net1028));
 sg13g2_nand2_1 _6474_ (.Y(_2531_),
    .A(net1459),
    .B(net1095));
 sg13g2_nand2_1 _6475_ (.Y(_2532_),
    .A(\led_controller.cpu.i_bus_data[2] ),
    .B(net1018));
 sg13g2_a21oi_1 _6476_ (.A1(_2531_),
    .A2(_2532_),
    .Y(_0345_),
    .B1(net1028));
 sg13g2_nand2_1 _6477_ (.Y(_2533_),
    .A(net1440),
    .B(net1095));
 sg13g2_nand2_1 _6478_ (.Y(_2534_),
    .A(\led_controller.cpu.i_bus_data[3] ),
    .B(net1018));
 sg13g2_a21oi_1 _6479_ (.A1(_2533_),
    .A2(_2534_),
    .Y(_0346_),
    .B1(net1028));
 sg13g2_nand2_1 _6480_ (.Y(_2535_),
    .A(net1541),
    .B(net1095));
 sg13g2_nand2_1 _6481_ (.Y(_2536_),
    .A(\led_controller.cpu.i_bus_data[4] ),
    .B(net1018));
 sg13g2_a21oi_1 _6482_ (.A1(_2535_),
    .A2(_2536_),
    .Y(_0347_),
    .B1(net1029));
 sg13g2_nand2_1 _6483_ (.Y(_2537_),
    .A(net1373),
    .B(net1095));
 sg13g2_nand2_1 _6484_ (.Y(_2538_),
    .A(\led_controller.cpu.i_bus_data[5] ),
    .B(net1018));
 sg13g2_a21oi_1 _6485_ (.A1(_2537_),
    .A2(_2538_),
    .Y(_0348_),
    .B1(net1028));
 sg13g2_nand2_1 _6486_ (.Y(_2539_),
    .A(net1416),
    .B(net1095));
 sg13g2_nand2_1 _6487_ (.Y(_2540_),
    .A(\led_controller.cpu.i_bus_data[6] ),
    .B(net1018));
 sg13g2_a21oi_1 _6488_ (.A1(_2539_),
    .A2(_2540_),
    .Y(_0349_),
    .B1(net1028));
 sg13g2_nand2_1 _6489_ (.Y(_2541_),
    .A(net1418),
    .B(net1095));
 sg13g2_nand2_1 _6490_ (.Y(_2542_),
    .A(\led_controller.cpu.i_bus_data[7] ),
    .B(net1018));
 sg13g2_a21oi_1 _6491_ (.A1(_2541_),
    .A2(_2542_),
    .Y(_0350_),
    .B1(net1028));
 sg13g2_o21ai_1 _6492_ (.B1(net1059),
    .Y(_2543_),
    .A1(\led_controller.cpu.fetch_instruction[4] ),
    .A2(net945));
 sg13g2_a21oi_1 _6493_ (.A1(_0851_),
    .A2(net946),
    .Y(_0355_),
    .B1(_2543_));
 sg13g2_o21ai_1 _6494_ (.B1(net1059),
    .Y(_2544_),
    .A1(\led_controller.cpu.fetch_instruction[5] ),
    .A2(net945));
 sg13g2_a21oi_1 _6495_ (.A1(_0850_),
    .A2(net945),
    .Y(_0356_),
    .B1(_2544_));
 sg13g2_o21ai_1 _6496_ (.B1(net1047),
    .Y(_2545_),
    .A1(\led_controller.cpu.fetch_instruction[6] ),
    .A2(net944));
 sg13g2_a21oi_1 _6497_ (.A1(_0849_),
    .A2(net944),
    .Y(_0357_),
    .B1(_2545_));
 sg13g2_o21ai_1 _6498_ (.B1(net1049),
    .Y(_2546_),
    .A1(\led_controller.cpu.fetch_instruction[7] ),
    .A2(net944));
 sg13g2_a21oi_1 _6499_ (.A1(_0848_),
    .A2(net944),
    .Y(_0358_),
    .B1(_2546_));
 sg13g2_o21ai_1 _6500_ (.B1(net1046),
    .Y(_2547_),
    .A1(net1573),
    .A2(net937));
 sg13g2_a21oi_1 _6501_ (.A1(_0847_),
    .A2(net937),
    .Y(_0359_),
    .B1(_2547_));
 sg13g2_o21ai_1 _6502_ (.B1(net1046),
    .Y(_2548_),
    .A1(net1453),
    .A2(net944));
 sg13g2_a21oi_1 _6503_ (.A1(_0846_),
    .A2(net937),
    .Y(_0360_),
    .B1(_2548_));
 sg13g2_o21ai_1 _6504_ (.B1(net1046),
    .Y(_2549_),
    .A1(net1459),
    .A2(net937));
 sg13g2_a21oi_1 _6505_ (.A1(_0845_),
    .A2(net937),
    .Y(_0361_),
    .B1(_2549_));
 sg13g2_o21ai_1 _6506_ (.B1(net1046),
    .Y(_2550_),
    .A1(net1440),
    .A2(net937));
 sg13g2_a21oi_1 _6507_ (.A1(_0844_),
    .A2(net937),
    .Y(_0362_),
    .B1(_2550_));
 sg13g2_o21ai_1 _6508_ (.B1(net1046),
    .Y(_2551_),
    .A1(net1541),
    .A2(net938));
 sg13g2_a21oi_1 _6509_ (.A1(_0843_),
    .A2(net937),
    .Y(_0363_),
    .B1(_2551_));
 sg13g2_o21ai_1 _6510_ (.B1(net1046),
    .Y(_2552_),
    .A1(\led_controller.cpu.fetch_instruction[13] ),
    .A2(net944));
 sg13g2_a21oi_1 _6511_ (.A1(_0842_),
    .A2(net944),
    .Y(_0364_),
    .B1(_2552_));
 sg13g2_o21ai_1 _6512_ (.B1(net1047),
    .Y(_2553_),
    .A1(\led_controller.cpu.fetch_instruction[14] ),
    .A2(net947));
 sg13g2_a21oi_1 _6513_ (.A1(_0841_),
    .A2(net944),
    .Y(_0365_),
    .B1(_2553_));
 sg13g2_o21ai_1 _6514_ (.B1(net1048),
    .Y(_2554_),
    .A1(\led_controller.cpu.fetch_instruction[15] ),
    .A2(net938));
 sg13g2_a21oi_1 _6515_ (.A1(_0840_),
    .A2(net938),
    .Y(_0366_),
    .B1(_2554_));
 sg13g2_nand2_1 _6516_ (.Y(_2555_),
    .A(net1551),
    .B(net942));
 sg13g2_a21oi_1 _6517_ (.A1(_2453_),
    .A2(_2555_),
    .Y(_0367_),
    .B1(net1029));
 sg13g2_nand2_1 _6518_ (.Y(_2556_),
    .A(net1651),
    .B(net943));
 sg13g2_a21oi_1 _6519_ (.A1(_1229_),
    .A2(_2556_),
    .Y(_0368_),
    .B1(net1039));
 sg13g2_o21ai_1 _6520_ (.B1(net1048),
    .Y(_2557_),
    .A1(\led_controller.cpu.fetch_pc[2] ),
    .A2(net942));
 sg13g2_a21oi_1 _6521_ (.A1(_0839_),
    .A2(net942),
    .Y(_0369_),
    .B1(_2557_));
 sg13g2_o21ai_1 _6522_ (.B1(net1044),
    .Y(_2558_),
    .A1(\led_controller.cpu.fetch_pc[3] ),
    .A2(net942));
 sg13g2_a21oi_1 _6523_ (.A1(_0838_),
    .A2(net942),
    .Y(_0370_),
    .B1(_2558_));
 sg13g2_o21ai_1 _6524_ (.B1(net1044),
    .Y(_2559_),
    .A1(\led_controller.cpu.fetch_pc[4] ),
    .A2(net942));
 sg13g2_a21oi_1 _6525_ (.A1(_0836_),
    .A2(net942),
    .Y(_0371_),
    .B1(_2559_));
 sg13g2_o21ai_1 _6526_ (.B1(net1044),
    .Y(_2560_),
    .A1(\led_controller.cpu.fetch_pc[5] ),
    .A2(net940));
 sg13g2_a21oi_1 _6527_ (.A1(_0835_),
    .A2(net940),
    .Y(_0372_),
    .B1(_2560_));
 sg13g2_o21ai_1 _6528_ (.B1(net1044),
    .Y(_2561_),
    .A1(\led_controller.cpu.fetch_pc[6] ),
    .A2(net940));
 sg13g2_a21oi_1 _6529_ (.A1(_0834_),
    .A2(net942),
    .Y(_0373_),
    .B1(_2561_));
 sg13g2_o21ai_1 _6530_ (.B1(net1044),
    .Y(_2562_),
    .A1(net1977),
    .A2(net948));
 sg13g2_a21oi_1 _6531_ (.A1(_0833_),
    .A2(net948),
    .Y(_0374_),
    .B1(_2562_));
 sg13g2_o21ai_1 _6532_ (.B1(net1043),
    .Y(_2563_),
    .A1(\led_controller.cpu.fetch_pc[8] ),
    .A2(net940));
 sg13g2_a21oi_1 _6533_ (.A1(_0832_),
    .A2(net941),
    .Y(_0375_),
    .B1(_2563_));
 sg13g2_o21ai_1 _6534_ (.B1(net1043),
    .Y(_2564_),
    .A1(\led_controller.cpu.fetch_pc[9] ),
    .A2(net941));
 sg13g2_a21oi_1 _6535_ (.A1(_0831_),
    .A2(net941),
    .Y(_0376_),
    .B1(_2564_));
 sg13g2_o21ai_1 _6536_ (.B1(net1043),
    .Y(_2565_),
    .A1(\led_controller.cpu.fetch_pc[10] ),
    .A2(net940));
 sg13g2_a21oi_1 _6537_ (.A1(_0830_),
    .A2(net943),
    .Y(_0377_),
    .B1(_2565_));
 sg13g2_o21ai_1 _6538_ (.B1(net1043),
    .Y(_2566_),
    .A1(\led_controller.cpu.fetch_pc[11] ),
    .A2(net939));
 sg13g2_a21oi_1 _6539_ (.A1(_0829_),
    .A2(net941),
    .Y(_0378_),
    .B1(_2566_));
 sg13g2_o21ai_1 _6540_ (.B1(net1043),
    .Y(_2567_),
    .A1(\led_controller.cpu.fetch_pc[12] ),
    .A2(net939));
 sg13g2_a21oi_1 _6541_ (.A1(_0828_),
    .A2(net941),
    .Y(_0379_),
    .B1(_2567_));
 sg13g2_o21ai_1 _6542_ (.B1(net1043),
    .Y(_2568_),
    .A1(\led_controller.cpu.fetch_pc[13] ),
    .A2(net940));
 sg13g2_a21oi_1 _6543_ (.A1(_0827_),
    .A2(net939),
    .Y(_0380_),
    .B1(_2568_));
 sg13g2_o21ai_1 _6544_ (.B1(net1043),
    .Y(_2569_),
    .A1(\led_controller.cpu.fetch_pc[14] ),
    .A2(net939));
 sg13g2_a21oi_1 _6545_ (.A1(_0826_),
    .A2(net939),
    .Y(_0381_),
    .B1(_2569_));
 sg13g2_o21ai_1 _6546_ (.B1(net1043),
    .Y(_2570_),
    .A1(\led_controller.cpu.fetch_pc[15] ),
    .A2(net941));
 sg13g2_a21oi_1 _6547_ (.A1(_0825_),
    .A2(net941),
    .Y(_0382_),
    .B1(_2570_));
 sg13g2_a21oi_1 _6548_ (.A1(_0824_),
    .A2(net945),
    .Y(_0383_),
    .B1(net1034));
 sg13g2_nor2_1 _6549_ (.A(\led_controller.cpu.i_bus_data_valid ),
    .B(net1617),
    .Y(_2571_));
 sg13g2_nor3_1 _6550_ (.A(net1029),
    .B(net1093),
    .C(net1618),
    .Y(_0384_));
 sg13g2_o21ai_1 _6551_ (.B1(net830),
    .Y(_2572_),
    .A1(net1836),
    .A2(net1094));
 sg13g2_inv_1 _6552_ (.Y(_0385_),
    .A(net1837));
 sg13g2_nor2_1 _6553_ (.A(net1971),
    .B(_1226_),
    .Y(_2573_));
 sg13g2_nor2b_1 _6554_ (.A(\led_controller.cpu.pc[0] ),
    .B_N(_1226_),
    .Y(_2574_));
 sg13g2_nor3_1 _6555_ (.A(net1029),
    .B(net1972),
    .C(_2574_),
    .Y(_0386_));
 sg13g2_nor4_1 _6556_ (.A(net1032),
    .B(_1064_),
    .C(_1095_),
    .D(_2444_),
    .Y(_0387_));
 sg13g2_nor4_1 _6557_ (.A(net1718),
    .B(\led_controller.flash.cs_delay_counter[4] ),
    .C(net1566),
    .D(net1605),
    .Y(_2575_));
 sg13g2_nor4_1 _6558_ (.A(_0886_),
    .B(net764),
    .C(\led_controller.flash.cs_delay_counter[3] ),
    .D(net1555),
    .Y(_2576_));
 sg13g2_nand4_1 _6559_ (.B(_0997_),
    .C(_2575_),
    .A(net1575),
    .Y(_2577_),
    .D(_2576_));
 sg13g2_nand2_1 _6560_ (.Y(_2578_),
    .A(net1942),
    .B(net854));
 sg13g2_nand3_1 _6561_ (.B(_2577_),
    .C(_2578_),
    .A(net1058),
    .Y(_0388_));
 sg13g2_o21ai_1 _6562_ (.B1(net1053),
    .Y(_2579_),
    .A1(\led_controller.cpu.o_bus_addr[0] ),
    .A2(net854));
 sg13g2_a21oi_1 _6563_ (.A1(_0822_),
    .A2(net853),
    .Y(_0389_),
    .B1(_2579_));
 sg13g2_o21ai_1 _6564_ (.B1(net1053),
    .Y(_2580_),
    .A1(\led_controller.cpu.o_bus_addr[1] ),
    .A2(net854));
 sg13g2_a21oi_1 _6565_ (.A1(_0821_),
    .A2(net853),
    .Y(_0390_),
    .B1(_2580_));
 sg13g2_o21ai_1 _6566_ (.B1(net1053),
    .Y(_2581_),
    .A1(\led_controller.cpu.o_bus_addr[2] ),
    .A2(net854));
 sg13g2_a21oi_1 _6567_ (.A1(_0820_),
    .A2(net853),
    .Y(_0391_),
    .B1(_2581_));
 sg13g2_o21ai_1 _6568_ (.B1(net1053),
    .Y(_2582_),
    .A1(\led_controller.cpu.o_bus_addr[3] ),
    .A2(net853));
 sg13g2_a21oi_1 _6569_ (.A1(_0819_),
    .A2(net853),
    .Y(_0392_),
    .B1(_2582_));
 sg13g2_o21ai_1 _6570_ (.B1(net1053),
    .Y(_2583_),
    .A1(\led_controller.cpu.o_bus_addr[4] ),
    .A2(net853));
 sg13g2_a21oi_1 _6571_ (.A1(_0818_),
    .A2(net852),
    .Y(_0393_),
    .B1(_2583_));
 sg13g2_o21ai_1 _6572_ (.B1(net1051),
    .Y(_2584_),
    .A1(\led_controller.cpu.o_bus_addr[5] ),
    .A2(net852));
 sg13g2_a21oi_1 _6573_ (.A1(_0817_),
    .A2(net852),
    .Y(_0394_),
    .B1(_2584_));
 sg13g2_o21ai_1 _6574_ (.B1(net1051),
    .Y(_2585_),
    .A1(\led_controller.cpu.o_bus_addr[6] ),
    .A2(net852));
 sg13g2_a21oi_1 _6575_ (.A1(_0816_),
    .A2(net855),
    .Y(_0395_),
    .B1(_2585_));
 sg13g2_o21ai_1 _6576_ (.B1(net1050),
    .Y(_2586_),
    .A1(\led_controller.cpu.o_bus_addr[7] ),
    .A2(net851));
 sg13g2_a21oi_1 _6577_ (.A1(_0815_),
    .A2(net851),
    .Y(_0396_),
    .B1(_2586_));
 sg13g2_o21ai_1 _6578_ (.B1(net1050),
    .Y(_2587_),
    .A1(\led_controller.cpu.o_bus_addr[8] ),
    .A2(net853));
 sg13g2_a21oi_1 _6579_ (.A1(_0814_),
    .A2(net853),
    .Y(_0397_),
    .B1(_2587_));
 sg13g2_o21ai_1 _6580_ (.B1(net1051),
    .Y(_2588_),
    .A1(\led_controller.cpu.o_bus_addr[9] ),
    .A2(net852));
 sg13g2_a21oi_1 _6581_ (.A1(_0813_),
    .A2(net852),
    .Y(_0398_),
    .B1(_2588_));
 sg13g2_o21ai_1 _6582_ (.B1(net1051),
    .Y(_2589_),
    .A1(\led_controller.cpu.o_bus_addr[10] ),
    .A2(net852));
 sg13g2_a21oi_1 _6583_ (.A1(_0811_),
    .A2(net852),
    .Y(_0399_),
    .B1(_2589_));
 sg13g2_o21ai_1 _6584_ (.B1(net1050),
    .Y(_2590_),
    .A1(\led_controller.cpu.o_bus_addr[11] ),
    .A2(net851));
 sg13g2_a21oi_1 _6585_ (.A1(_0810_),
    .A2(net850),
    .Y(_0400_),
    .B1(_2590_));
 sg13g2_o21ai_1 _6586_ (.B1(net1050),
    .Y(_2591_),
    .A1(\led_controller.cpu.o_bus_addr[12] ),
    .A2(net850));
 sg13g2_a21oi_1 _6587_ (.A1(_0809_),
    .A2(net850),
    .Y(_0401_),
    .B1(_2591_));
 sg13g2_o21ai_1 _6588_ (.B1(net1050),
    .Y(_2592_),
    .A1(\led_controller.cpu.o_bus_addr[13] ),
    .A2(net850));
 sg13g2_a21oi_1 _6589_ (.A1(_0808_),
    .A2(net850),
    .Y(_0402_),
    .B1(_2592_));
 sg13g2_o21ai_1 _6590_ (.B1(net1050),
    .Y(_2593_),
    .A1(\led_controller.cpu.o_bus_addr[14] ),
    .A2(net850));
 sg13g2_a21oi_1 _6591_ (.A1(_0807_),
    .A2(net850),
    .Y(_0403_),
    .B1(_2593_));
 sg13g2_o21ai_1 _6592_ (.B1(net1050),
    .Y(_2594_),
    .A1(\led_controller.cpu.o_bus_addr[15] ),
    .A2(net850));
 sg13g2_a21oi_1 _6593_ (.A1(_0806_),
    .A2(net851),
    .Y(_0404_),
    .B1(_2594_));
 sg13g2_a21oi_1 _6594_ (.A1(_0889_),
    .A2(_0991_),
    .Y(_2595_),
    .B1(_0990_));
 sg13g2_a221oi_1 _6595_ (.B2(net1343),
    .C1(_0991_),
    .B1(net2087),
    .A1(net1437),
    .Y(_2596_),
    .A2(net1193));
 sg13g2_o21ai_1 _6596_ (.B1(net1056),
    .Y(_2597_),
    .A1(net1522),
    .A2(net833));
 sg13g2_a21oi_1 _6597_ (.A1(net833),
    .A2(_2596_),
    .Y(_0405_),
    .B1(_2597_));
 sg13g2_a221oi_1 _6598_ (.B2(net1384),
    .C1(_0991_),
    .B1(net2087),
    .A1(net1400),
    .Y(_2598_),
    .A2(net1193));
 sg13g2_o21ai_1 _6599_ (.B1(net1054),
    .Y(_2599_),
    .A1(net2243),
    .A2(net833));
 sg13g2_a21oi_1 _6600_ (.A1(net833),
    .A2(_2598_),
    .Y(_0406_),
    .B1(_2599_));
 sg13g2_a22oi_1 _6601_ (.Y(_2600_),
    .B1(net2087),
    .B2(net1378),
    .A2(net1936),
    .A1(net1474));
 sg13g2_o21ai_1 _6602_ (.B1(net1054),
    .Y(_2601_),
    .A1(net1610),
    .A2(net833));
 sg13g2_a21oi_1 _6603_ (.A1(_2595_),
    .A2(_2600_),
    .Y(_0407_),
    .B1(_2601_));
 sg13g2_a22oi_1 _6604_ (.Y(_2602_),
    .B1(net1192),
    .B2(net1325),
    .A2(net1193),
    .A1(net1492));
 sg13g2_o21ai_1 _6605_ (.B1(net1054),
    .Y(_2603_),
    .A1(net2100),
    .A2(net833));
 sg13g2_a21oi_1 _6606_ (.A1(net833),
    .A2(_2602_),
    .Y(_0408_),
    .B1(_2603_));
 sg13g2_a22oi_1 _6607_ (.Y(_2604_),
    .B1(net1192),
    .B2(net1329),
    .A2(net1193),
    .A1(net1430));
 sg13g2_o21ai_1 _6608_ (.B1(net1054),
    .Y(_2605_),
    .A1(net2154),
    .A2(net832));
 sg13g2_a21oi_1 _6609_ (.A1(net832),
    .A2(_2604_),
    .Y(_0409_),
    .B1(_2605_));
 sg13g2_a22oi_1 _6610_ (.Y(_2606_),
    .B1(net1192),
    .B2(net1356),
    .A2(net1193),
    .A1(net1382));
 sg13g2_o21ai_1 _6611_ (.B1(net1054),
    .Y(_2607_),
    .A1(net1584),
    .A2(net832));
 sg13g2_a21oi_1 _6612_ (.A1(net832),
    .A2(_2606_),
    .Y(_0410_),
    .B1(_2607_));
 sg13g2_a22oi_1 _6613_ (.Y(_2608_),
    .B1(net1192),
    .B2(net1321),
    .A2(net1193),
    .A1(net1398));
 sg13g2_o21ai_1 _6614_ (.B1(net1054),
    .Y(_2609_),
    .A1(net2136),
    .A2(net832));
 sg13g2_a21oi_1 _6615_ (.A1(net832),
    .A2(_2608_),
    .Y(_0411_),
    .B1(_2609_));
 sg13g2_a22oi_1 _6616_ (.Y(_2610_),
    .B1(net1192),
    .B2(net1389),
    .A2(net1193),
    .A1(net1370));
 sg13g2_o21ai_1 _6617_ (.B1(net1054),
    .Y(_2611_),
    .A1(net2089),
    .A2(net832));
 sg13g2_a21oi_1 _6618_ (.A1(net832),
    .A2(_2610_),
    .Y(_0412_),
    .B1(_2611_));
 sg13g2_and2_1 _6619_ (.A(net1353),
    .B(_0908_),
    .X(_0413_));
 sg13g2_and2_1 _6620_ (.A(net1803),
    .B(_1775_),
    .X(_2612_));
 sg13g2_o21ai_1 _6621_ (.B1(net1055),
    .Y(_2613_),
    .A1(net1176),
    .A2(_1010_));
 sg13g2_nor2_1 _6622_ (.A(net1803),
    .B(_1775_),
    .Y(_2614_));
 sg13g2_nor3_1 _6623_ (.A(_2612_),
    .B(net970),
    .C(net1804),
    .Y(_0414_));
 sg13g2_xnor2_1 _6624_ (.Y(_2615_),
    .A(net2079),
    .B(_2612_));
 sg13g2_nor2_1 _6625_ (.A(net970),
    .B(net2080),
    .Y(_0415_));
 sg13g2_a21oi_1 _6626_ (.A1(\led_controller.flash.master.bit_counter[2] ),
    .A2(_2612_),
    .Y(_2616_),
    .B1(net1683));
 sg13g2_and3_1 _6627_ (.X(_2617_),
    .A(net1683),
    .B(\led_controller.flash.master.bit_counter[2] ),
    .C(_2612_));
 sg13g2_nor2_1 _6628_ (.A(net1333),
    .B(_1783_),
    .Y(_2618_));
 sg13g2_nor4_1 _6629_ (.A(net970),
    .B(net1684),
    .C(_2617_),
    .D(_2618_),
    .Y(_0416_));
 sg13g2_and2_1 _6630_ (.A(net1176),
    .B(net1563),
    .X(_2619_));
 sg13g2_nor2_1 _6631_ (.A(net1176),
    .B(net1563),
    .Y(_2620_));
 sg13g2_nor4_1 _6632_ (.A(_1772_),
    .B(net970),
    .C(_2619_),
    .D(net1564),
    .Y(_0417_));
 sg13g2_xnor2_1 _6633_ (.Y(_2621_),
    .A(net1899),
    .B(_2619_));
 sg13g2_nor2_1 _6634_ (.A(net971),
    .B(_2621_),
    .Y(_0418_));
 sg13g2_a21oi_1 _6635_ (.A1(\led_controller.flash.master.sck_counter[1] ),
    .A2(_2619_),
    .Y(_2622_),
    .B1(net1525));
 sg13g2_and3_1 _6636_ (.X(_2623_),
    .A(net1525),
    .B(\led_controller.flash.master.sck_counter[1] ),
    .C(_2619_));
 sg13g2_nor3_1 _6637_ (.A(net971),
    .B(net1526),
    .C(_2623_),
    .Y(_0419_));
 sg13g2_nor2_1 _6638_ (.A(net1823),
    .B(_2623_),
    .Y(_2624_));
 sg13g2_and2_1 _6639_ (.A(net1823),
    .B(_2623_),
    .X(_2625_));
 sg13g2_nor3_1 _6640_ (.A(net971),
    .B(net1824),
    .C(_2625_),
    .Y(_0420_));
 sg13g2_a21oi_1 _6641_ (.A1(net2167),
    .A2(_2625_),
    .Y(_2626_),
    .B1(net970));
 sg13g2_o21ai_1 _6642_ (.B1(_2626_),
    .Y(_2627_),
    .A1(net2167),
    .A2(_2625_));
 sg13g2_inv_1 _6643_ (.Y(_0421_),
    .A(_2627_));
 sg13g2_a21oi_1 _6644_ (.A1(\led_controller.flash.master.sck_counter[4] ),
    .A2(_2625_),
    .Y(_2628_),
    .B1(net1519));
 sg13g2_and3_1 _6645_ (.X(_2629_),
    .A(net1519),
    .B(net2387),
    .C(_2625_));
 sg13g2_nor3_1 _6646_ (.A(net970),
    .B(net1520),
    .C(_2629_),
    .Y(_0422_));
 sg13g2_nor2_1 _6647_ (.A(net1926),
    .B(_2629_),
    .Y(_2630_));
 sg13g2_and2_1 _6648_ (.A(net1926),
    .B(_2629_),
    .X(_2631_));
 sg13g2_nor3_1 _6649_ (.A(net970),
    .B(net1927),
    .C(_2631_),
    .Y(_0423_));
 sg13g2_a21oi_1 _6650_ (.A1(net2161),
    .A2(_2631_),
    .Y(_2632_),
    .B1(net970));
 sg13g2_o21ai_1 _6651_ (.B1(_2632_),
    .Y(_2633_),
    .A1(net2161),
    .A2(_2631_));
 sg13g2_inv_1 _6652_ (.Y(_0424_),
    .A(_2633_));
 sg13g2_a221oi_1 _6653_ (.B2(_1006_),
    .C1(net1040),
    .B1(_0991_),
    .A1(_0804_),
    .Y(_0425_),
    .A2(net1608));
 sg13g2_o21ai_1 _6654_ (.B1(_1009_),
    .Y(_2634_),
    .A1(_0804_),
    .A2(_1010_));
 sg13g2_and3_1 _6655_ (.X(_2635_),
    .A(net1176),
    .B(net1055),
    .C(_2634_));
 sg13g2_or2_1 _6656_ (.X(_0426_),
    .B(_2635_),
    .A(_1778_));
 sg13g2_o21ai_1 _6657_ (.B1(net1058),
    .Y(_2636_),
    .A1(net5),
    .A2(_1774_));
 sg13g2_a21oi_1 _6658_ (.A1(_0803_),
    .A2(_1774_),
    .Y(_0427_),
    .B1(_2636_));
 sg13g2_o21ai_1 _6659_ (.B1(net1048),
    .Y(_2637_),
    .A1(\led_controller.cpu.i_bus_data[0] ),
    .A2(net966));
 sg13g2_a21oi_1 _6660_ (.A1(_0802_),
    .A2(net966),
    .Y(_0428_),
    .B1(_2637_));
 sg13g2_o21ai_1 _6661_ (.B1(net1048),
    .Y(_2638_),
    .A1(net1769),
    .A2(net968));
 sg13g2_a21oi_1 _6662_ (.A1(_0802_),
    .A2(net968),
    .Y(_0429_),
    .B1(_2638_));
 sg13g2_o21ai_1 _6663_ (.B1(net1049),
    .Y(_2639_),
    .A1(\led_controller.cpu.i_bus_data[2] ),
    .A2(net966));
 sg13g2_a21oi_1 _6664_ (.A1(_0801_),
    .A2(net966),
    .Y(_0430_),
    .B1(_2639_));
 sg13g2_o21ai_1 _6665_ (.B1(net1048),
    .Y(_2640_),
    .A1(net1628),
    .A2(net966));
 sg13g2_a21oi_1 _6666_ (.A1(_0800_),
    .A2(net966),
    .Y(_0431_),
    .B1(_2640_));
 sg13g2_o21ai_1 _6667_ (.B1(net1048),
    .Y(_2641_),
    .A1(net1806),
    .A2(net968));
 sg13g2_a21oi_1 _6668_ (.A1(_0800_),
    .A2(net968),
    .Y(_0432_),
    .B1(_2641_));
 sg13g2_o21ai_1 _6669_ (.B1(net1048),
    .Y(_2642_),
    .A1(\led_controller.cpu.i_bus_data[5] ),
    .A2(net966));
 sg13g2_a21oi_1 _6670_ (.A1(_0799_),
    .A2(net966),
    .Y(_0433_),
    .B1(_2642_));
 sg13g2_o21ai_1 _6671_ (.B1(net1048),
    .Y(_2643_),
    .A1(net1766),
    .A2(net968));
 sg13g2_a21oi_1 _6672_ (.A1(_0799_),
    .A2(net968),
    .Y(_0434_),
    .B1(_2643_));
 sg13g2_xnor2_1 _6673_ (.Y(_2644_),
    .A(_0798_),
    .B(_1009_));
 sg13g2_and2_1 _6674_ (.A(_2635_),
    .B(_2644_),
    .X(_0435_));
 sg13g2_o21ai_1 _6675_ (.B1(net1056),
    .Y(_2645_),
    .A1(net1566),
    .A2(_0987_));
 sg13g2_nor2_1 _6676_ (.A(net764),
    .B(_2645_),
    .Y(_0436_));
 sg13g2_nand2_1 _6677_ (.Y(_2646_),
    .A(net2343),
    .B(net764));
 sg13g2_a21o_1 _6678_ (.A2(_2646_),
    .A1(_0982_),
    .B1(_2645_),
    .X(_2647_));
 sg13g2_o21ai_1 _6679_ (.B1(_2647_),
    .Y(_0437_),
    .A1(net1041),
    .A2(net854));
 sg13g2_nand2_1 _6680_ (.Y(_2648_),
    .A(net1555),
    .B(_0982_));
 sg13g2_a221oi_1 _6681_ (.B2(_0983_),
    .C1(net1041),
    .B1(net1556),
    .A1(\led_controller.cpu.o_bus_addr_valid ),
    .Y(_0438_),
    .A2(_0988_));
 sg13g2_xor2_1 _6682_ (.B(_0983_),
    .A(net2117),
    .X(_2649_));
 sg13g2_nor2_1 _6683_ (.A(_2645_),
    .B(_2649_),
    .Y(_0439_));
 sg13g2_xnor2_1 _6684_ (.Y(_2650_),
    .A(net1956),
    .B(_0984_));
 sg13g2_nor2_1 _6685_ (.A(_2645_),
    .B(net1957),
    .Y(_0440_));
 sg13g2_nand2b_1 _6686_ (.Y(_2651_),
    .B(net1718),
    .A_N(_0985_));
 sg13g2_a21oi_1 _6687_ (.A1(_0986_),
    .A2(net1719),
    .Y(_0441_),
    .B1(_2645_));
 sg13g2_nand2_1 _6688_ (.Y(_2652_),
    .A(net1605),
    .B(_0986_));
 sg13g2_a21oi_1 _6689_ (.A1(_0987_),
    .A2(net1606),
    .Y(_0442_),
    .B1(_2645_));
 sg13g2_and3_1 _6690_ (.X(_0443_),
    .A(net1566),
    .B(net1057),
    .C(_0987_));
 sg13g2_nor3_1 _6691_ (.A(\led_controller.flash.master.bit_counter[3] ),
    .B(\led_controller.flash.master.bit_counter[2] ),
    .C(\led_controller.flash.master.bit_counter[1] ),
    .Y(_2653_));
 sg13g2_a21oi_1 _6692_ (.A1(\led_controller.flash.master.bit_counter[0] ),
    .A2(_2653_),
    .Y(_2654_),
    .B1(_1776_));
 sg13g2_mux2_1 _6693_ (.A0(\led_controller.flash.master.i_tx_data[7] ),
    .A1(\led_controller.flash.master.tx_data[7] ),
    .S(_2654_),
    .X(_2655_));
 sg13g2_o21ai_1 _6694_ (.B1(net1055),
    .Y(_2656_),
    .A1(_1781_),
    .A2(_2655_));
 sg13g2_a21oi_1 _6695_ (.A1(_0797_),
    .A2(_1781_),
    .Y(_0444_),
    .B1(_2656_));
 sg13g2_a22oi_1 _6696_ (.Y(_2657_),
    .B1(_2618_),
    .B2(net1522),
    .A2(_1784_),
    .A1(net1688));
 sg13g2_nor2_1 _6697_ (.A(net971),
    .B(net1689),
    .Y(_0445_));
 sg13g2_nand2b_2 _6698_ (.Y(_2658_),
    .B(_1124_),
    .A_N(_1101_));
 sg13g2_and2_1 _6699_ (.A(net1060),
    .B(net821),
    .X(_2659_));
 sg13g2_nand2_1 _6700_ (.Y(_2660_),
    .A(net1319),
    .B(_2659_));
 sg13g2_o21ai_1 _6701_ (.B1(_2660_),
    .Y(_0446_),
    .A1(net934),
    .A2(net821));
 sg13g2_nand2_1 _6702_ (.Y(_2661_),
    .A(net1295),
    .B(_2659_));
 sg13g2_o21ai_1 _6703_ (.B1(_2661_),
    .Y(_0447_),
    .A1(net933),
    .A2(_2658_));
 sg13g2_nand2_1 _6704_ (.Y(_2662_),
    .A(net1253),
    .B(_2659_));
 sg13g2_o21ai_1 _6705_ (.B1(_2662_),
    .Y(_0448_),
    .A1(net929),
    .A2(net821));
 sg13g2_nand2_1 _6706_ (.Y(_2663_),
    .A(net814),
    .B(_2659_));
 sg13g2_o21ai_1 _6707_ (.B1(_2663_),
    .Y(_0449_),
    .A1(net927),
    .A2(net821));
 sg13g2_nand2_1 _6708_ (.Y(_2664_),
    .A(net1246),
    .B(_2659_));
 sg13g2_o21ai_1 _6709_ (.B1(_2664_),
    .Y(_0450_),
    .A1(net925),
    .A2(net821));
 sg13g2_nand2_1 _6710_ (.Y(_2665_),
    .A(net1272),
    .B(_2659_));
 sg13g2_o21ai_1 _6711_ (.B1(_2665_),
    .Y(_0451_),
    .A1(net922),
    .A2(net821));
 sg13g2_nand2_1 _6712_ (.Y(_2666_),
    .A(net1318),
    .B(_2659_));
 sg13g2_o21ai_1 _6713_ (.B1(_2666_),
    .Y(_0452_),
    .A1(net919),
    .A2(net821));
 sg13g2_nand2_1 _6714_ (.Y(_2667_),
    .A(net1283),
    .B(_2659_));
 sg13g2_o21ai_1 _6715_ (.B1(_2667_),
    .Y(_0453_),
    .A1(net917),
    .A2(net821));
 sg13g2_nor3_2 _6716_ (.A(net2059),
    .B(net2118),
    .C(net2137),
    .Y(_2668_));
 sg13g2_nand2b_1 _6717_ (.Y(_2669_),
    .B(_0910_),
    .A_N(net2137));
 sg13g2_a21oi_1 _6718_ (.A1(_0890_),
    .A2(_2668_),
    .Y(_2670_),
    .B1(net1599));
 sg13g2_nor3_1 _6719_ (.A(\led_controller.led_effect_chase.finished ),
    .B(net1098),
    .C(_2669_),
    .Y(_2671_));
 sg13g2_o21ai_1 _6720_ (.B1(net1157),
    .Y(_2672_),
    .A1(_0890_),
    .A2(_2668_));
 sg13g2_nor3_1 _6721_ (.A(net1600),
    .B(_2671_),
    .C(_2672_),
    .Y(_0454_));
 sg13g2_nand2_1 _6722_ (.Y(_2673_),
    .A(net2379),
    .B(_1382_));
 sg13g2_nand3_1 _6723_ (.B(_0917_),
    .C(_2668_),
    .A(\led_controller.effect_chase_led_strb ),
    .Y(_2674_));
 sg13g2_nand2_1 _6724_ (.Y(_2675_),
    .A(_0890_),
    .B(_2674_));
 sg13g2_and2_1 _6725_ (.A(_2673_),
    .B(_2675_),
    .X(_2676_));
 sg13g2_xnor2_1 _6726_ (.Y(_2677_),
    .A(\led_controller.cpu.i_num_colors[1] ),
    .B(\led_controller.cpu.i_num_colors[0] ));
 sg13g2_xnor2_1 _6727_ (.Y(_2678_),
    .A(net2290),
    .B(_2677_));
 sg13g2_xor2_1 _6728_ (.B(\led_controller.effect_chase_led_color[0] ),
    .A(\led_controller.cpu.i_num_colors[0] ),
    .X(_2679_));
 sg13g2_a21oi_1 _6729_ (.A1(_2678_),
    .A2(_2679_),
    .Y(_2680_),
    .B1(\led_controller.led_effect_chase.finished ));
 sg13g2_nand3_1 _6730_ (.B(\led_controller.led_effect_chase.finished ),
    .C(_2668_),
    .A(net2162),
    .Y(_2681_));
 sg13g2_nor2_1 _6731_ (.A(net2290),
    .B(\led_controller.effect_chase_led_color[0] ),
    .Y(_2682_));
 sg13g2_a21oi_1 _6732_ (.A1(\led_controller.cpu.i_num_colors[0] ),
    .A2(_2682_),
    .Y(_2683_),
    .B1(_2681_));
 sg13g2_o21ai_1 _6733_ (.B1(_2676_),
    .Y(_2684_),
    .A1(_2680_),
    .A2(_2683_));
 sg13g2_mux2_1 _6734_ (.A0(_2684_),
    .A1(_2676_),
    .S(net2293),
    .X(_2685_));
 sg13g2_nor2_1 _6735_ (.A(net1120),
    .B(net2294),
    .Y(_0455_));
 sg13g2_and2_1 _6736_ (.A(net2290),
    .B(\led_controller.effect_chase_led_color[0] ),
    .X(_2686_));
 sg13g2_nor2_1 _6737_ (.A(_2682_),
    .B(_2686_),
    .Y(_2687_));
 sg13g2_a21oi_1 _6738_ (.A1(_2677_),
    .A2(_2682_),
    .Y(_2688_),
    .B1(_2686_));
 sg13g2_o21ai_1 _6739_ (.B1(_2676_),
    .Y(_2689_),
    .A1(_2681_),
    .A2(_2688_));
 sg13g2_a21oi_1 _6740_ (.A1(_2680_),
    .A2(_2687_),
    .Y(_2690_),
    .B1(_2689_));
 sg13g2_o21ai_1 _6741_ (.B1(net1157),
    .Y(_2691_),
    .A1(net2290),
    .A2(_2676_));
 sg13g2_nor2_1 _6742_ (.A(_2690_),
    .B(_2691_),
    .Y(_0456_));
 sg13g2_nor3_1 _6743_ (.A(net1333),
    .B(net1041),
    .C(_1783_),
    .Y(_0457_));
 sg13g2_or2_1 _6744_ (.X(_2692_),
    .B(\led_controller.cpu.i_num_leds[0] ),
    .A(\led_controller.cpu.i_num_leds[1] ));
 sg13g2_nor2_1 _6745_ (.A(\led_controller.cpu.i_num_leds[2] ),
    .B(_2692_),
    .Y(_2693_));
 sg13g2_nor3_1 _6746_ (.A(\led_controller.cpu.i_num_leds[3] ),
    .B(\led_controller.cpu.i_num_leds[2] ),
    .C(_2692_),
    .Y(_2694_));
 sg13g2_nor2b_1 _6747_ (.A(\led_controller.cpu.i_num_leds[4] ),
    .B_N(_2694_),
    .Y(_2695_));
 sg13g2_nor2b_1 _6748_ (.A(\led_controller.cpu.i_num_leds[5] ),
    .B_N(_2695_),
    .Y(_2696_));
 sg13g2_nor2b_1 _6749_ (.A(\led_controller.cpu.i_num_leds[6] ),
    .B_N(_2696_),
    .Y(_2697_));
 sg13g2_nand2b_2 _6750_ (.Y(_2698_),
    .B(\led_controller.cpu.i_num_leds[7] ),
    .A_N(_2697_));
 sg13g2_xnor2_1 _6751_ (.Y(_2699_),
    .A(\led_controller.cpu.i_num_leds[6] ),
    .B(_2696_));
 sg13g2_xor2_1 _6752_ (.B(_2695_),
    .A(\led_controller.cpu.i_num_leds[5] ),
    .X(_2700_));
 sg13g2_inv_1 _6753_ (.Y(_2701_),
    .A(_2700_));
 sg13g2_xor2_1 _6754_ (.B(_2700_),
    .A(\led_controller.led_effect_chase.current_led[5] ),
    .X(_2702_));
 sg13g2_xnor2_1 _6755_ (.Y(_2703_),
    .A(\led_controller.cpu.i_num_leds[4] ),
    .B(_2694_));
 sg13g2_nor2_1 _6756_ (.A(\led_controller.led_effect_chase.current_led[4] ),
    .B(_2703_),
    .Y(_2704_));
 sg13g2_xor2_1 _6757_ (.B(_2692_),
    .A(\led_controller.cpu.i_num_leds[2] ),
    .X(_2705_));
 sg13g2_nor2b_1 _6758_ (.A(\led_controller.cpu.i_num_leds[7] ),
    .B_N(_2697_),
    .Y(_2706_));
 sg13g2_xnor2_1 _6759_ (.Y(_2707_),
    .A(\led_controller.cpu.i_num_leds[3] ),
    .B(_2693_));
 sg13g2_xor2_1 _6760_ (.B(\led_controller.cpu.i_num_leds[0] ),
    .A(\led_controller.cpu.i_num_leds[1] ),
    .X(_2708_));
 sg13g2_xor2_1 _6761_ (.B(\led_controller.led_effect_chase.current_led[0] ),
    .A(\led_controller.cpu.i_num_leds[0] ),
    .X(_2709_));
 sg13g2_nor2_1 _6762_ (.A(net1653),
    .B(_2698_),
    .Y(_2710_));
 sg13g2_xnor2_1 _6763_ (.Y(_2711_),
    .A(net2330),
    .B(_2708_));
 sg13g2_a21oi_1 _6764_ (.A1(net2107),
    .A2(_2703_),
    .Y(_2712_),
    .B1(_2711_));
 sg13g2_xnor2_1 _6765_ (.Y(_2713_),
    .A(net2050),
    .B(_2707_));
 sg13g2_nor3_1 _6766_ (.A(_2702_),
    .B(_2706_),
    .C(_2713_),
    .Y(_2714_));
 sg13g2_xnor2_1 _6767_ (.Y(_2715_),
    .A(net1543),
    .B(_2699_));
 sg13g2_a21oi_1 _6768_ (.A1(net1653),
    .A2(_2698_),
    .Y(_2716_),
    .B1(_2715_));
 sg13g2_xnor2_1 _6769_ (.Y(_2717_),
    .A(\led_controller.led_effect_chase.current_led[2] ),
    .B(_2705_));
 sg13g2_nand3_1 _6770_ (.B(_2671_),
    .C(_2709_),
    .A(net1599),
    .Y(_2718_));
 sg13g2_nor4_1 _6771_ (.A(_2704_),
    .B(_2710_),
    .C(_2717_),
    .D(_2718_),
    .Y(_2719_));
 sg13g2_nand4_1 _6772_ (.B(_2714_),
    .C(_2716_),
    .A(_2712_),
    .Y(_2720_),
    .D(_2719_));
 sg13g2_o21ai_1 _6773_ (.B1(_2720_),
    .Y(_2721_),
    .A1(_2669_),
    .A2(_2673_));
 sg13g2_nand2b_2 _6774_ (.Y(_2722_),
    .B(_2675_),
    .A_N(_2721_));
 sg13g2_inv_1 _6775_ (.Y(_2723_),
    .A(_2722_));
 sg13g2_nor2_2 _6776_ (.A(\led_controller.led_effect_chase.finished ),
    .B(_2722_),
    .Y(_2724_));
 sg13g2_nand2_1 _6777_ (.Y(_2725_),
    .A(net2240),
    .B(_2723_));
 sg13g2_o21ai_1 _6778_ (.B1(_2725_),
    .Y(_2726_),
    .A1(net2240),
    .A2(_2724_));
 sg13g2_nor2_1 _6779_ (.A(net1120),
    .B(net2241),
    .Y(_0458_));
 sg13g2_nand2b_1 _6780_ (.Y(_2727_),
    .B(_2725_),
    .A_N(net2330));
 sg13g2_and2_1 _6781_ (.A(net2330),
    .B(net2240),
    .X(_2728_));
 sg13g2_o21ai_1 _6782_ (.B1(_2723_),
    .Y(_2729_),
    .A1(\led_controller.led_effect_chase.finished ),
    .A2(_2728_));
 sg13g2_and3_1 _6783_ (.X(_0459_),
    .A(net1157),
    .B(_2727_),
    .C(_2729_));
 sg13g2_nor2b_1 _6784_ (.A(net2130),
    .B_N(_2728_),
    .Y(_2730_));
 sg13g2_a22oi_1 _6785_ (.Y(_2731_),
    .B1(_2730_),
    .B2(_2724_),
    .A2(_2729_),
    .A1(net2130));
 sg13g2_nor2_1 _6786_ (.A(net1120),
    .B(net2131),
    .Y(_0460_));
 sg13g2_nand3_1 _6787_ (.B(\led_controller.led_effect_chase.current_led[2] ),
    .C(_2728_),
    .A(net2050),
    .Y(_2732_));
 sg13g2_a21o_1 _6788_ (.A2(_2728_),
    .A1(\led_controller.led_effect_chase.current_led[2] ),
    .B1(net2050),
    .X(_2733_));
 sg13g2_and2_1 _6789_ (.A(_2732_),
    .B(_2733_),
    .X(_2734_));
 sg13g2_a22oi_1 _6790_ (.Y(_2735_),
    .B1(_2724_),
    .B2(_2734_),
    .A2(_2722_),
    .A1(net2050));
 sg13g2_nor2_1 _6791_ (.A(net1120),
    .B(net2051),
    .Y(_0461_));
 sg13g2_nor2_1 _6792_ (.A(_0796_),
    .B(_2732_),
    .Y(_2736_));
 sg13g2_xnor2_1 _6793_ (.Y(_2737_),
    .A(net2107),
    .B(_2732_));
 sg13g2_a22oi_1 _6794_ (.Y(_2738_),
    .B1(_2724_),
    .B2(_2737_),
    .A2(_2722_),
    .A1(net2107));
 sg13g2_nor2_1 _6795_ (.A(net1121),
    .B(net2108),
    .Y(_0462_));
 sg13g2_and2_1 _6796_ (.A(net2114),
    .B(_2736_),
    .X(_2739_));
 sg13g2_inv_1 _6797_ (.Y(_2740_),
    .A(_2739_));
 sg13g2_a22oi_1 _6798_ (.Y(_2741_),
    .B1(_2724_),
    .B2(_2740_),
    .A2(_2722_),
    .A1(net2114));
 sg13g2_o21ai_1 _6799_ (.B1(net1157),
    .Y(_2742_),
    .A1(net2114),
    .A2(_2736_));
 sg13g2_nor2_1 _6800_ (.A(net2115),
    .B(_2742_),
    .Y(_0463_));
 sg13g2_a21oi_1 _6801_ (.A1(net1543),
    .A2(_2739_),
    .Y(_2743_),
    .B1(\led_controller.led_effect_chase.finished ));
 sg13g2_o21ai_1 _6802_ (.B1(net1157),
    .Y(_2744_),
    .A1(_2722_),
    .A2(_2743_));
 sg13g2_a21oi_1 _6803_ (.A1(_2724_),
    .A2(_2739_),
    .Y(_2745_),
    .B1(net1543));
 sg13g2_nor2_1 _6804_ (.A(_2744_),
    .B(net1544),
    .Y(_0464_));
 sg13g2_nor2_1 _6805_ (.A(net1653),
    .B(net1121),
    .Y(_2746_));
 sg13g2_nand4_1 _6806_ (.B(_2724_),
    .C(_2739_),
    .A(net1543),
    .Y(_2747_),
    .D(_2746_));
 sg13g2_o21ai_1 _6807_ (.B1(_2747_),
    .Y(_0465_),
    .A1(_0795_),
    .A2(_2744_));
 sg13g2_or2_1 _6808_ (.X(_2748_),
    .B(_1137_),
    .A(_1101_));
 sg13g2_and2_1 _6809_ (.A(net1060),
    .B(_2748_),
    .X(_2749_));
 sg13g2_nand2_1 _6810_ (.Y(_2750_),
    .A(net790),
    .B(_2749_));
 sg13g2_o21ai_1 _6811_ (.B1(_2750_),
    .Y(_0466_),
    .A1(net934),
    .A2(_2748_));
 sg13g2_nand2_1 _6812_ (.Y(_2751_),
    .A(net1247),
    .B(_2749_));
 sg13g2_o21ai_1 _6813_ (.B1(_2751_),
    .Y(_0467_),
    .A1(net933),
    .A2(_2748_));
 sg13g2_nand2_1 _6814_ (.Y(_2752_),
    .A(net1323),
    .B(_2749_));
 sg13g2_o21ai_1 _6815_ (.B1(_2752_),
    .Y(_0468_),
    .A1(_1113_),
    .A2(_2748_));
 sg13g2_nor3_1 _6816_ (.A(_1097_),
    .B(net927),
    .C(_1137_),
    .Y(_2753_));
 sg13g2_a21o_1 _6817_ (.A2(_2749_),
    .A1(net1571),
    .B1(_2753_),
    .X(_0469_));
 sg13g2_nand2_1 _6818_ (.Y(_2754_),
    .A(net1386),
    .B(_2749_));
 sg13g2_o21ai_1 _6819_ (.B1(_2754_),
    .Y(_0470_),
    .A1(net925),
    .A2(_2748_));
 sg13g2_nand2_1 _6820_ (.Y(_2755_),
    .A(net1293),
    .B(_2749_));
 sg13g2_o21ai_1 _6821_ (.B1(_2755_),
    .Y(_0471_),
    .A1(net922),
    .A2(_2748_));
 sg13g2_nand2_1 _6822_ (.Y(_2756_),
    .A(net1305),
    .B(_2749_));
 sg13g2_o21ai_1 _6823_ (.B1(_2756_),
    .Y(_0472_),
    .A1(net919),
    .A2(_2748_));
 sg13g2_nand2_1 _6824_ (.Y(_2757_),
    .A(net1224),
    .B(_2749_));
 sg13g2_o21ai_1 _6825_ (.B1(_2757_),
    .Y(_0473_),
    .A1(net917),
    .A2(_2748_));
 sg13g2_nand2b_2 _6826_ (.Y(_2758_),
    .B(_1158_),
    .A_N(_1137_));
 sg13g2_and2_1 _6827_ (.A(net1060),
    .B(net826),
    .X(_2759_));
 sg13g2_nand2_1 _6828_ (.Y(_2760_),
    .A(net1288),
    .B(_2759_));
 sg13g2_o21ai_1 _6829_ (.B1(_2760_),
    .Y(_0474_),
    .A1(net934),
    .A2(net826));
 sg13g2_nand2_1 _6830_ (.Y(_2761_),
    .A(net1252),
    .B(_2759_));
 sg13g2_o21ai_1 _6831_ (.B1(_2761_),
    .Y(_0475_),
    .A1(net933),
    .A2(net826));
 sg13g2_nand2_1 _6832_ (.Y(_2762_),
    .A(net789),
    .B(_2759_));
 sg13g2_o21ai_1 _6833_ (.B1(_2762_),
    .Y(_0476_),
    .A1(net930),
    .A2(net826));
 sg13g2_nand2_1 _6834_ (.Y(_2763_),
    .A(net805),
    .B(_2759_));
 sg13g2_o21ai_1 _6835_ (.B1(_2763_),
    .Y(_0477_),
    .A1(net926),
    .A2(net826));
 sg13g2_nand2_1 _6836_ (.Y(_2764_),
    .A(net1314),
    .B(_2759_));
 sg13g2_o21ai_1 _6837_ (.B1(_2764_),
    .Y(_0478_),
    .A1(net925),
    .A2(net826));
 sg13g2_nand2_1 _6838_ (.Y(_2765_),
    .A(net1289),
    .B(_2759_));
 sg13g2_o21ai_1 _6839_ (.B1(_2765_),
    .Y(_0479_),
    .A1(net921),
    .A2(net826));
 sg13g2_nand2_1 _6840_ (.Y(_2766_),
    .A(net808),
    .B(_2759_));
 sg13g2_o21ai_1 _6841_ (.B1(_2766_),
    .Y(_0480_),
    .A1(net919),
    .A2(_2758_));
 sg13g2_nand2_1 _6842_ (.Y(_2767_),
    .A(net818),
    .B(_2759_));
 sg13g2_o21ai_1 _6843_ (.B1(_2767_),
    .Y(_0481_),
    .A1(_1123_),
    .A2(net826));
 sg13g2_nor2_1 _6844_ (.A(\led_controller.led_effect_pulse.finished ),
    .B(\led_controller.effect_pulse_led_strb ),
    .Y(_2768_));
 sg13g2_nand4_1 _6845_ (.B(_0916_),
    .C(_1013_),
    .A(\led_controller.led_effect_pulse.calc_color_valid ),
    .Y(_2769_),
    .D(_2768_));
 sg13g2_nor2_2 _6846_ (.A(net1708),
    .B(_0919_),
    .Y(_2770_));
 sg13g2_nand2_2 _6847_ (.Y(_2771_),
    .A(_0918_),
    .B(_1013_));
 sg13g2_nand2_1 _6848_ (.Y(_2772_),
    .A(net1845),
    .B(_2771_));
 sg13g2_a21oi_1 _6849_ (.A1(net956),
    .A2(_2772_),
    .Y(_0482_),
    .B1(_0915_));
 sg13g2_o21ai_1 _6850_ (.B1(net989),
    .Y(_2773_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[0] ),
    .A2(net962));
 sg13g2_a21oi_1 _6851_ (.A1(_0793_),
    .A2(net962),
    .Y(_0483_),
    .B1(_2773_));
 sg13g2_o21ai_1 _6852_ (.B1(net988),
    .Y(_2774_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[1] ),
    .A2(net960));
 sg13g2_a21oi_1 _6853_ (.A1(_0792_),
    .A2(net960),
    .Y(_0484_),
    .B1(_2774_));
 sg13g2_o21ai_1 _6854_ (.B1(net985),
    .Y(_2775_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[2] ),
    .A2(net956));
 sg13g2_a21oi_1 _6855_ (.A1(_0791_),
    .A2(net956),
    .Y(_0485_),
    .B1(_2775_));
 sg13g2_o21ai_1 _6856_ (.B1(net986),
    .Y(_2776_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[3] ),
    .A2(net956));
 sg13g2_a21oi_1 _6857_ (.A1(_0790_),
    .A2(net956),
    .Y(_0486_),
    .B1(_2776_));
 sg13g2_o21ai_1 _6858_ (.B1(net987),
    .Y(_2777_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[4] ),
    .A2(net957));
 sg13g2_a21oi_1 _6859_ (.A1(_0789_),
    .A2(net957),
    .Y(_0487_),
    .B1(_2777_));
 sg13g2_o21ai_1 _6860_ (.B1(net988),
    .Y(_2778_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[5] ),
    .A2(net957));
 sg13g2_a21oi_1 _6861_ (.A1(_0788_),
    .A2(net957),
    .Y(_0488_),
    .B1(_2778_));
 sg13g2_o21ai_1 _6862_ (.B1(net988),
    .Y(_2779_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[6] ),
    .A2(net957));
 sg13g2_a21oi_1 _6863_ (.A1(_0787_),
    .A2(net957),
    .Y(_0489_),
    .B1(_2779_));
 sg13g2_o21ai_1 _6864_ (.B1(net987),
    .Y(_2780_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[7] ),
    .A2(net957));
 sg13g2_a21oi_1 _6865_ (.A1(_0786_),
    .A2(net959),
    .Y(_0490_),
    .B1(_2780_));
 sg13g2_o21ai_1 _6866_ (.B1(net990),
    .Y(_2781_),
    .A1(net1236),
    .A2(net961));
 sg13g2_a21oi_1 _6867_ (.A1(_0785_),
    .A2(net960),
    .Y(_0491_),
    .B1(_2781_));
 sg13g2_o21ai_1 _6868_ (.B1(net986),
    .Y(_2782_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[9] ),
    .A2(net956));
 sg13g2_a21oi_1 _6869_ (.A1(_0784_),
    .A2(_2769_),
    .Y(_0492_),
    .B1(_2782_));
 sg13g2_o21ai_1 _6870_ (.B1(net990),
    .Y(_2783_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[10] ),
    .A2(net961));
 sg13g2_a21oi_1 _6871_ (.A1(_0783_),
    .A2(net961),
    .Y(_0493_),
    .B1(_2783_));
 sg13g2_o21ai_1 _6872_ (.B1(net990),
    .Y(_2784_),
    .A1(net1320),
    .A2(net960));
 sg13g2_a21oi_1 _6873_ (.A1(_0782_),
    .A2(net960),
    .Y(_0494_),
    .B1(_2784_));
 sg13g2_o21ai_1 _6874_ (.B1(net989),
    .Y(_2785_),
    .A1(net1294),
    .A2(net960));
 sg13g2_a21oi_1 _6875_ (.A1(_0781_),
    .A2(net962),
    .Y(_0495_),
    .B1(_2785_));
 sg13g2_o21ai_1 _6876_ (.B1(net989),
    .Y(_2786_),
    .A1(net1411),
    .A2(net964));
 sg13g2_a21oi_1 _6877_ (.A1(_0780_),
    .A2(net964),
    .Y(_0496_),
    .B1(_2786_));
 sg13g2_o21ai_1 _6878_ (.B1(net989),
    .Y(_2787_),
    .A1(net1355),
    .A2(net962));
 sg13g2_a21oi_1 _6879_ (.A1(_0779_),
    .A2(net963),
    .Y(_0497_),
    .B1(_2787_));
 sg13g2_o21ai_1 _6880_ (.B1(net990),
    .Y(_2788_),
    .A1(net1358),
    .A2(net961));
 sg13g2_a21oi_1 _6881_ (.A1(_0778_),
    .A2(net962),
    .Y(_0498_),
    .B1(_2788_));
 sg13g2_o21ai_1 _6882_ (.B1(net989),
    .Y(_2789_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[16] ),
    .A2(net964));
 sg13g2_a21oi_1 _6883_ (.A1(_0777_),
    .A2(net964),
    .Y(_0499_),
    .B1(_2789_));
 sg13g2_o21ai_1 _6884_ (.B1(net990),
    .Y(_2790_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[17] ),
    .A2(net960));
 sg13g2_a21oi_1 _6885_ (.A1(_0776_),
    .A2(net960),
    .Y(_0500_),
    .B1(_2790_));
 sg13g2_o21ai_1 _6886_ (.B1(net990),
    .Y(_2791_),
    .A1(net1464),
    .A2(net961));
 sg13g2_a21oi_1 _6887_ (.A1(_0775_),
    .A2(net961),
    .Y(_0501_),
    .B1(_2791_));
 sg13g2_o21ai_1 _6888_ (.B1(net988),
    .Y(_2792_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[19] ),
    .A2(net956));
 sg13g2_a21oi_1 _6889_ (.A1(_0774_),
    .A2(net956),
    .Y(_0502_),
    .B1(_2792_));
 sg13g2_o21ai_1 _6890_ (.B1(net988),
    .Y(_2793_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[20] ),
    .A2(net957));
 sg13g2_a21oi_1 _6891_ (.A1(_0773_),
    .A2(net959),
    .Y(_0503_),
    .B1(_2793_));
 sg13g2_o21ai_1 _6892_ (.B1(net987),
    .Y(_2794_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[21] ),
    .A2(net958));
 sg13g2_a21oi_1 _6893_ (.A1(_0772_),
    .A2(net959),
    .Y(_0504_),
    .B1(_2794_));
 sg13g2_o21ai_1 _6894_ (.B1(net987),
    .Y(_2795_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[22] ),
    .A2(net958));
 sg13g2_a21oi_1 _6895_ (.A1(_0771_),
    .A2(net959),
    .Y(_0505_),
    .B1(_2795_));
 sg13g2_o21ai_1 _6896_ (.B1(net987),
    .Y(_2796_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[23] ),
    .A2(net964));
 sg13g2_a21oi_1 _6897_ (.A1(_0770_),
    .A2(net959),
    .Y(_0506_),
    .B1(_2796_));
 sg13g2_o21ai_1 _6898_ (.B1(net989),
    .Y(_2797_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[24] ),
    .A2(net962));
 sg13g2_a21oi_1 _6899_ (.A1(_0769_),
    .A2(net963),
    .Y(_0507_),
    .B1(_2797_));
 sg13g2_o21ai_1 _6900_ (.B1(net989),
    .Y(_2798_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[25] ),
    .A2(net962));
 sg13g2_a21oi_1 _6901_ (.A1(_0768_),
    .A2(net962),
    .Y(_0508_),
    .B1(_2798_));
 sg13g2_o21ai_1 _6902_ (.B1(net987),
    .Y(_2799_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[26] ),
    .A2(net958));
 sg13g2_a21oi_1 _6903_ (.A1(_0767_),
    .A2(net958),
    .Y(_0509_),
    .B1(_2799_));
 sg13g2_o21ai_1 _6904_ (.B1(net988),
    .Y(_2800_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[27] ),
    .A2(net965));
 sg13g2_a21oi_1 _6905_ (.A1(_0766_),
    .A2(net965),
    .Y(_0510_),
    .B1(_2800_));
 sg13g2_o21ai_1 _6906_ (.B1(net989),
    .Y(_2801_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[28] ),
    .A2(net963));
 sg13g2_a21oi_1 _6907_ (.A1(_0765_),
    .A2(net963),
    .Y(_0511_),
    .B1(_2801_));
 sg13g2_o21ai_1 _6908_ (.B1(net987),
    .Y(_2802_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[29] ),
    .A2(net958));
 sg13g2_a21oi_1 _6909_ (.A1(_0764_),
    .A2(net958),
    .Y(_0512_),
    .B1(_2802_));
 sg13g2_o21ai_1 _6910_ (.B1(net987),
    .Y(_2803_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[30] ),
    .A2(net958));
 sg13g2_a21oi_1 _6911_ (.A1(_0763_),
    .A2(net959),
    .Y(_0513_),
    .B1(_2803_));
 sg13g2_o21ai_1 _6912_ (.B1(net990),
    .Y(_2804_),
    .A1(\led_controller.led_effect_pulse.calc_color_out[31] ),
    .A2(net963));
 sg13g2_a21oi_1 _6913_ (.A1(_0762_),
    .A2(net963),
    .Y(_0514_),
    .B1(_2804_));
 sg13g2_nand2b_1 _6914_ (.Y(_2805_),
    .B(net2238),
    .A_N(_1014_));
 sg13g2_nor2_1 _6915_ (.A(\led_controller.led_effect_pulse.current_led[1] ),
    .B(_2708_),
    .Y(_2806_));
 sg13g2_o21ai_1 _6916_ (.B1(_2692_),
    .Y(_2807_),
    .A1(_0749_),
    .A2(\led_controller.led_effect_pulse.current_led[1] ));
 sg13g2_a21oi_1 _6917_ (.A1(_0761_),
    .A2(_2807_),
    .Y(_2808_),
    .B1(_2806_));
 sg13g2_o21ai_1 _6918_ (.B1(_2808_),
    .Y(_2809_),
    .A1(\led_controller.led_effect_pulse.current_led[2] ),
    .A2(_2705_));
 sg13g2_a22oi_1 _6919_ (.Y(_2810_),
    .B1(_2707_),
    .B2(\led_controller.led_effect_pulse.current_led[3] ),
    .A2(_2705_),
    .A1(\led_controller.led_effect_pulse.current_led[2] ));
 sg13g2_nor2_1 _6920_ (.A(\led_controller.led_effect_pulse.current_led[4] ),
    .B(_2703_),
    .Y(_2811_));
 sg13g2_a21oi_1 _6921_ (.A1(_2809_),
    .A2(_2810_),
    .Y(_2812_),
    .B1(_2811_));
 sg13g2_o21ai_1 _6922_ (.B1(_2812_),
    .Y(_2813_),
    .A1(\led_controller.led_effect_pulse.current_led[3] ),
    .A2(_2707_));
 sg13g2_a22oi_1 _6923_ (.Y(_2814_),
    .B1(_2703_),
    .B2(\led_controller.led_effect_pulse.current_led[4] ),
    .A2(_2701_),
    .A1(\led_controller.led_effect_pulse.current_led[5] ));
 sg13g2_nand2b_1 _6924_ (.Y(_2815_),
    .B(_2700_),
    .A_N(\led_controller.led_effect_pulse.current_led[5] ));
 sg13g2_o21ai_1 _6925_ (.B1(_2815_),
    .Y(_2816_),
    .A1(\led_controller.led_effect_pulse.current_led[6] ),
    .A2(_2699_));
 sg13g2_a21oi_1 _6926_ (.A1(_2813_),
    .A2(_2814_),
    .Y(_2817_),
    .B1(_2816_));
 sg13g2_a221oi_1 _6927_ (.B2(net1882),
    .C1(_2817_),
    .B1(_2699_),
    .A1(net1738),
    .Y(_2818_),
    .A2(_2698_));
 sg13g2_o21ai_1 _6928_ (.B1(_2770_),
    .Y(_2819_),
    .A1(net1738),
    .A2(_2698_));
 sg13g2_or3_1 _6929_ (.A(_2706_),
    .B(_2818_),
    .C(_2819_),
    .X(_2820_));
 sg13g2_a21oi_1 _6930_ (.A1(_2805_),
    .A2(_2820_),
    .Y(_0515_),
    .B1(_0915_));
 sg13g2_a21oi_1 _6931_ (.A1(net951),
    .A2(_2771_),
    .Y(_2821_),
    .B1(_0761_));
 sg13g2_o21ai_1 _6932_ (.B1(net985),
    .Y(_2822_),
    .A1(net1921),
    .A2(_2770_));
 sg13g2_nor2_1 _6933_ (.A(_2821_),
    .B(_2822_),
    .Y(_0516_));
 sg13g2_and2_1 _6934_ (.A(net1775),
    .B(_2821_),
    .X(_2823_));
 sg13g2_nand2_2 _6935_ (.Y(_2824_),
    .A(net985),
    .B(net951));
 sg13g2_nor2_1 _6936_ (.A(net1775),
    .B(_2821_),
    .Y(_2825_));
 sg13g2_nor3_1 _6937_ (.A(_2823_),
    .B(_2824_),
    .C(net1776),
    .Y(_0517_));
 sg13g2_and2_1 _6938_ (.A(net1860),
    .B(_2823_),
    .X(_2826_));
 sg13g2_or2_1 _6939_ (.X(_2827_),
    .B(_2826_),
    .A(_2824_));
 sg13g2_nor2_1 _6940_ (.A(net1860),
    .B(_2823_),
    .Y(_2828_));
 sg13g2_nor2_1 _6941_ (.A(_2827_),
    .B(net1861),
    .Y(_0518_));
 sg13g2_a21oi_1 _6942_ (.A1(_0918_),
    .A2(_2826_),
    .Y(_2829_),
    .B1(net1592));
 sg13g2_nand2b_1 _6943_ (.Y(_2830_),
    .B(net985),
    .A_N(net1592));
 sg13g2_a21oi_1 _6944_ (.A1(_2827_),
    .A2(_2830_),
    .Y(_0519_),
    .B1(net1593));
 sg13g2_a21oi_1 _6945_ (.A1(\led_controller.led_effect_pulse.current_led[3] ),
    .A2(_2826_),
    .Y(_2831_),
    .B1(net1580));
 sg13g2_and3_1 _6946_ (.X(_2832_),
    .A(net1580),
    .B(net1592),
    .C(_2826_));
 sg13g2_nor3_1 _6947_ (.A(_2824_),
    .B(net1581),
    .C(_2832_),
    .Y(_0520_));
 sg13g2_a22oi_1 _6948_ (.Y(_2833_),
    .B1(_2832_),
    .B2(_0918_),
    .A2(net951),
    .A1(net2147));
 sg13g2_and2_1 _6949_ (.A(net2147),
    .B(_2832_),
    .X(_2834_));
 sg13g2_nor3_1 _6950_ (.A(_0915_),
    .B(net2148),
    .C(_2834_),
    .Y(_0521_));
 sg13g2_nor2_1 _6951_ (.A(net1882),
    .B(_2834_),
    .Y(_2835_));
 sg13g2_and2_1 _6952_ (.A(net1882),
    .B(_2834_),
    .X(_2836_));
 sg13g2_nor3_1 _6953_ (.A(_2824_),
    .B(net1883),
    .C(_2836_),
    .Y(_0522_));
 sg13g2_nand4_1 _6954_ (.B(net985),
    .C(_0918_),
    .A(_0760_),
    .Y(_2837_),
    .D(_2836_));
 sg13g2_nand3_1 _6955_ (.B(net985),
    .C(net951),
    .A(net1738),
    .Y(_2838_));
 sg13g2_o21ai_1 _6956_ (.B1(_2837_),
    .Y(_0523_),
    .A1(_2836_),
    .A2(_2838_));
 sg13g2_xnor2_1 _6957_ (.Y(_2839_),
    .A(net2002),
    .B(_2677_));
 sg13g2_xor2_1 _6958_ (.B(net1736),
    .A(\led_controller.cpu.i_num_colors[0] ),
    .X(_2840_));
 sg13g2_a21oi_1 _6959_ (.A1(_2839_),
    .A2(_2840_),
    .Y(_2841_),
    .B1(_2771_));
 sg13g2_o21ai_1 _6960_ (.B1(net985),
    .Y(_2842_),
    .A1(net1736),
    .A2(_2841_));
 sg13g2_a21oi_1 _6961_ (.A1(net1736),
    .A2(_2770_),
    .Y(_0524_),
    .B1(_2842_));
 sg13g2_nand2_1 _6962_ (.Y(_2843_),
    .A(net2002),
    .B(_2771_));
 sg13g2_nor2b_2 _6963_ (.A(\led_controller.led_effect_pulse.color_index[0] ),
    .B_N(\led_controller.led_effect_pulse.color_index[1] ),
    .Y(_2844_));
 sg13g2_nor2b_2 _6964_ (.A(\led_controller.led_effect_pulse.color_index[1] ),
    .B_N(\led_controller.led_effect_pulse.color_index[0] ),
    .Y(_2845_));
 sg13g2_o21ai_1 _6965_ (.B1(_2841_),
    .Y(_2846_),
    .A1(net1090),
    .A2(net1085));
 sg13g2_a21oi_1 _6966_ (.A1(_2843_),
    .A2(_2846_),
    .Y(_0525_),
    .B1(_0915_));
 sg13g2_o21ai_1 _6967_ (.B1(_1015_),
    .Y(_2847_),
    .A1(net2283),
    .A2(_1018_));
 sg13g2_nor2_1 _6968_ (.A(net1175),
    .B(_1020_),
    .Y(_2848_));
 sg13g2_o21ai_1 _6969_ (.B1(net986),
    .Y(_2849_),
    .A1(_2847_),
    .A2(_2848_));
 sg13g2_a21oi_1 _6970_ (.A1(_2847_),
    .A2(_2848_),
    .Y(_0526_),
    .B1(_2849_));
 sg13g2_and2_1 _6971_ (.A(net1174),
    .B(net1175),
    .X(_2850_));
 sg13g2_nor2_1 _6972_ (.A(_1017_),
    .B(_2850_),
    .Y(_2851_));
 sg13g2_o21ai_1 _6973_ (.B1(net2283),
    .Y(_2852_),
    .A1(net1168),
    .A2(_1018_));
 sg13g2_nor2_1 _6974_ (.A(_2851_),
    .B(_2852_),
    .Y(_2853_));
 sg13g2_nor3_1 _6975_ (.A(net2283),
    .B(_1017_),
    .C(_2850_),
    .Y(_2854_));
 sg13g2_nor3_1 _6976_ (.A(net951),
    .B(_2853_),
    .C(_2854_),
    .Y(_2855_));
 sg13g2_o21ai_1 _6977_ (.B1(net986),
    .Y(_2856_),
    .A1(net1174),
    .A2(_1015_));
 sg13g2_nor2_1 _6978_ (.A(_2855_),
    .B(_2856_),
    .Y(_0527_));
 sg13g2_nor2_1 _6979_ (.A(_0882_),
    .B(_1017_),
    .Y(_2857_));
 sg13g2_nor2b_1 _6980_ (.A(_2850_),
    .B_N(_2852_),
    .Y(_2858_));
 sg13g2_nor3_1 _6981_ (.A(net951),
    .B(_2857_),
    .C(_2858_),
    .Y(_2859_));
 sg13g2_o21ai_1 _6982_ (.B1(net986),
    .Y(_2860_),
    .A1(net1172),
    .A2(_2859_));
 sg13g2_a21oi_1 _6983_ (.A1(net1172),
    .A2(_2859_),
    .Y(_0528_),
    .B1(_2860_));
 sg13g2_nand2_1 _6984_ (.Y(_2861_),
    .A(net1172),
    .B(_2850_));
 sg13g2_xnor2_1 _6985_ (.Y(_2862_),
    .A(net1170),
    .B(_2861_));
 sg13g2_a21o_1 _6986_ (.A2(_1017_),
    .A1(_0758_),
    .B1(_0757_),
    .X(_2863_));
 sg13g2_a21oi_1 _6987_ (.A1(_1018_),
    .A2(_2863_),
    .Y(_2864_),
    .B1(_2852_));
 sg13g2_a21oi_1 _6988_ (.A1(_0882_),
    .A2(_2862_),
    .Y(_2865_),
    .B1(_2864_));
 sg13g2_a21oi_1 _6989_ (.A1(net1170),
    .A2(_1016_),
    .Y(_2866_),
    .B1(_0915_));
 sg13g2_o21ai_1 _6990_ (.B1(_2866_),
    .Y(_0529_),
    .A1(_1016_),
    .A2(_2865_));
 sg13g2_nor4_1 _6991_ (.A(_0757_),
    .B(\led_controller.led_effect_pulse.fade_out ),
    .C(_1016_),
    .D(_2861_),
    .Y(_2867_));
 sg13g2_a21o_1 _6992_ (.A2(_1019_),
    .A1(\led_controller.led_effect_pulse.fade_out ),
    .B1(_2867_),
    .X(_2868_));
 sg13g2_o21ai_1 _6993_ (.B1(net986),
    .Y(_2869_),
    .A1(net1168),
    .A2(_2867_));
 sg13g2_a21oi_1 _6994_ (.A1(net1168),
    .A2(_2868_),
    .Y(_0530_),
    .B1(_2869_));
 sg13g2_a21oi_1 _6995_ (.A1(net2228),
    .A2(_0913_),
    .Y(_2870_),
    .B1(_0915_));
 sg13g2_nand2_1 _6996_ (.Y(_0531_),
    .A(_2771_),
    .B(net2229));
 sg13g2_nand2_2 _6997_ (.Y(_2871_),
    .A(net1159),
    .B(net1096));
 sg13g2_nand2b_2 _6998_ (.Y(_2872_),
    .B(net2228),
    .A_N(net1187));
 sg13g2_and2_1 _6999_ (.A(net1159),
    .B(net1082),
    .X(_2873_));
 sg13g2_nand2_2 _7000_ (.Y(_2874_),
    .A(net1159),
    .B(net1082));
 sg13g2_o21ai_1 _7001_ (.B1(_2871_),
    .Y(_0532_),
    .A1(_0887_),
    .A2(_2874_));
 sg13g2_a21oi_1 _7002_ (.A1(\led_controller.colors[43] ),
    .A2(net1085),
    .Y(_2875_),
    .B1(net1167));
 sg13g2_nor2_2 _7003_ (.A(\led_controller.led_effect_pulse.color_index[1] ),
    .B(\led_controller.led_effect_pulse.color_index[0] ),
    .Y(_2876_));
 sg13g2_a22oi_1 _7004_ (.Y(_2877_),
    .B1(net1079),
    .B2(\led_controller.colors[75] ),
    .A2(net1090),
    .A1(\led_controller.colors[11] ));
 sg13g2_a22oi_1 _7005_ (.Y(_2878_),
    .B1(net1081),
    .B2(\led_controller.colors[67] ),
    .A2(net1090),
    .A1(\led_controller.colors[3] ));
 sg13g2_a21oi_1 _7006_ (.A1(\led_controller.colors[35] ),
    .A2(net1085),
    .Y(_2879_),
    .B1(_0885_));
 sg13g2_a221oi_1 _7007_ (.B2(_2879_),
    .C1(_0902_),
    .B1(_2878_),
    .A1(_2875_),
    .Y(_2880_),
    .A2(_2877_));
 sg13g2_nor2_2 _7008_ (.A(net1165),
    .B(net1163),
    .Y(_2881_));
 sg13g2_or2_1 _7009_ (.X(_2882_),
    .B(net1163),
    .A(net1165));
 sg13g2_nand2_1 _7010_ (.Y(_2883_),
    .A(\led_controller.colors[27] ),
    .B(net1090));
 sg13g2_a22oi_1 _7011_ (.Y(_2884_),
    .B1(net1079),
    .B2(\led_controller.colors[91] ),
    .A2(net1085),
    .A1(\led_controller.colors[59] ));
 sg13g2_a21oi_1 _7012_ (.A1(_2883_),
    .A2(_2884_),
    .Y(_2885_),
    .B1(net1076));
 sg13g2_nor2_1 _7013_ (.A(_0885_),
    .B(net1163),
    .Y(_2886_));
 sg13g2_nand2b_2 _7014_ (.Y(_2887_),
    .B(net1167),
    .A_N(net1164));
 sg13g2_nand2_1 _7015_ (.Y(_2888_),
    .A(\led_controller.colors[83] ),
    .B(net1079));
 sg13g2_a22oi_1 _7016_ (.Y(_2889_),
    .B1(net1085),
    .B2(\led_controller.colors[51] ),
    .A2(net1090),
    .A1(\led_controller.colors[19] ));
 sg13g2_a21oi_1 _7017_ (.A1(_2888_),
    .A2(_2889_),
    .Y(_2890_),
    .B1(_2887_));
 sg13g2_or3_1 _7018_ (.A(_2880_),
    .B(_2885_),
    .C(_2890_),
    .X(_2891_));
 sg13g2_nand2_1 _7019_ (.Y(_2892_),
    .A(net1174),
    .B(_2891_));
 sg13g2_inv_1 _7020_ (.Y(_2893_),
    .A(_2892_));
 sg13g2_nand2_1 _7021_ (.Y(_2894_),
    .A(\led_controller.colors[88] ),
    .B(net1080));
 sg13g2_a22oi_1 _7022_ (.Y(_2895_),
    .B1(net1086),
    .B2(\led_controller.colors[56] ),
    .A2(net1091),
    .A1(\led_controller.colors[24] ));
 sg13g2_a21oi_1 _7023_ (.A1(_2894_),
    .A2(_2895_),
    .Y(_2896_),
    .B1(net1076));
 sg13g2_nor2b_2 _7024_ (.A(net1165),
    .B_N(net1163),
    .Y(_2897_));
 sg13g2_nand2b_2 _7025_ (.Y(_2898_),
    .B(net1164),
    .A_N(net1167));
 sg13g2_nor2_1 _7026_ (.A(net1014),
    .B(_2897_),
    .Y(_2899_));
 sg13g2_xor2_1 _7027_ (.B(net1164),
    .A(net1166),
    .X(_2900_));
 sg13g2_a22oi_1 _7028_ (.Y(_2901_),
    .B1(net1087),
    .B2(\led_controller.colors[32] ),
    .A2(net1091),
    .A1(\led_controller.colors[0] ));
 sg13g2_a21oi_1 _7029_ (.A1(\led_controller.colors[64] ),
    .A2(net1080),
    .Y(_2902_),
    .B1(_2900_));
 sg13g2_a21oi_1 _7030_ (.A1(\led_controller.colors[80] ),
    .A2(net1080),
    .Y(_2903_),
    .B1(net1164));
 sg13g2_a22oi_1 _7031_ (.Y(_2904_),
    .B1(net1086),
    .B2(\led_controller.colors[48] ),
    .A2(net1091),
    .A1(\led_controller.colors[16] ));
 sg13g2_a22oi_1 _7032_ (.Y(_2905_),
    .B1(net1087),
    .B2(\led_controller.colors[40] ),
    .A2(net1092),
    .A1(\led_controller.colors[8] ));
 sg13g2_a21oi_1 _7033_ (.A1(\led_controller.colors[72] ),
    .A2(net1080),
    .Y(_2906_),
    .B1(net1166));
 sg13g2_a21oi_1 _7034_ (.A1(_2901_),
    .A2(_2902_),
    .Y(_2907_),
    .B1(_2881_));
 sg13g2_a22oi_1 _7035_ (.Y(_2908_),
    .B1(_2905_),
    .B2(_2906_),
    .A2(_2904_),
    .A1(_2903_));
 sg13g2_a21o_2 _7036_ (.A2(_2908_),
    .A1(_2907_),
    .B1(_2896_),
    .X(_2909_));
 sg13g2_nand2_1 _7037_ (.Y(_2910_),
    .A(net1170),
    .B(_2909_));
 sg13g2_inv_1 _7038_ (.Y(_2911_),
    .A(_2910_));
 sg13g2_nand2_1 _7039_ (.Y(_2912_),
    .A(net1175),
    .B(_2891_));
 sg13g2_inv_1 _7040_ (.Y(_2913_),
    .A(_2912_));
 sg13g2_a21oi_1 _7041_ (.A1(\led_controller.colors[41] ),
    .A2(net1085),
    .Y(_2914_),
    .B1(net1166));
 sg13g2_a22oi_1 _7042_ (.Y(_2915_),
    .B1(net1081),
    .B2(\led_controller.colors[73] ),
    .A2(net1090),
    .A1(\led_controller.colors[9] ));
 sg13g2_a22oi_1 _7043_ (.Y(_2916_),
    .B1(net1079),
    .B2(\led_controller.colors[65] ),
    .A2(net1090),
    .A1(\led_controller.colors[1] ));
 sg13g2_a21oi_1 _7044_ (.A1(\led_controller.colors[33] ),
    .A2(net1087),
    .Y(_2917_),
    .B1(_0885_));
 sg13g2_a221oi_1 _7045_ (.B2(_2917_),
    .C1(_0902_),
    .B1(_2916_),
    .A1(_2914_),
    .Y(_2918_),
    .A2(_2915_));
 sg13g2_nand2_1 _7046_ (.Y(_2919_),
    .A(\led_controller.colors[25] ),
    .B(net1090));
 sg13g2_a22oi_1 _7047_ (.Y(_2920_),
    .B1(net1079),
    .B2(\led_controller.colors[89] ),
    .A2(net1085),
    .A1(\led_controller.colors[57] ));
 sg13g2_a21oi_1 _7048_ (.A1(_2919_),
    .A2(_2920_),
    .Y(_2921_),
    .B1(_2882_));
 sg13g2_nand2_1 _7049_ (.Y(_2922_),
    .A(\led_controller.colors[81] ),
    .B(net1079));
 sg13g2_a22oi_1 _7050_ (.Y(_2923_),
    .B1(net1085),
    .B2(\led_controller.colors[49] ),
    .A2(net1092),
    .A1(\led_controller.colors[17] ));
 sg13g2_a21oi_1 _7051_ (.A1(_2922_),
    .A2(_2923_),
    .Y(_2924_),
    .B1(_2887_));
 sg13g2_or3_1 _7052_ (.A(_2918_),
    .B(_2921_),
    .C(_2924_),
    .X(_2925_));
 sg13g2_nand2_1 _7053_ (.Y(_2926_),
    .A(net1172),
    .B(_2925_));
 sg13g2_nor2_1 _7054_ (.A(_2912_),
    .B(_2926_),
    .Y(_2927_));
 sg13g2_xor2_1 _7055_ (.B(_2926_),
    .A(_2912_),
    .X(_2928_));
 sg13g2_xnor2_1 _7056_ (.Y(_2929_),
    .A(_2910_),
    .B(_2928_));
 sg13g2_a21oi_1 _7057_ (.A1(\led_controller.colors[10] ),
    .A2(net1091),
    .Y(_2930_),
    .B1(_2898_));
 sg13g2_a22oi_1 _7058_ (.Y(_2931_),
    .B1(net1079),
    .B2(\led_controller.colors[74] ),
    .A2(net1086),
    .A1(\led_controller.colors[42] ));
 sg13g2_a21oi_1 _7059_ (.A1(\led_controller.colors[2] ),
    .A2(net1091),
    .Y(_2932_),
    .B1(_2897_));
 sg13g2_a22oi_1 _7060_ (.Y(_2933_),
    .B1(net1079),
    .B2(\led_controller.colors[66] ),
    .A2(net1086),
    .A1(\led_controller.colors[34] ));
 sg13g2_a22oi_1 _7061_ (.Y(_2934_),
    .B1(_2932_),
    .B2(_2933_),
    .A2(_2931_),
    .A1(_2930_));
 sg13g2_nor2_1 _7062_ (.A(_0902_),
    .B(_2934_),
    .Y(_2935_));
 sg13g2_a22oi_1 _7063_ (.Y(_2936_),
    .B1(net1086),
    .B2(\led_controller.colors[58] ),
    .A2(net1091),
    .A1(\led_controller.colors[26] ));
 sg13g2_a21oi_1 _7064_ (.A1(\led_controller.colors[90] ),
    .A2(net1081),
    .Y(_2937_),
    .B1(_2882_));
 sg13g2_a22oi_1 _7065_ (.Y(_2938_),
    .B1(net1087),
    .B2(\led_controller.colors[50] ),
    .A2(net1092),
    .A1(\led_controller.colors[18] ));
 sg13g2_a21oi_1 _7066_ (.A1(\led_controller.colors[82] ),
    .A2(net1080),
    .Y(_2939_),
    .B1(_2887_));
 sg13g2_a22oi_1 _7067_ (.Y(_2940_),
    .B1(_2938_),
    .B2(_2939_),
    .A2(_2937_),
    .A1(_2936_));
 sg13g2_nor2b_2 _7068_ (.A(_2935_),
    .B_N(_2940_),
    .Y(_2941_));
 sg13g2_o21ai_1 _7069_ (.B1(_2940_),
    .Y(_2942_),
    .A1(_0902_),
    .A2(_2934_));
 sg13g2_nor2_1 _7070_ (.A(_0759_),
    .B(_2942_),
    .Y(_2943_));
 sg13g2_nand2_1 _7071_ (.Y(_2944_),
    .A(net1172),
    .B(_2909_));
 sg13g2_nor3_1 _7072_ (.A(_0759_),
    .B(_2942_),
    .C(_2944_),
    .Y(_2945_));
 sg13g2_and2_1 _7073_ (.A(_2929_),
    .B(_2945_),
    .X(_2946_));
 sg13g2_and2_1 _7074_ (.A(net1168),
    .B(_2909_),
    .X(_2947_));
 sg13g2_a21oi_1 _7075_ (.A1(_2911_),
    .A2(_2928_),
    .Y(_2948_),
    .B1(_2927_));
 sg13g2_nand2_1 _7076_ (.Y(_2949_),
    .A(net1170),
    .B(_2925_));
 sg13g2_a21oi_1 _7077_ (.A1(\led_controller.colors[12] ),
    .A2(net1089),
    .Y(_2950_),
    .B1(_2898_));
 sg13g2_a22oi_1 _7078_ (.Y(_2951_),
    .B1(net1078),
    .B2(\led_controller.colors[76] ),
    .A2(net1084),
    .A1(\led_controller.colors[44] ));
 sg13g2_a21oi_1 _7079_ (.A1(\led_controller.colors[4] ),
    .A2(net1089),
    .Y(_2952_),
    .B1(_2897_));
 sg13g2_a22oi_1 _7080_ (.Y(_2953_),
    .B1(net1080),
    .B2(\led_controller.colors[68] ),
    .A2(net1086),
    .A1(\led_controller.colors[36] ));
 sg13g2_a22oi_1 _7081_ (.Y(_2954_),
    .B1(_2952_),
    .B2(_2953_),
    .A2(_2951_),
    .A1(_2950_));
 sg13g2_nand2b_1 _7082_ (.Y(_2955_),
    .B(net1163),
    .A_N(_2954_));
 sg13g2_a22oi_1 _7083_ (.Y(_2956_),
    .B1(net1086),
    .B2(\led_controller.colors[60] ),
    .A2(net1091),
    .A1(\led_controller.colors[28] ));
 sg13g2_a21oi_1 _7084_ (.A1(\led_controller.colors[92] ),
    .A2(net1080),
    .Y(_2957_),
    .B1(net1076));
 sg13g2_a22oi_1 _7085_ (.Y(_2958_),
    .B1(net1086),
    .B2(\led_controller.colors[52] ),
    .A2(net1091),
    .A1(\led_controller.colors[20] ));
 sg13g2_a21oi_1 _7086_ (.A1(\led_controller.colors[84] ),
    .A2(net1080),
    .Y(_2959_),
    .B1(_2887_));
 sg13g2_a22oi_1 _7087_ (.Y(_2960_),
    .B1(_2958_),
    .B2(_2959_),
    .A2(_2957_),
    .A1(_2956_));
 sg13g2_and2_1 _7088_ (.A(_2955_),
    .B(_2960_),
    .X(_2961_));
 sg13g2_nand2_1 _7089_ (.Y(_2962_),
    .A(net1172),
    .B(_2961_));
 sg13g2_and3_1 _7090_ (.X(_2963_),
    .A(net1175),
    .B(_2955_),
    .C(_2960_));
 sg13g2_nor2_1 _7091_ (.A(_0758_),
    .B(_2942_),
    .Y(_2964_));
 sg13g2_nand2_1 _7092_ (.Y(_2965_),
    .A(_2963_),
    .B(_2964_));
 sg13g2_xnor2_1 _7093_ (.Y(_2966_),
    .A(_2963_),
    .B(_2964_));
 sg13g2_xnor2_1 _7094_ (.Y(_2967_),
    .A(_2949_),
    .B(_2966_));
 sg13g2_nor2_1 _7095_ (.A(_2948_),
    .B(_2967_),
    .Y(_2968_));
 sg13g2_xor2_1 _7096_ (.B(_2967_),
    .A(_2948_),
    .X(_2969_));
 sg13g2_xor2_1 _7097_ (.B(_2969_),
    .A(_2947_),
    .X(_2970_));
 sg13g2_and2_1 _7098_ (.A(_2946_),
    .B(_2970_),
    .X(_2971_));
 sg13g2_xor2_1 _7099_ (.B(_2970_),
    .A(_2946_),
    .X(_2972_));
 sg13g2_xnor2_1 _7100_ (.Y(_2973_),
    .A(_2892_),
    .B(_2972_));
 sg13g2_xor2_1 _7101_ (.B(_2945_),
    .A(_2929_),
    .X(_2974_));
 sg13g2_and3_2 _7102_ (.X(_2975_),
    .A(net1174),
    .B(_2941_),
    .C(_2974_));
 sg13g2_and2_1 _7103_ (.A(_2973_),
    .B(_2975_),
    .X(_2976_));
 sg13g2_xnor2_1 _7104_ (.Y(_2977_),
    .A(_2973_),
    .B(_2975_));
 sg13g2_xnor2_1 _7105_ (.Y(_2978_),
    .A(_2943_),
    .B(_2944_));
 sg13g2_o21ai_1 _7106_ (.B1(net1174),
    .Y(_2979_),
    .A1(_2929_),
    .A2(_2941_));
 sg13g2_o21ai_1 _7107_ (.B1(_2978_),
    .Y(_2980_),
    .A1(_2975_),
    .A2(_2979_));
 sg13g2_nand3_1 _7108_ (.B(_2909_),
    .C(_2929_),
    .A(_2850_),
    .Y(_2981_));
 sg13g2_nand2b_1 _7109_ (.Y(_2982_),
    .B(_2981_),
    .A_N(_2978_));
 sg13g2_nand3_1 _7110_ (.B(_2980_),
    .C(_2982_),
    .A(_2925_),
    .Y(_2983_));
 sg13g2_nor2_1 _7111_ (.A(_2977_),
    .B(_2983_),
    .Y(_2984_));
 sg13g2_xnor2_1 _7112_ (.Y(_2985_),
    .A(_2977_),
    .B(_2983_));
 sg13g2_o21ai_1 _7113_ (.B1(net1015),
    .Y(_2986_),
    .A1(net1898),
    .A2(net1096));
 sg13g2_a21oi_1 _7114_ (.A1(net1096),
    .A2(_2985_),
    .Y(_0533_),
    .B1(_2986_));
 sg13g2_nor2_1 _7115_ (.A(_2976_),
    .B(_2984_),
    .Y(_2987_));
 sg13g2_a21oi_1 _7116_ (.A1(_2893_),
    .A2(_2972_),
    .Y(_2988_),
    .B1(_2971_));
 sg13g2_and2_1 _7117_ (.A(net1174),
    .B(_2961_),
    .X(_2989_));
 sg13g2_a21oi_1 _7118_ (.A1(_2947_),
    .A2(_2969_),
    .Y(_2990_),
    .B1(_2968_));
 sg13g2_nand2_1 _7119_ (.Y(_2991_),
    .A(net1168),
    .B(_2925_));
 sg13g2_o21ai_1 _7120_ (.B1(_2965_),
    .Y(_2992_),
    .A1(_2949_),
    .A2(_2966_));
 sg13g2_nand2_1 _7121_ (.Y(_2993_),
    .A(net1170),
    .B(_2941_));
 sg13g2_a21oi_1 _7122_ (.A1(\led_controller.colors[13] ),
    .A2(net1088),
    .Y(_2994_),
    .B1(_2898_));
 sg13g2_a22oi_1 _7123_ (.Y(_2995_),
    .B1(net1077),
    .B2(\led_controller.colors[77] ),
    .A2(net1083),
    .A1(\led_controller.colors[45] ));
 sg13g2_a21oi_1 _7124_ (.A1(\led_controller.colors[5] ),
    .A2(net1088),
    .Y(_2996_),
    .B1(_2897_));
 sg13g2_a22oi_1 _7125_ (.Y(_2997_),
    .B1(net1077),
    .B2(\led_controller.colors[69] ),
    .A2(net1083),
    .A1(\led_controller.colors[37] ));
 sg13g2_a22oi_1 _7126_ (.Y(_2998_),
    .B1(_2996_),
    .B2(_2997_),
    .A2(_2995_),
    .A1(_2994_));
 sg13g2_nand2b_1 _7127_ (.Y(_2999_),
    .B(net1163),
    .A_N(_2998_));
 sg13g2_a22oi_1 _7128_ (.Y(_3000_),
    .B1(net1083),
    .B2(\led_controller.colors[53] ),
    .A2(net1088),
    .A1(\led_controller.colors[21] ));
 sg13g2_a21oi_1 _7129_ (.A1(\led_controller.colors[85] ),
    .A2(net1077),
    .Y(_3001_),
    .B1(_2887_));
 sg13g2_a22oi_1 _7130_ (.Y(_3002_),
    .B1(net1083),
    .B2(\led_controller.colors[61] ),
    .A2(net1088),
    .A1(\led_controller.colors[29] ));
 sg13g2_a21oi_1 _7131_ (.A1(\led_controller.colors[93] ),
    .A2(net1077),
    .Y(_3003_),
    .B1(net1076));
 sg13g2_a22oi_1 _7132_ (.Y(_3004_),
    .B1(_3002_),
    .B2(_3003_),
    .A2(_3001_),
    .A1(_3000_));
 sg13g2_and2_1 _7133_ (.A(_2999_),
    .B(_3004_),
    .X(_3005_));
 sg13g2_and2_1 _7134_ (.A(net1172),
    .B(_3005_),
    .X(_3006_));
 sg13g2_and3_1 _7135_ (.X(_3007_),
    .A(net1175),
    .B(_2999_),
    .C(_3004_));
 sg13g2_nand2_1 _7136_ (.Y(_3008_),
    .A(net1173),
    .B(_2891_));
 sg13g2_xor2_1 _7137_ (.B(_3008_),
    .A(_3007_),
    .X(_3009_));
 sg13g2_nor2_1 _7138_ (.A(_2993_),
    .B(_3009_),
    .Y(_3010_));
 sg13g2_xnor2_1 _7139_ (.Y(_3011_),
    .A(_2993_),
    .B(_3009_));
 sg13g2_nand2b_1 _7140_ (.Y(_3012_),
    .B(_2992_),
    .A_N(_3011_));
 sg13g2_xor2_1 _7141_ (.B(_3011_),
    .A(_2992_),
    .X(_3013_));
 sg13g2_xnor2_1 _7142_ (.Y(_3014_),
    .A(_2991_),
    .B(_3013_));
 sg13g2_nor2_1 _7143_ (.A(_2990_),
    .B(_3014_),
    .Y(_3015_));
 sg13g2_xor2_1 _7144_ (.B(_3014_),
    .A(_2990_),
    .X(_3016_));
 sg13g2_xnor2_1 _7145_ (.Y(_3017_),
    .A(_2989_),
    .B(_3016_));
 sg13g2_nor2_1 _7146_ (.A(_2988_),
    .B(_3017_),
    .Y(_3018_));
 sg13g2_nand2_1 _7147_ (.Y(_3019_),
    .A(_2988_),
    .B(_3017_));
 sg13g2_nor2b_1 _7148_ (.A(_3018_),
    .B_N(_3019_),
    .Y(_3020_));
 sg13g2_xor2_1 _7149_ (.B(_3020_),
    .A(_2987_),
    .X(_3021_));
 sg13g2_o21ai_1 _7150_ (.B1(net1015),
    .Y(_3022_),
    .A1(net1944),
    .A2(net1096));
 sg13g2_a21oi_1 _7151_ (.A1(net1096),
    .A2(_3021_),
    .Y(_0534_),
    .B1(_3022_));
 sg13g2_or2_1 _7152_ (.X(_3023_),
    .B(_3018_),
    .A(_2976_));
 sg13g2_a22oi_1 _7153_ (.Y(_3024_),
    .B1(_3023_),
    .B2(_3019_),
    .A2(_3020_),
    .A1(_2984_));
 sg13g2_a21oi_1 _7154_ (.A1(_2989_),
    .A2(_3016_),
    .Y(_3025_),
    .B1(_3015_));
 sg13g2_nand2_1 _7155_ (.Y(_3026_),
    .A(net1174),
    .B(_3005_));
 sg13g2_o21ai_1 _7156_ (.B1(_3012_),
    .Y(_3027_),
    .A1(_2991_),
    .A2(_3013_));
 sg13g2_and2_1 _7157_ (.A(net1168),
    .B(_2941_),
    .X(_3028_));
 sg13g2_a21oi_1 _7158_ (.A1(_2913_),
    .A2(_3006_),
    .Y(_3029_),
    .B1(_3010_));
 sg13g2_nand2_1 _7159_ (.Y(_3030_),
    .A(net1170),
    .B(_2891_));
 sg13g2_nand2_1 _7160_ (.Y(_3031_),
    .A(\led_controller.colors[94] ),
    .B(net1077));
 sg13g2_a22oi_1 _7161_ (.Y(_3032_),
    .B1(net1083),
    .B2(\led_controller.colors[62] ),
    .A2(net1088),
    .A1(\led_controller.colors[30] ));
 sg13g2_a21oi_1 _7162_ (.A1(_3031_),
    .A2(_3032_),
    .Y(_3033_),
    .B1(net1076));
 sg13g2_a21oi_1 _7163_ (.A1(\led_controller.colors[70] ),
    .A2(net1077),
    .Y(_3034_),
    .B1(_2900_));
 sg13g2_a22oi_1 _7164_ (.Y(_3035_),
    .B1(net1083),
    .B2(\led_controller.colors[38] ),
    .A2(net1088),
    .A1(\led_controller.colors[6] ));
 sg13g2_a21oi_1 _7165_ (.A1(_3034_),
    .A2(_3035_),
    .Y(_3036_),
    .B1(_2881_));
 sg13g2_a22oi_1 _7166_ (.Y(_3037_),
    .B1(net1084),
    .B2(\led_controller.colors[54] ),
    .A2(net1089),
    .A1(\led_controller.colors[22] ));
 sg13g2_a21oi_1 _7167_ (.A1(\led_controller.colors[86] ),
    .A2(net1078),
    .Y(_3038_),
    .B1(net1164));
 sg13g2_a22oi_1 _7168_ (.Y(_3039_),
    .B1(net1084),
    .B2(\led_controller.colors[46] ),
    .A2(net1089),
    .A1(\led_controller.colors[14] ));
 sg13g2_a21oi_1 _7169_ (.A1(\led_controller.colors[78] ),
    .A2(net1078),
    .Y(_3040_),
    .B1(net1167));
 sg13g2_a22oi_1 _7170_ (.Y(_3041_),
    .B1(_3039_),
    .B2(_3040_),
    .A2(_3038_),
    .A1(_3037_));
 sg13g2_a21o_2 _7171_ (.A2(_3041_),
    .A1(_3036_),
    .B1(_3033_),
    .X(_3042_));
 sg13g2_nand2_1 _7172_ (.Y(_3043_),
    .A(net1173),
    .B(_3042_));
 sg13g2_nand2_1 _7173_ (.Y(_3044_),
    .A(net1175),
    .B(_3042_));
 sg13g2_xnor2_1 _7174_ (.Y(_3045_),
    .A(_2962_),
    .B(_3044_));
 sg13g2_or2_1 _7175_ (.X(_3046_),
    .B(_3045_),
    .A(_3030_));
 sg13g2_xor2_1 _7176_ (.B(_3045_),
    .A(_3030_),
    .X(_3047_));
 sg13g2_nor2b_1 _7177_ (.A(_3029_),
    .B_N(_3047_),
    .Y(_3048_));
 sg13g2_xnor2_1 _7178_ (.Y(_3049_),
    .A(_3029_),
    .B(_3047_));
 sg13g2_xnor2_1 _7179_ (.Y(_3050_),
    .A(_3028_),
    .B(_3049_));
 sg13g2_nor2b_1 _7180_ (.A(_3050_),
    .B_N(_3027_),
    .Y(_3051_));
 sg13g2_xor2_1 _7181_ (.B(_3050_),
    .A(_3027_),
    .X(_3052_));
 sg13g2_nor2_1 _7182_ (.A(_3026_),
    .B(_3052_),
    .Y(_3053_));
 sg13g2_xnor2_1 _7183_ (.Y(_3054_),
    .A(_3026_),
    .B(_3052_));
 sg13g2_or2_1 _7184_ (.X(_3055_),
    .B(_3054_),
    .A(_3025_));
 sg13g2_and2_1 _7185_ (.A(_3025_),
    .B(_3054_),
    .X(_3056_));
 sg13g2_xor2_1 _7186_ (.B(_3054_),
    .A(_3025_),
    .X(_3057_));
 sg13g2_xnor2_1 _7187_ (.Y(_3058_),
    .A(_3024_),
    .B(_3057_));
 sg13g2_nand2b_1 _7188_ (.Y(_3059_),
    .B(_3058_),
    .A_N(_1519_));
 sg13g2_nand2_2 _7189_ (.Y(_3060_),
    .A(net1187),
    .B(net1076));
 sg13g2_nand2_1 _7190_ (.Y(_3061_),
    .A(net1879),
    .B(net1082));
 sg13g2_nand3_1 _7191_ (.B(_1519_),
    .C(net1082),
    .A(net1879),
    .Y(_3062_));
 sg13g2_nor2b_1 _7192_ (.A(_3060_),
    .B_N(_3062_),
    .Y(_3063_));
 sg13g2_a221oi_1 _7193_ (.B2(_3059_),
    .C1(net1131),
    .B1(_3063_),
    .A1(_3060_),
    .Y(_0535_),
    .A2(net1880));
 sg13g2_and2_1 _7194_ (.A(net2366),
    .B(net1082),
    .X(_3064_));
 sg13g2_nand2_1 _7195_ (.Y(_3065_),
    .A(_2900_),
    .B(_3064_));
 sg13g2_o21ai_1 _7196_ (.B1(_3055_),
    .Y(_3066_),
    .A1(_3024_),
    .A2(_3056_));
 sg13g2_nor2_1 _7197_ (.A(_3051_),
    .B(_3053_),
    .Y(_3067_));
 sg13g2_nand2_1 _7198_ (.Y(_3068_),
    .A(\led_controller.led_effect_pulse.brightness[1] ),
    .B(_3042_));
 sg13g2_a21o_1 _7199_ (.A2(_3049_),
    .A1(_3028_),
    .B1(_3048_),
    .X(_3069_));
 sg13g2_nand2_1 _7200_ (.Y(_3070_),
    .A(net1168),
    .B(_2891_));
 sg13g2_o21ai_1 _7201_ (.B1(_3046_),
    .Y(_3071_),
    .A1(_2962_),
    .A2(_3044_));
 sg13g2_nand2_1 _7202_ (.Y(_3072_),
    .A(net1170),
    .B(_2961_));
 sg13g2_a22oi_1 _7203_ (.Y(_3073_),
    .B1(net1078),
    .B2(\led_controller.colors[87] ),
    .A2(net1089),
    .A1(\led_controller.colors[23] ));
 sg13g2_a21oi_1 _7204_ (.A1(\led_controller.colors[55] ),
    .A2(net1083),
    .Y(_3074_),
    .B1(_2887_));
 sg13g2_a21oi_1 _7205_ (.A1(\led_controller.colors[15] ),
    .A2(net1088),
    .Y(_3075_),
    .B1(_2898_));
 sg13g2_a22oi_1 _7206_ (.Y(_3076_),
    .B1(net1078),
    .B2(\led_controller.colors[79] ),
    .A2(net1084),
    .A1(\led_controller.colors[47] ));
 sg13g2_nand2_1 _7207_ (.Y(_3077_),
    .A(_3075_),
    .B(_3076_));
 sg13g2_a21oi_1 _7208_ (.A1(\led_controller.colors[71] ),
    .A2(net1077),
    .Y(_3078_),
    .B1(_2900_));
 sg13g2_a22oi_1 _7209_ (.Y(_3079_),
    .B1(net1084),
    .B2(\led_controller.colors[39] ),
    .A2(net1089),
    .A1(\led_controller.colors[7] ));
 sg13g2_a22oi_1 _7210_ (.Y(_3080_),
    .B1(net1077),
    .B2(\led_controller.colors[95] ),
    .A2(net1083),
    .A1(\led_controller.colors[63] ));
 sg13g2_a21oi_1 _7211_ (.A1(\led_controller.colors[31] ),
    .A2(net1088),
    .Y(_3081_),
    .B1(net1076));
 sg13g2_a22oi_1 _7212_ (.Y(_3082_),
    .B1(_3078_),
    .B2(_3079_),
    .A2(_3074_),
    .A1(_3073_));
 sg13g2_nand2_1 _7213_ (.Y(_3083_),
    .A(_3077_),
    .B(_3082_));
 sg13g2_a22oi_1 _7214_ (.Y(_3084_),
    .B1(_3083_),
    .B2(net1076),
    .A2(_3081_),
    .A1(_3080_));
 sg13g2_and2_1 _7215_ (.A(net1173),
    .B(_3084_),
    .X(_3085_));
 sg13g2_nand2_1 _7216_ (.Y(_3086_),
    .A(net1173),
    .B(_3084_));
 sg13g2_nand2_1 _7217_ (.Y(_3087_),
    .A(\led_controller.led_effect_pulse.brightness[0] ),
    .B(_3084_));
 sg13g2_xor2_1 _7218_ (.B(_3087_),
    .A(_3006_),
    .X(_3088_));
 sg13g2_nor2_1 _7219_ (.A(_3072_),
    .B(_3088_),
    .Y(_3089_));
 sg13g2_xnor2_1 _7220_ (.Y(_3090_),
    .A(_3072_),
    .B(_3088_));
 sg13g2_nand2b_1 _7221_ (.Y(_3091_),
    .B(_3071_),
    .A_N(_3090_));
 sg13g2_xor2_1 _7222_ (.B(_3090_),
    .A(_3071_),
    .X(_3092_));
 sg13g2_xor2_1 _7223_ (.B(_3092_),
    .A(_3070_),
    .X(_3093_));
 sg13g2_xor2_1 _7224_ (.B(_3093_),
    .A(_3069_),
    .X(_3094_));
 sg13g2_nor2b_1 _7225_ (.A(_3068_),
    .B_N(_3094_),
    .Y(_3095_));
 sg13g2_xnor2_1 _7226_ (.Y(_3096_),
    .A(_3068_),
    .B(_3094_));
 sg13g2_nor2b_1 _7227_ (.A(_3067_),
    .B_N(_3096_),
    .Y(_3097_));
 sg13g2_xnor2_1 _7228_ (.Y(_3098_),
    .A(_3067_),
    .B(_3096_));
 sg13g2_xnor2_1 _7229_ (.Y(_3099_),
    .A(_3066_),
    .B(_3098_));
 sg13g2_o21ai_1 _7230_ (.B1(_3065_),
    .Y(_3100_),
    .A1(_1519_),
    .A2(_3099_));
 sg13g2_a22oi_1 _7231_ (.Y(_3101_),
    .B1(_3100_),
    .B2(net1187),
    .A2(_3064_),
    .A1(_3060_));
 sg13g2_nor2_1 _7232_ (.A(net1128),
    .B(net2367),
    .Y(_0536_));
 sg13g2_a21oi_1 _7233_ (.A1(_3066_),
    .A2(_3098_),
    .Y(_3102_),
    .B1(_3097_));
 sg13g2_a21o_1 _7234_ (.A2(_3093_),
    .A1(_3069_),
    .B1(_3095_),
    .X(_3103_));
 sg13g2_nand2_1 _7235_ (.Y(_3104_),
    .A(\led_controller.led_effect_pulse.brightness[1] ),
    .B(_3084_));
 sg13g2_o21ai_1 _7236_ (.B1(_3091_),
    .Y(_3105_),
    .A1(_3070_),
    .A2(_3092_));
 sg13g2_and2_1 _7237_ (.A(net1169),
    .B(_2961_),
    .X(_3106_));
 sg13g2_nand2_1 _7238_ (.Y(_3107_),
    .A(net1171),
    .B(_3042_));
 sg13g2_nand2_1 _7239_ (.Y(_3108_),
    .A(net1171),
    .B(_3005_));
 sg13g2_xor2_1 _7240_ (.B(_3108_),
    .A(_3043_),
    .X(_3109_));
 sg13g2_a21oi_1 _7241_ (.A1(_3007_),
    .A2(_3085_),
    .Y(_3110_),
    .B1(_3089_));
 sg13g2_nor2b_1 _7242_ (.A(_3110_),
    .B_N(_3109_),
    .Y(_3111_));
 sg13g2_xnor2_1 _7243_ (.Y(_3112_),
    .A(_3109_),
    .B(_3110_));
 sg13g2_xnor2_1 _7244_ (.Y(_3113_),
    .A(_3106_),
    .B(_3112_));
 sg13g2_nand2b_1 _7245_ (.Y(_3114_),
    .B(_3105_),
    .A_N(_3113_));
 sg13g2_xor2_1 _7246_ (.B(_3113_),
    .A(_3105_),
    .X(_3115_));
 sg13g2_xor2_1 _7247_ (.B(_3115_),
    .A(_3104_),
    .X(_3116_));
 sg13g2_nand2_1 _7248_ (.Y(_3117_),
    .A(_3103_),
    .B(_3116_));
 sg13g2_xnor2_1 _7249_ (.Y(_3118_),
    .A(_3103_),
    .B(_3116_));
 sg13g2_xnor2_1 _7250_ (.Y(_3119_),
    .A(_3102_),
    .B(_3118_));
 sg13g2_nand2_1 _7251_ (.Y(_3120_),
    .A(net1540),
    .B(net1015));
 sg13g2_a22oi_1 _7252_ (.Y(_0537_),
    .B1(_3120_),
    .B2(_2871_),
    .A2(_3119_),
    .A1(net1096));
 sg13g2_a21oi_1 _7253_ (.A1(_3106_),
    .A2(_3112_),
    .Y(_3121_),
    .B1(_3111_));
 sg13g2_and2_1 _7254_ (.A(net1169),
    .B(_3005_),
    .X(_3122_));
 sg13g2_nor2_1 _7255_ (.A(_3006_),
    .B(_3107_),
    .Y(_3123_));
 sg13g2_nand2_1 _7256_ (.Y(_3124_),
    .A(net1171),
    .B(_3084_));
 sg13g2_nand4_1 _7257_ (.B(_3006_),
    .C(_3042_),
    .A(net1171),
    .Y(_3125_),
    .D(_3086_));
 sg13g2_xnor2_1 _7258_ (.Y(_3126_),
    .A(_3086_),
    .B(_3123_));
 sg13g2_nand2_1 _7259_ (.Y(_3127_),
    .A(_3122_),
    .B(_3126_));
 sg13g2_xor2_1 _7260_ (.B(_3126_),
    .A(_3122_),
    .X(_3128_));
 sg13g2_nor2b_1 _7261_ (.A(_3121_),
    .B_N(_3128_),
    .Y(_3129_));
 sg13g2_xnor2_1 _7262_ (.Y(_3130_),
    .A(_3121_),
    .B(_3128_));
 sg13g2_o21ai_1 _7263_ (.B1(_3114_),
    .Y(_3131_),
    .A1(_3104_),
    .A2(_3115_));
 sg13g2_and2_1 _7264_ (.A(_3130_),
    .B(_3131_),
    .X(_3132_));
 sg13g2_xor2_1 _7265_ (.B(_3131_),
    .A(_3130_),
    .X(_3133_));
 sg13g2_o21ai_1 _7266_ (.B1(_3117_),
    .Y(_3134_),
    .A1(_3102_),
    .A2(_3118_));
 sg13g2_xnor2_1 _7267_ (.Y(_3135_),
    .A(_3133_),
    .B(_3134_));
 sg13g2_nand2_1 _7268_ (.Y(_3136_),
    .A(net1439),
    .B(net1015));
 sg13g2_a22oi_1 _7269_ (.Y(_0538_),
    .B1(_3136_),
    .B2(_2871_),
    .A2(_3135_),
    .A1(net1096));
 sg13g2_nand3_1 _7270_ (.B(_3043_),
    .C(_3084_),
    .A(net1171),
    .Y(_3137_));
 sg13g2_nand2_1 _7271_ (.Y(_3138_),
    .A(net1169),
    .B(_3042_));
 sg13g2_xnor2_1 _7272_ (.Y(_3139_),
    .A(_3137_),
    .B(_3138_));
 sg13g2_a21oi_1 _7273_ (.A1(_3125_),
    .A2(_3127_),
    .Y(_3140_),
    .B1(_3139_));
 sg13g2_nand3_1 _7274_ (.B(_3127_),
    .C(_3139_),
    .A(_3125_),
    .Y(_3141_));
 sg13g2_nor2b_1 _7275_ (.A(_3140_),
    .B_N(_3141_),
    .Y(_3142_));
 sg13g2_nand2_1 _7276_ (.Y(_3143_),
    .A(_3129_),
    .B(_3142_));
 sg13g2_xnor2_1 _7277_ (.Y(_3144_),
    .A(_3129_),
    .B(_3142_));
 sg13g2_a21oi_1 _7278_ (.A1(_3133_),
    .A2(_3134_),
    .Y(_3145_),
    .B1(_3132_));
 sg13g2_xnor2_1 _7279_ (.Y(_3146_),
    .A(_3144_),
    .B(_3145_));
 sg13g2_nand2_1 _7280_ (.Y(_3147_),
    .A(net1463),
    .B(net1015));
 sg13g2_a22oi_1 _7281_ (.Y(_0539_),
    .B1(_3147_),
    .B2(_2871_),
    .A2(_3146_),
    .A1(_1520_));
 sg13g2_o21ai_1 _7282_ (.B1(_3143_),
    .Y(_3148_),
    .A1(_3144_),
    .A2(_3145_));
 sg13g2_a21oi_1 _7283_ (.A1(_3043_),
    .A2(_3138_),
    .Y(_3149_),
    .B1(_3124_));
 sg13g2_nand2_1 _7284_ (.Y(_3150_),
    .A(net1169),
    .B(_3084_));
 sg13g2_xor2_1 _7285_ (.B(_3150_),
    .A(_3149_),
    .X(_3151_));
 sg13g2_xnor2_1 _7286_ (.Y(_3152_),
    .A(_3140_),
    .B(_3151_));
 sg13g2_xnor2_1 _7287_ (.Y(_3153_),
    .A(_3148_),
    .B(_3152_));
 sg13g2_nand3b_1 _7288_ (.B(net1015),
    .C(net1616),
    .Y(_3154_),
    .A_N(_1520_));
 sg13g2_o21ai_1 _7289_ (.B1(_3154_),
    .Y(_0540_),
    .A1(_2871_),
    .A2(_3153_));
 sg13g2_and2_1 _7290_ (.A(net1187),
    .B(_2897_),
    .X(_3155_));
 sg13g2_nand2_2 _7291_ (.Y(_3156_),
    .A(net1159),
    .B(_3155_));
 sg13g2_inv_1 _7292_ (.Y(_3157_),
    .A(_3156_));
 sg13g2_nor2_2 _7293_ (.A(_2874_),
    .B(_3155_),
    .Y(_3158_));
 sg13g2_nand2_1 _7294_ (.Y(_3159_),
    .A(net1236),
    .B(_3158_));
 sg13g2_o21ai_1 _7295_ (.B1(_3159_),
    .Y(_0541_),
    .A1(_2985_),
    .A2(_3156_));
 sg13g2_nand2_1 _7296_ (.Y(_3160_),
    .A(net1808),
    .B(net1082));
 sg13g2_a22oi_1 _7297_ (.Y(_3161_),
    .B1(_3160_),
    .B2(net1165),
    .A2(_3021_),
    .A1(_2897_));
 sg13g2_o21ai_1 _7298_ (.B1(net1159),
    .Y(_3162_),
    .A1(_3060_),
    .A2(_3161_));
 sg13g2_a21oi_1 _7299_ (.A1(_3060_),
    .A2(net1809),
    .Y(_0542_),
    .B1(_3162_));
 sg13g2_a22oi_1 _7300_ (.Y(_3163_),
    .B1(_3158_),
    .B2(net1491),
    .A2(_3157_),
    .A1(_3058_));
 sg13g2_inv_1 _7301_ (.Y(_0543_),
    .A(_3163_));
 sg13g2_nand2_1 _7302_ (.Y(_3164_),
    .A(net1320),
    .B(_3158_));
 sg13g2_o21ai_1 _7303_ (.B1(_3164_),
    .Y(_0544_),
    .A1(_3099_),
    .A2(_3156_));
 sg13g2_nand2_1 _7304_ (.Y(_3165_),
    .A(net1294),
    .B(_3158_));
 sg13g2_o21ai_1 _7305_ (.B1(_3165_),
    .Y(_0545_),
    .A1(_3119_),
    .A2(_3156_));
 sg13g2_nand2_1 _7306_ (.Y(_3166_),
    .A(net1411),
    .B(net1015));
 sg13g2_a22oi_1 _7307_ (.Y(_0546_),
    .B1(_3156_),
    .B2(_3166_),
    .A2(_3155_),
    .A1(_3135_));
 sg13g2_nand2_1 _7308_ (.Y(_3167_),
    .A(net1355),
    .B(net1016));
 sg13g2_a22oi_1 _7309_ (.Y(_0547_),
    .B1(_3156_),
    .B2(_3167_),
    .A2(_3155_),
    .A1(_3146_));
 sg13g2_nand2_1 _7310_ (.Y(_3168_),
    .A(net1358),
    .B(net1016));
 sg13g2_a22oi_1 _7311_ (.Y(_0548_),
    .B1(_3156_),
    .B2(_3168_),
    .A2(_3155_),
    .A1(_3153_));
 sg13g2_and2_1 _7312_ (.A(net1187),
    .B(net1013),
    .X(_3169_));
 sg13g2_o21ai_1 _7313_ (.B1(net1188),
    .Y(_3170_),
    .A1(net1655),
    .A2(net1012));
 sg13g2_a21oi_1 _7314_ (.A1(net1012),
    .A2(_2985_),
    .Y(_3171_),
    .B1(_3170_));
 sg13g2_a21oi_1 _7315_ (.A1(net1655),
    .A2(_1521_),
    .Y(_3172_),
    .B1(_3171_));
 sg13g2_nor2_1 _7316_ (.A(net1129),
    .B(net1656),
    .Y(_0549_));
 sg13g2_a22oi_1 _7317_ (.Y(_3173_),
    .B1(_3169_),
    .B2(net1159),
    .A2(net1015),
    .A1(net1778));
 sg13g2_a21oi_1 _7318_ (.A1(_3021_),
    .A2(_3169_),
    .Y(_0550_),
    .B1(_3173_));
 sg13g2_nand3_1 _7319_ (.B(_3058_),
    .C(_3169_),
    .A(net1161),
    .Y(_3174_));
 sg13g2_nand2_1 _7320_ (.Y(_3175_),
    .A(net1464),
    .B(net1016));
 sg13g2_o21ai_1 _7321_ (.B1(_3174_),
    .Y(_0551_),
    .A1(_3169_),
    .A2(_3175_));
 sg13g2_o21ai_1 _7322_ (.B1(net1187),
    .Y(_3176_),
    .A1(net1644),
    .A2(net1014));
 sg13g2_a21oi_1 _7323_ (.A1(net1014),
    .A2(_3099_),
    .Y(_3177_),
    .B1(_3176_));
 sg13g2_a21oi_1 _7324_ (.A1(net1644),
    .A2(_1521_),
    .Y(_3178_),
    .B1(_3177_));
 sg13g2_nor2_1 _7325_ (.A(net1131),
    .B(net1645),
    .Y(_0552_));
 sg13g2_o21ai_1 _7326_ (.B1(net1188),
    .Y(_3179_),
    .A1(net1657),
    .A2(net1012));
 sg13g2_a21oi_1 _7327_ (.A1(net1012),
    .A2(_3119_),
    .Y(_3180_),
    .B1(_3179_));
 sg13g2_a21oi_1 _7328_ (.A1(net1657),
    .A2(_1521_),
    .Y(_3181_),
    .B1(_3180_));
 sg13g2_nor2_1 _7329_ (.A(net1130),
    .B(net1658),
    .Y(_0553_));
 sg13g2_o21ai_1 _7330_ (.B1(net1188),
    .Y(_3182_),
    .A1(net1950),
    .A2(net1012));
 sg13g2_a21oi_1 _7331_ (.A1(net1012),
    .A2(_3135_),
    .Y(_3183_),
    .B1(_3182_));
 sg13g2_a21oi_1 _7332_ (.A1(net1950),
    .A2(_1521_),
    .Y(_3184_),
    .B1(_3183_));
 sg13g2_nor2_1 _7333_ (.A(net1129),
    .B(net1951),
    .Y(_0554_));
 sg13g2_o21ai_1 _7334_ (.B1(net1188),
    .Y(_3185_),
    .A1(net1758),
    .A2(net1012));
 sg13g2_a21oi_1 _7335_ (.A1(net1012),
    .A2(_3146_),
    .Y(_3186_),
    .B1(_3185_));
 sg13g2_a21oi_1 _7336_ (.A1(net1758),
    .A2(_1521_),
    .Y(_3187_),
    .B1(_3186_));
 sg13g2_nor2_1 _7337_ (.A(net1129),
    .B(net1759),
    .Y(_0555_));
 sg13g2_o21ai_1 _7338_ (.B1(net1188),
    .Y(_3188_),
    .A1(net1690),
    .A2(net1013));
 sg13g2_a21o_1 _7339_ (.A2(_3153_),
    .A1(net1013),
    .B1(_3188_),
    .X(_3189_));
 sg13g2_nand2_1 _7340_ (.Y(_3190_),
    .A(net1690),
    .B(_1521_));
 sg13g2_a21oi_1 _7341_ (.A1(_3189_),
    .A2(net1691),
    .Y(_0556_),
    .B1(net1130));
 sg13g2_and2_1 _7342_ (.A(net1188),
    .B(_2881_),
    .X(_3191_));
 sg13g2_nand2_2 _7343_ (.Y(_3192_),
    .A(net1188),
    .B(_2881_));
 sg13g2_o21ai_1 _7344_ (.B1(net1016),
    .Y(_3193_),
    .A1(net1847),
    .A2(net1011));
 sg13g2_a21oi_1 _7345_ (.A1(_2985_),
    .A2(net1011),
    .Y(_0557_),
    .B1(_3193_));
 sg13g2_o21ai_1 _7346_ (.B1(net1016),
    .Y(_3194_),
    .A1(net1870),
    .A2(_3191_));
 sg13g2_a21oi_1 _7347_ (.A1(_3021_),
    .A2(_3191_),
    .Y(_0558_),
    .B1(_3194_));
 sg13g2_nand2_1 _7348_ (.Y(_3195_),
    .A(_3058_),
    .B(net1011));
 sg13g2_nand3_1 _7349_ (.B(net1082),
    .C(_3192_),
    .A(net1578),
    .Y(_3196_));
 sg13g2_a21oi_1 _7350_ (.A1(_3195_),
    .A2(net1579),
    .Y(_0559_),
    .B1(net1130));
 sg13g2_and2_1 _7351_ (.A(net2327),
    .B(net1082),
    .X(_3197_));
 sg13g2_o21ai_1 _7352_ (.B1(net1161),
    .Y(_3198_),
    .A1(net1011),
    .A2(_3197_));
 sg13g2_a21oi_1 _7353_ (.A1(_3099_),
    .A2(net1011),
    .Y(_0560_),
    .B1(_3198_));
 sg13g2_o21ai_1 _7354_ (.B1(net1016),
    .Y(_3199_),
    .A1(net1931),
    .A2(net1011));
 sg13g2_a21oi_1 _7355_ (.A1(_3119_),
    .A2(_3191_),
    .Y(_0561_),
    .B1(_3199_));
 sg13g2_nand3_1 _7356_ (.B(_2872_),
    .C(_3192_),
    .A(net2284),
    .Y(_3200_));
 sg13g2_o21ai_1 _7357_ (.B1(_3200_),
    .Y(_3201_),
    .A1(_3135_),
    .A2(_3192_));
 sg13g2_and2_1 _7358_ (.A(net1159),
    .B(net2285),
    .X(_0562_));
 sg13g2_nand3_1 _7359_ (.B(_2872_),
    .C(_3192_),
    .A(net2311),
    .Y(_3202_));
 sg13g2_o21ai_1 _7360_ (.B1(_3202_),
    .Y(_3203_),
    .A1(_3146_),
    .A2(_3192_));
 sg13g2_and2_1 _7361_ (.A(net1159),
    .B(net2312),
    .X(_0563_));
 sg13g2_o21ai_1 _7362_ (.B1(net1016),
    .Y(_3204_),
    .A1(net1853),
    .A2(net1011));
 sg13g2_a21oi_1 _7363_ (.A1(_3153_),
    .A2(net1011),
    .Y(_0564_),
    .B1(_3204_));
 sg13g2_nor2_1 _7364_ (.A(net1165),
    .B(_2874_),
    .Y(_0565_));
 sg13g2_nor2_1 _7365_ (.A(_2874_),
    .B(_2899_),
    .Y(_0566_));
 sg13g2_and2_1 _7366_ (.A(net1157),
    .B(net2380),
    .X(_0567_));
 sg13g2_a22oi_1 _7367_ (.Y(_3205_),
    .B1(net1850),
    .B2(net1093),
    .A2(net1954),
    .A1(_0756_));
 sg13g2_nor2_1 _7368_ (.A(net1034),
    .B(net1955),
    .Y(_0568_));
 sg13g2_a22oi_1 _7369_ (.Y(_3206_),
    .B1(net1706),
    .B2(net1093),
    .A2(net1756),
    .A1(net1133));
 sg13g2_nor2_1 _7370_ (.A(net1034),
    .B(net1757),
    .Y(_0569_));
 sg13g2_a22oi_1 _7371_ (.Y(_3207_),
    .B1(net1769),
    .B2(net1093),
    .A2(net1969),
    .A1(net1133));
 sg13g2_nor2_1 _7372_ (.A(net1034),
    .B(net1970),
    .Y(_0570_));
 sg13g2_a22oi_1 _7373_ (.Y(_3208_),
    .B1(net1628),
    .B2(net1093),
    .A2(net1767),
    .A1(net1133));
 sg13g2_nor2_1 _7374_ (.A(net1034),
    .B(net1768),
    .Y(_0571_));
 sg13g2_a22oi_1 _7375_ (.Y(_3209_),
    .B1(net1796),
    .B2(net1093),
    .A2(net1851),
    .A1(net1133));
 sg13g2_nor2_1 _7376_ (.A(net1034),
    .B(net1852),
    .Y(_0572_));
 sg13g2_a22oi_1 _7377_ (.Y(_3210_),
    .B1(net1806),
    .B2(net1094),
    .A2(net1908),
    .A1(net1133));
 sg13g2_nor2_1 _7378_ (.A(net1034),
    .B(net1909),
    .Y(_0573_));
 sg13g2_a22oi_1 _7379_ (.Y(_3211_),
    .B1(net1734),
    .B2(net1093),
    .A2(net1864),
    .A1(net1133));
 sg13g2_nor2_1 _7380_ (.A(net1028),
    .B(net1865),
    .Y(_0574_));
 sg13g2_a22oi_1 _7381_ (.Y(_3212_),
    .B1(\led_controller.cpu.i_bus_data[7] ),
    .B2(net1093),
    .A2(net1133),
    .A1(net1742));
 sg13g2_nor2_1 _7382_ (.A(net1029),
    .B(net1743),
    .Y(_0575_));
 sg13g2_or3_1 _7383_ (.A(net1583),
    .B(_0903_),
    .C(_0917_),
    .X(_3213_));
 sg13g2_nand2_1 _7384_ (.Y(_3214_),
    .A(net1583),
    .B(_0917_));
 sg13g2_nor2_1 _7385_ (.A(\led_controller.register_address[6] ),
    .B(net2082),
    .Y(_3215_));
 sg13g2_and2_1 _7386_ (.A(net2305),
    .B(_3215_),
    .X(_3216_));
 sg13g2_nor2_2 _7387_ (.A(_0750_),
    .B(net1135),
    .Y(_3217_));
 sg13g2_nand2_1 _7388_ (.Y(_3218_),
    .A(net2128),
    .B(net1194));
 sg13g2_nor2_2 _7389_ (.A(net1136),
    .B(net1140),
    .Y(_3219_));
 sg13g2_and2_1 _7390_ (.A(\led_controller.register_address[1] ),
    .B(\led_controller.register_address[0] ),
    .X(_3220_));
 sg13g2_and2_1 _7391_ (.A(_3219_),
    .B(net1072),
    .X(_3221_));
 sg13g2_nand3_1 _7392_ (.B(_3217_),
    .C(_3221_),
    .A(_3216_),
    .Y(_3222_));
 sg13g2_nor2_2 _7393_ (.A(\led_controller.register_address[1] ),
    .B(\led_controller.register_address[0] ),
    .Y(_3223_));
 sg13g2_nor2b_1 _7394_ (.A(net1136),
    .B_N(net1138),
    .Y(_3224_));
 sg13g2_nand4_1 _7395_ (.B(_3217_),
    .C(net1068),
    .A(_3216_),
    .Y(_3225_),
    .D(_3224_));
 sg13g2_and2_1 _7396_ (.A(_3222_),
    .B(_3225_),
    .X(_3226_));
 sg13g2_nand2_1 _7397_ (.Y(_3227_),
    .A(net1144),
    .B(_3226_));
 sg13g2_a21oi_1 _7398_ (.A1(_3213_),
    .A2(_3214_),
    .Y(_0576_),
    .B1(_3227_));
 sg13g2_or2_1 _7399_ (.X(_3228_),
    .B(_3213_),
    .A(\led_controller.cpu_reset_counter[1] ));
 sg13g2_xor2_1 _7400_ (.B(_3213_),
    .A(net2321),
    .X(_3229_));
 sg13g2_a21oi_1 _7401_ (.A1(_3226_),
    .A2(_3229_),
    .Y(_0577_),
    .B1(net1105));
 sg13g2_xor2_1 _7402_ (.B(_3228_),
    .A(net2152),
    .X(_3230_));
 sg13g2_nor2_1 _7403_ (.A(_3227_),
    .B(net2153),
    .Y(_0578_));
 sg13g2_o21ai_1 _7404_ (.B1(net1568),
    .Y(_3231_),
    .A1(\led_controller.cpu_reset_counter[2] ),
    .A2(_3228_));
 sg13g2_a21oi_1 _7405_ (.A1(_3226_),
    .A2(net1569),
    .Y(_0579_),
    .B1(net1105));
 sg13g2_nor2_1 _7406_ (.A(net1134),
    .B(net1105),
    .Y(_0580_));
 sg13g2_a21oi_1 _7407_ (.A1(net2308),
    .A2(_3222_),
    .Y(_3232_),
    .B1(net1106));
 sg13g2_o21ai_1 _7408_ (.B1(_3232_),
    .Y(_0581_),
    .A1(_0747_),
    .A2(_3222_));
 sg13g2_nand2_1 _7409_ (.Y(_3233_),
    .A(net1134),
    .B(net1498));
 sg13g2_nor3_2 _7410_ (.A(\led_controller.register_address[6] ),
    .B(\led_controller.register_address[5] ),
    .C(\led_controller.register_address[4] ),
    .Y(_3234_));
 sg13g2_nand2b_2 _7411_ (.Y(_3235_),
    .B(_3215_),
    .A_N(\led_controller.register_address[4] ));
 sg13g2_nor2_2 _7412_ (.A(_3219_),
    .B(_3235_),
    .Y(_3236_));
 sg13g2_nand2b_2 _7413_ (.Y(_3237_),
    .B(_3234_),
    .A_N(_3219_));
 sg13g2_xor2_1 _7414_ (.B(\led_controller.register_address[4] ),
    .A(\led_controller.register_address[5] ),
    .X(_3238_));
 sg13g2_nor2b_2 _7415_ (.A(\led_controller.register_address[1] ),
    .B_N(\led_controller.register_address[0] ),
    .Y(_3239_));
 sg13g2_a22oi_1 _7416_ (.Y(_3240_),
    .B1(net1065),
    .B2(\led_controller.colors[80] ),
    .A2(net1070),
    .A1(\led_controller.colors[88] ));
 sg13g2_nor2_1 _7417_ (.A(_0752_),
    .B(\led_controller.register_address[0] ),
    .Y(_3241_));
 sg13g2_nand2b_2 _7418_ (.Y(_3242_),
    .B(\led_controller.register_address[1] ),
    .A_N(\led_controller.register_address[0] ));
 sg13g2_a22oi_1 _7419_ (.Y(_3243_),
    .B1(net1008),
    .B2(\led_controller.colors[72] ),
    .A2(net1074),
    .A1(\led_controller.colors[64] ));
 sg13g2_a21oi_1 _7420_ (.A1(_3240_),
    .A2(_3243_),
    .Y(_3244_),
    .B1(net1137));
 sg13g2_nand2_2 _7421_ (.Y(_3245_),
    .A(net1136),
    .B(net1140));
 sg13g2_a22oi_1 _7422_ (.Y(_3246_),
    .B1(net1066),
    .B2(\led_controller.colors[16] ),
    .A2(net1073),
    .A1(\led_controller.colors[0] ));
 sg13g2_a22oi_1 _7423_ (.Y(_3247_),
    .B1(net1007),
    .B2(\led_controller.colors[8] ),
    .A2(net1069),
    .A1(\led_controller.colors[24] ));
 sg13g2_a21oi_1 _7424_ (.A1(_3246_),
    .A2(_3247_),
    .Y(_3248_),
    .B1(net1061));
 sg13g2_a22oi_1 _7425_ (.Y(_3249_),
    .B1(net1007),
    .B2(\led_controller.colors[40] ),
    .A2(net1065),
    .A1(\led_controller.colors[48] ));
 sg13g2_a22oi_1 _7426_ (.Y(_3250_),
    .B1(net1069),
    .B2(\led_controller.colors[56] ),
    .A2(net1073),
    .A1(\led_controller.colors[32] ));
 sg13g2_a21oi_1 _7427_ (.A1(_3249_),
    .A2(_3250_),
    .Y(_3251_),
    .B1(net1141));
 sg13g2_nor3_2 _7428_ (.A(_3244_),
    .B(_3248_),
    .C(_3251_),
    .Y(_3252_));
 sg13g2_o21ai_1 _7429_ (.B1(net969),
    .Y(_3253_),
    .A1(_3238_),
    .A2(_3252_));
 sg13g2_nand3_1 _7430_ (.B(net1138),
    .C(net1072),
    .A(net1136),
    .Y(_3254_));
 sg13g2_and2_1 _7431_ (.A(_3234_),
    .B(net1064),
    .X(_3255_));
 sg13g2_and2_1 _7432_ (.A(_3219_),
    .B(net1004),
    .X(_3256_));
 sg13g2_nand3_1 _7433_ (.B(_3216_),
    .C(_3221_),
    .A(\led_controller.flash.i_addr_width_24 ),
    .Y(_3257_));
 sg13g2_nand2_1 _7434_ (.Y(_3258_),
    .A(_3216_),
    .B(_3219_));
 sg13g2_nor2_1 _7435_ (.A(net1062),
    .B(_3258_),
    .Y(_3259_));
 sg13g2_nor2_2 _7436_ (.A(net1010),
    .B(net1062),
    .Y(_3260_));
 sg13g2_nor2_1 _7437_ (.A(net969),
    .B(_3260_),
    .Y(_3261_));
 sg13g2_a21oi_1 _7438_ (.A1(\led_controller.register_address[1] ),
    .A2(_3234_),
    .Y(_3262_),
    .B1(net969));
 sg13g2_and3_2 _7439_ (.X(_3263_),
    .A(_3216_),
    .B(_3219_),
    .C(net1064));
 sg13g2_nor3_2 _7440_ (.A(\led_controller.register_address[1] ),
    .B(\led_controller.register_address[0] ),
    .C(_3258_),
    .Y(_3264_));
 sg13g2_a22oi_1 _7441_ (.Y(_3265_),
    .B1(_3263_),
    .B2(\led_controller.cpu.i_num_colors[0] ),
    .A2(_3256_),
    .A1(\led_controller.effect[0] ));
 sg13g2_a22oi_1 _7442_ (.Y(_3266_),
    .B1(net954),
    .B2(\led_controller.cpu.i_num_leds[0] ),
    .A2(net955),
    .A1(\led_controller.clock_divider[0] ));
 sg13g2_nand4_1 _7443_ (.B(_3262_),
    .C(_3265_),
    .A(_3257_),
    .Y(_3267_),
    .D(_3266_));
 sg13g2_nor2_2 _7444_ (.A(\led_controller.register_address[7] ),
    .B(net1134),
    .Y(_3268_));
 sg13g2_nand2_2 _7445_ (.Y(_3269_),
    .A(_0750_),
    .B(net1194));
 sg13g2_nand3_1 _7446_ (.B(_3267_),
    .C(_3268_),
    .A(_3253_),
    .Y(_3270_));
 sg13g2_a21oi_1 _7447_ (.A1(_3233_),
    .A2(_3270_),
    .Y(_0582_),
    .B1(net1106));
 sg13g2_and2_1 _7448_ (.A(\led_controller.effect[1] ),
    .B(_3256_),
    .X(_3271_));
 sg13g2_a21oi_1 _7449_ (.A1(\led_controller.cpu.i_num_colors[1] ),
    .A2(_3263_),
    .Y(_3272_),
    .B1(_3236_));
 sg13g2_a221oi_1 _7450_ (.B2(\led_controller.cpu.i_num_leds[1] ),
    .C1(_3271_),
    .B1(net954),
    .A1(\led_controller.clock_divider[1] ),
    .Y(_3273_),
    .A2(net955));
 sg13g2_a22oi_1 _7451_ (.Y(_3274_),
    .B1(net1008),
    .B2(\led_controller.colors[41] ),
    .A2(net1066),
    .A1(\led_controller.colors[49] ));
 sg13g2_a22oi_1 _7452_ (.Y(_3275_),
    .B1(net1070),
    .B2(\led_controller.colors[57] ),
    .A2(net1074),
    .A1(\led_controller.colors[33] ));
 sg13g2_a21oi_1 _7453_ (.A1(_3274_),
    .A2(_3275_),
    .Y(_3276_),
    .B1(net1141));
 sg13g2_a22oi_1 _7454_ (.Y(_3277_),
    .B1(net1066),
    .B2(\led_controller.colors[17] ),
    .A2(net1074),
    .A1(\led_controller.colors[1] ));
 sg13g2_a22oi_1 _7455_ (.Y(_3278_),
    .B1(net1008),
    .B2(\led_controller.colors[9] ),
    .A2(net1070),
    .A1(\led_controller.colors[25] ));
 sg13g2_a21oi_1 _7456_ (.A1(_3277_),
    .A2(_3278_),
    .Y(_3279_),
    .B1(net1061));
 sg13g2_a22oi_1 _7457_ (.Y(_3280_),
    .B1(net1070),
    .B2(\led_controller.colors[89] ),
    .A2(net1074),
    .A1(\led_controller.colors[65] ));
 sg13g2_a22oi_1 _7458_ (.Y(_3281_),
    .B1(net1008),
    .B2(\led_controller.colors[73] ),
    .A2(net1066),
    .A1(\led_controller.colors[81] ));
 sg13g2_a21oi_1 _7459_ (.A1(_3280_),
    .A2(_3281_),
    .Y(_3282_),
    .B1(net1137));
 sg13g2_nor4_1 _7460_ (.A(_3237_),
    .B(_3276_),
    .C(_3279_),
    .D(_3282_),
    .Y(_3283_));
 sg13g2_a21oi_1 _7461_ (.A1(_3272_),
    .A2(_3273_),
    .Y(_3284_),
    .B1(_3283_));
 sg13g2_a22oi_1 _7462_ (.Y(_3285_),
    .B1(_3268_),
    .B2(_3284_),
    .A2(net1744),
    .A1(net1134));
 sg13g2_nor2_1 _7463_ (.A(net1105),
    .B(net1745),
    .Y(_0583_));
 sg13g2_a22oi_1 _7464_ (.Y(_3286_),
    .B1(net1007),
    .B2(\led_controller.colors[42] ),
    .A2(net1069),
    .A1(\led_controller.colors[58] ));
 sg13g2_a22oi_1 _7465_ (.Y(_3287_),
    .B1(net1065),
    .B2(\led_controller.colors[50] ),
    .A2(net1073),
    .A1(\led_controller.colors[34] ));
 sg13g2_a21oi_1 _7466_ (.A1(_3286_),
    .A2(_3287_),
    .Y(_3288_),
    .B1(net1141));
 sg13g2_a22oi_1 _7467_ (.Y(_3289_),
    .B1(net1007),
    .B2(\led_controller.colors[10] ),
    .A2(net1065),
    .A1(\led_controller.colors[18] ));
 sg13g2_a22oi_1 _7468_ (.Y(_3290_),
    .B1(net1069),
    .B2(\led_controller.colors[26] ),
    .A2(net1073),
    .A1(\led_controller.colors[2] ));
 sg13g2_a21oi_1 _7469_ (.A1(_3289_),
    .A2(_3290_),
    .Y(_3291_),
    .B1(net1061));
 sg13g2_a22oi_1 _7470_ (.Y(_3292_),
    .B1(net1007),
    .B2(\led_controller.colors[74] ),
    .A2(net1073),
    .A1(\led_controller.colors[66] ));
 sg13g2_a22oi_1 _7471_ (.Y(_3293_),
    .B1(net1065),
    .B2(\led_controller.colors[82] ),
    .A2(net1069),
    .A1(\led_controller.colors[90] ));
 sg13g2_a21oi_1 _7472_ (.A1(_3292_),
    .A2(_3293_),
    .Y(_3294_),
    .B1(net1137));
 sg13g2_nor3_2 _7473_ (.A(_3288_),
    .B(_3291_),
    .C(_3294_),
    .Y(_3295_));
 sg13g2_o21ai_1 _7474_ (.B1(net969),
    .Y(_3296_),
    .A1(_3238_),
    .A2(_3295_));
 sg13g2_a221oi_1 _7475_ (.B2(\led_controller.cpu.i_num_leds[2] ),
    .C1(_3236_),
    .B1(_3264_),
    .A1(net1072),
    .Y(_3297_),
    .A2(_3234_));
 sg13g2_a22oi_1 _7476_ (.Y(_3298_),
    .B1(_3259_),
    .B2(\led_controller.clock_divider[2] ),
    .A2(_3256_),
    .A1(\led_controller.effect[2] ));
 sg13g2_a21oi_1 _7477_ (.A1(_3297_),
    .A2(_3298_),
    .Y(_3299_),
    .B1(_3269_));
 sg13g2_a22oi_1 _7478_ (.Y(_3300_),
    .B1(_3296_),
    .B2(_3299_),
    .A2(net2019),
    .A1(net1135));
 sg13g2_nor2_1 _7479_ (.A(net1106),
    .B(net2020),
    .Y(_0584_));
 sg13g2_a22oi_1 _7480_ (.Y(_3301_),
    .B1(net1008),
    .B2(\led_controller.colors[75] ),
    .A2(net1074),
    .A1(\led_controller.colors[67] ));
 sg13g2_a22oi_1 _7481_ (.Y(_3302_),
    .B1(net1066),
    .B2(\led_controller.colors[83] ),
    .A2(net1070),
    .A1(\led_controller.colors[91] ));
 sg13g2_a21oi_1 _7482_ (.A1(_3301_),
    .A2(_3302_),
    .Y(_3303_),
    .B1(\led_controller.register_address[3] ));
 sg13g2_a22oi_1 _7483_ (.Y(_3304_),
    .B1(net1008),
    .B2(\led_controller.colors[43] ),
    .A2(net1066),
    .A1(\led_controller.colors[51] ));
 sg13g2_a22oi_1 _7484_ (.Y(_3305_),
    .B1(net1070),
    .B2(\led_controller.colors[59] ),
    .A2(net1074),
    .A1(\led_controller.colors[35] ));
 sg13g2_a21oi_1 _7485_ (.A1(_3304_),
    .A2(_3305_),
    .Y(_3306_),
    .B1(net1141));
 sg13g2_a22oi_1 _7486_ (.Y(_3307_),
    .B1(net1008),
    .B2(\led_controller.colors[11] ),
    .A2(net1070),
    .A1(\led_controller.colors[27] ));
 sg13g2_a22oi_1 _7487_ (.Y(_3308_),
    .B1(net1066),
    .B2(\led_controller.colors[19] ),
    .A2(net1074),
    .A1(\led_controller.colors[3] ));
 sg13g2_a21oi_1 _7488_ (.A1(_3307_),
    .A2(_3308_),
    .Y(_3309_),
    .B1(_3245_));
 sg13g2_nor3_2 _7489_ (.A(_3303_),
    .B(_3306_),
    .C(_3309_),
    .Y(_3310_));
 sg13g2_o21ai_1 _7490_ (.B1(net969),
    .Y(_3311_),
    .A1(_3238_),
    .A2(_3310_));
 sg13g2_a221oi_1 _7491_ (.B2(\led_controller.clock_divider[3] ),
    .C1(_3236_),
    .B1(net955),
    .A1(_3234_),
    .Y(_3312_),
    .A2(net1009));
 sg13g2_a22oi_1 _7492_ (.Y(_3313_),
    .B1(net954),
    .B2(\led_controller.cpu.i_num_leds[3] ),
    .A2(_3256_),
    .A1(\led_controller.effect[3] ));
 sg13g2_a21oi_1 _7493_ (.A1(_3312_),
    .A2(_3313_),
    .Y(_3314_),
    .B1(_3269_));
 sg13g2_a22oi_1 _7494_ (.Y(_3315_),
    .B1(_3311_),
    .B2(_3314_),
    .A2(net2040),
    .A1(net1135));
 sg13g2_nor2_1 _7495_ (.A(net1106),
    .B(net2041),
    .Y(_0585_));
 sg13g2_a22oi_1 _7496_ (.Y(_3316_),
    .B1(net1007),
    .B2(\led_controller.colors[44] ),
    .A2(net1069),
    .A1(\led_controller.colors[60] ));
 sg13g2_a22oi_1 _7497_ (.Y(_3317_),
    .B1(net1065),
    .B2(\led_controller.colors[52] ),
    .A2(net1073),
    .A1(\led_controller.colors[36] ));
 sg13g2_a21oi_1 _7498_ (.A1(_3316_),
    .A2(_3317_),
    .Y(_3318_),
    .B1(net1141));
 sg13g2_a22oi_1 _7499_ (.Y(_3319_),
    .B1(net1007),
    .B2(\led_controller.colors[12] ),
    .A2(net1065),
    .A1(\led_controller.colors[20] ));
 sg13g2_a22oi_1 _7500_ (.Y(_3320_),
    .B1(net1069),
    .B2(\led_controller.colors[28] ),
    .A2(net1073),
    .A1(\led_controller.colors[4] ));
 sg13g2_a21oi_1 _7501_ (.A1(_3319_),
    .A2(_3320_),
    .Y(_3321_),
    .B1(net1061));
 sg13g2_a22oi_1 _7502_ (.Y(_3322_),
    .B1(net1007),
    .B2(\led_controller.colors[76] ),
    .A2(net1073),
    .A1(\led_controller.colors[68] ));
 sg13g2_a22oi_1 _7503_ (.Y(_3323_),
    .B1(net1065),
    .B2(\led_controller.colors[84] ),
    .A2(net1069),
    .A1(\led_controller.colors[92] ));
 sg13g2_a21oi_1 _7504_ (.A1(_3322_),
    .A2(_3323_),
    .Y(_3324_),
    .B1(net1137));
 sg13g2_nor3_1 _7505_ (.A(_3318_),
    .B(_3321_),
    .C(_3324_),
    .Y(_3325_));
 sg13g2_a22oi_1 _7506_ (.Y(_3326_),
    .B1(net954),
    .B2(\led_controller.cpu.i_num_leds[4] ),
    .A2(net955),
    .A1(\led_controller.clock_divider[4] ));
 sg13g2_o21ai_1 _7507_ (.B1(_3326_),
    .Y(_3327_),
    .A1(_3237_),
    .A2(_3325_));
 sg13g2_a22oi_1 _7508_ (.Y(_3328_),
    .B1(_3268_),
    .B2(_3327_),
    .A2(net1821),
    .A1(net1134));
 sg13g2_nor2_1 _7509_ (.A(net1105),
    .B(net1822),
    .Y(_0586_));
 sg13g2_a22oi_1 _7510_ (.Y(_3329_),
    .B1(net1006),
    .B2(\led_controller.colors[77] ),
    .A2(net1063),
    .A1(\led_controller.colors[85] ));
 sg13g2_a22oi_1 _7511_ (.Y(_3330_),
    .B1(net1067),
    .B2(\led_controller.colors[93] ),
    .A2(net1071),
    .A1(\led_controller.colors[69] ));
 sg13g2_a21oi_1 _7512_ (.A1(_3329_),
    .A2(_3330_),
    .Y(_3331_),
    .B1(net1137));
 sg13g2_a22oi_1 _7513_ (.Y(_3332_),
    .B1(net1006),
    .B2(\led_controller.colors[13] ),
    .A2(net1063),
    .A1(\led_controller.colors[21] ));
 sg13g2_a22oi_1 _7514_ (.Y(_3333_),
    .B1(net1067),
    .B2(\led_controller.colors[29] ),
    .A2(net1071),
    .A1(\led_controller.colors[5] ));
 sg13g2_a21oi_1 _7515_ (.A1(_3332_),
    .A2(_3333_),
    .Y(_3334_),
    .B1(net1061));
 sg13g2_a22oi_1 _7516_ (.Y(_3335_),
    .B1(net1006),
    .B2(\led_controller.colors[45] ),
    .A2(net1067),
    .A1(\led_controller.colors[61] ));
 sg13g2_a22oi_1 _7517_ (.Y(_3336_),
    .B1(net1063),
    .B2(\led_controller.colors[53] ),
    .A2(net1071),
    .A1(\led_controller.colors[37] ));
 sg13g2_a21oi_1 _7518_ (.A1(_3335_),
    .A2(_3336_),
    .Y(_3337_),
    .B1(net1140));
 sg13g2_nor3_1 _7519_ (.A(_3331_),
    .B(_3334_),
    .C(_3337_),
    .Y(_3338_));
 sg13g2_o21ai_1 _7520_ (.B1(net969),
    .Y(_3339_),
    .A1(_3238_),
    .A2(_3338_));
 sg13g2_a22oi_1 _7521_ (.Y(_3340_),
    .B1(net954),
    .B2(\led_controller.cpu.i_num_leds[5] ),
    .A2(net955),
    .A1(net1995));
 sg13g2_a21oi_1 _7522_ (.A1(_3262_),
    .A2(_3340_),
    .Y(_3341_),
    .B1(_3269_));
 sg13g2_a22oi_1 _7523_ (.Y(_3342_),
    .B1(_3339_),
    .B2(_3341_),
    .A2(net2075),
    .A1(net1135));
 sg13g2_nor2_1 _7524_ (.A(net1106),
    .B(net2076),
    .Y(_0587_));
 sg13g2_a22oi_1 _7525_ (.Y(_3343_),
    .B1(net1006),
    .B2(\led_controller.colors[46] ),
    .A2(net1067),
    .A1(\led_controller.colors[62] ));
 sg13g2_a22oi_1 _7526_ (.Y(_3344_),
    .B1(net1063),
    .B2(\led_controller.colors[54] ),
    .A2(net1071),
    .A1(\led_controller.colors[38] ));
 sg13g2_a21oi_1 _7527_ (.A1(_3343_),
    .A2(_3344_),
    .Y(_3345_),
    .B1(net1140));
 sg13g2_a22oi_1 _7528_ (.Y(_3346_),
    .B1(net1006),
    .B2(\led_controller.colors[14] ),
    .A2(net1063),
    .A1(\led_controller.colors[22] ));
 sg13g2_a22oi_1 _7529_ (.Y(_3347_),
    .B1(net1068),
    .B2(\led_controller.colors[30] ),
    .A2(net1071),
    .A1(\led_controller.colors[6] ));
 sg13g2_a21oi_1 _7530_ (.A1(_3346_),
    .A2(_3347_),
    .Y(_3348_),
    .B1(net1061));
 sg13g2_a22oi_1 _7531_ (.Y(_3349_),
    .B1(net1009),
    .B2(\led_controller.colors[78] ),
    .A2(net1064),
    .A1(\led_controller.colors[86] ));
 sg13g2_a22oi_1 _7532_ (.Y(_3350_),
    .B1(net1067),
    .B2(\led_controller.colors[94] ),
    .A2(net1075),
    .A1(\led_controller.colors[70] ));
 sg13g2_a21oi_1 _7533_ (.A1(_3349_),
    .A2(_3350_),
    .Y(_3351_),
    .B1(net1137));
 sg13g2_nor3_1 _7534_ (.A(_3345_),
    .B(_3348_),
    .C(_3351_),
    .Y(_3352_));
 sg13g2_o21ai_1 _7535_ (.B1(net969),
    .Y(_3353_),
    .A1(_3238_),
    .A2(_3352_));
 sg13g2_a22oi_1 _7536_ (.Y(_3354_),
    .B1(net954),
    .B2(\led_controller.cpu.i_num_leds[6] ),
    .A2(net955),
    .A1(\led_controller.clock_divider[6] ));
 sg13g2_a21oi_1 _7537_ (.A1(_3261_),
    .A2(_3354_),
    .Y(_3355_),
    .B1(_3269_));
 sg13g2_a22oi_1 _7538_ (.Y(_3356_),
    .B1(_3353_),
    .B2(_3355_),
    .A2(net2012),
    .A1(net1135));
 sg13g2_nor2_1 _7539_ (.A(net1109),
    .B(net2013),
    .Y(_0588_));
 sg13g2_a22oi_1 _7540_ (.Y(_3357_),
    .B1(net1063),
    .B2(\led_controller.colors[87] ),
    .A2(net1071),
    .A1(\led_controller.colors[71] ));
 sg13g2_a22oi_1 _7541_ (.Y(_3358_),
    .B1(net1006),
    .B2(\led_controller.colors[79] ),
    .A2(net1067),
    .A1(\led_controller.colors[95] ));
 sg13g2_a21oi_1 _7542_ (.A1(_3357_),
    .A2(_3358_),
    .Y(_3359_),
    .B1(net1137));
 sg13g2_a22oi_1 _7543_ (.Y(_3360_),
    .B1(net1006),
    .B2(\led_controller.colors[15] ),
    .A2(net1067),
    .A1(\led_controller.colors[31] ));
 sg13g2_a22oi_1 _7544_ (.Y(_3361_),
    .B1(net1063),
    .B2(\led_controller.colors[23] ),
    .A2(net1071),
    .A1(\led_controller.colors[7] ));
 sg13g2_a21oi_1 _7545_ (.A1(_3360_),
    .A2(_3361_),
    .Y(_3362_),
    .B1(net1061));
 sg13g2_a22oi_1 _7546_ (.Y(_3363_),
    .B1(net1006),
    .B2(\led_controller.colors[47] ),
    .A2(net1067),
    .A1(\led_controller.colors[63] ));
 sg13g2_a22oi_1 _7547_ (.Y(_3364_),
    .B1(net1063),
    .B2(\led_controller.colors[55] ),
    .A2(net1071),
    .A1(\led_controller.colors[39] ));
 sg13g2_a21oi_1 _7548_ (.A1(_3363_),
    .A2(_3364_),
    .Y(_3365_),
    .B1(net1140));
 sg13g2_nor3_2 _7549_ (.A(_3359_),
    .B(_3362_),
    .C(_3365_),
    .Y(_3366_));
 sg13g2_a22oi_1 _7550_ (.Y(_3367_),
    .B1(net954),
    .B2(\led_controller.cpu.i_num_leds[7] ),
    .A2(net955),
    .A1(\led_controller.clock_divider[7] ));
 sg13g2_o21ai_1 _7551_ (.B1(_3367_),
    .Y(_3368_),
    .A1(_3237_),
    .A2(_3366_));
 sg13g2_a22oi_1 _7552_ (.Y(_3369_),
    .B1(_3268_),
    .B2(_3368_),
    .A2(net1134),
    .A1(net1614));
 sg13g2_nor2_1 _7553_ (.A(net1105),
    .B(net1615),
    .Y(_0589_));
 sg13g2_o21ai_1 _7554_ (.B1(net1144),
    .Y(_3370_),
    .A1(net1994),
    .A2(net984));
 sg13g2_a21oi_1 _7555_ (.A1(_0747_),
    .A2(net983),
    .Y(_0590_),
    .B1(_3370_));
 sg13g2_o21ai_1 _7556_ (.B1(net1146),
    .Y(_3371_),
    .A1(net1952),
    .A2(net983));
 sg13g2_a21oi_1 _7557_ (.A1(_0746_),
    .A2(net983),
    .Y(_0591_),
    .B1(_3371_));
 sg13g2_o21ai_1 _7558_ (.B1(net1146),
    .Y(_3372_),
    .A1(net1785),
    .A2(net983));
 sg13g2_a21oi_1 _7559_ (.A1(_0745_),
    .A2(net983),
    .Y(_0592_),
    .B1(_3372_));
 sg13g2_o21ai_1 _7560_ (.B1(net1146),
    .Y(_3373_),
    .A1(net1797),
    .A2(net983));
 sg13g2_a21oi_1 _7561_ (.A1(_0744_),
    .A2(net983),
    .Y(_0593_),
    .B1(_3373_));
 sg13g2_o21ai_1 _7562_ (.B1(net1146),
    .Y(_3374_),
    .A1(net1906),
    .A2(net983));
 sg13g2_a21oi_1 _7563_ (.A1(_0743_),
    .A2(net984),
    .Y(_0594_),
    .B1(_3374_));
 sg13g2_o21ai_1 _7564_ (.B1(net1144),
    .Y(_3375_),
    .A1(net1695),
    .A2(net984));
 sg13g2_a21oi_1 _7565_ (.A1(_0742_),
    .A2(net984),
    .Y(_0595_),
    .B1(_3375_));
 sg13g2_o21ai_1 _7566_ (.B1(net1144),
    .Y(_3376_),
    .A1(net1633),
    .A2(net984));
 sg13g2_a21oi_1 _7567_ (.A1(_0741_),
    .A2(_0980_),
    .Y(_0596_),
    .B1(_3376_));
 sg13g2_o21ai_1 _7568_ (.B1(net1145),
    .Y(_3377_),
    .A1(net1916),
    .A2(net984));
 sg13g2_a21oi_1 _7569_ (.A1(_0740_),
    .A2(net984),
    .Y(_0597_),
    .B1(_3377_));
 sg13g2_nor2_2 _7570_ (.A(net1194),
    .B(_0975_),
    .Y(_3378_));
 sg13g2_a21oi_2 _7571_ (.B1(net1194),
    .Y(_3379_),
    .A2(_0973_),
    .A1(net2317));
 sg13g2_nor2_1 _7572_ (.A(net2319),
    .B(net1135),
    .Y(_3380_));
 sg13g2_a221oi_1 _7573_ (.B2(net2319),
    .C1(_3380_),
    .B1(_3379_),
    .A1(net1994),
    .Y(_3381_),
    .A2(_3378_));
 sg13g2_nor2_1 _7574_ (.A(net1104),
    .B(net2320),
    .Y(_0598_));
 sg13g2_o21ai_1 _7575_ (.B1(net1194),
    .Y(_3382_),
    .A1(net1072),
    .A2(net1068));
 sg13g2_nand2_1 _7576_ (.Y(_3383_),
    .A(net1144),
    .B(_3382_));
 sg13g2_a221oi_1 _7577_ (.B2(_0752_),
    .C1(_3383_),
    .B1(_3379_),
    .A1(_0754_),
    .Y(_0599_),
    .A2(_3378_));
 sg13g2_nand2_1 _7578_ (.Y(_3384_),
    .A(net1785),
    .B(_3378_));
 sg13g2_xor2_1 _7579_ (.B(net1072),
    .A(net1138),
    .X(_3385_));
 sg13g2_inv_2 _7580_ (.Y(_3386_),
    .A(_3385_));
 sg13g2_a22oi_1 _7581_ (.Y(_3387_),
    .B1(_3385_),
    .B2(\led_controller.spi_state[2] ),
    .A2(_3379_),
    .A1(net1138));
 sg13g2_a21oi_1 _7582_ (.A1(net1786),
    .A2(_3387_),
    .Y(_0600_),
    .B1(net1108));
 sg13g2_a21o_1 _7583_ (.A2(net1072),
    .A1(net1138),
    .B1(net1136),
    .X(_3388_));
 sg13g2_and2_1 _7584_ (.A(_3254_),
    .B(_3388_),
    .X(_3389_));
 sg13g2_inv_1 _7585_ (.Y(_3390_),
    .A(_3389_));
 sg13g2_nand2_1 _7586_ (.Y(_3391_),
    .A(net1797),
    .B(_3378_));
 sg13g2_a22oi_1 _7587_ (.Y(_3392_),
    .B1(_3389_),
    .B2(\led_controller.spi_state[2] ),
    .A2(_3379_),
    .A1(net1136));
 sg13g2_a21oi_1 _7588_ (.A1(net1798),
    .A2(_3392_),
    .Y(_0601_),
    .B1(net1108));
 sg13g2_a22oi_1 _7589_ (.Y(_3393_),
    .B1(_3379_),
    .B2(net2305),
    .A2(_3378_),
    .A1(net1906));
 sg13g2_nand4_1 _7590_ (.B(net1136),
    .C(net1138),
    .A(\led_controller.register_address[4] ),
    .Y(_3394_),
    .D(net1072));
 sg13g2_xor2_1 _7591_ (.B(_3254_),
    .A(net2305),
    .X(_3395_));
 sg13g2_or2_1 _7592_ (.X(_3396_),
    .B(_3395_),
    .A(net1135));
 sg13g2_a21oi_1 _7593_ (.A1(net2306),
    .A2(_3396_),
    .Y(_0602_),
    .B1(net1109));
 sg13g2_nor2_1 _7594_ (.A(_0751_),
    .B(_3394_),
    .Y(_3397_));
 sg13g2_nand2_1 _7595_ (.Y(_3398_),
    .A(net1194),
    .B(_3397_));
 sg13g2_nand2_1 _7596_ (.Y(_3399_),
    .A(net2082),
    .B(_0975_));
 sg13g2_a22oi_1 _7597_ (.Y(_3400_),
    .B1(net2083),
    .B2(net1134),
    .A2(_3394_),
    .A1(_0751_));
 sg13g2_a22oi_1 _7598_ (.Y(_3401_),
    .B1(_3398_),
    .B2(net2084),
    .A2(_3378_),
    .A1(net1695));
 sg13g2_nor2_1 _7599_ (.A(net1104),
    .B(net2085),
    .Y(_0603_));
 sg13g2_or2_1 _7600_ (.X(_3402_),
    .B(_3398_),
    .A(\led_controller.register_address[6] ));
 sg13g2_o21ai_1 _7601_ (.B1(_3398_),
    .Y(_3403_),
    .A1(\led_controller.register_address[6] ),
    .A2(_3378_));
 sg13g2_a221oi_1 _7602_ (.B2(_3403_),
    .C1(net1104),
    .B1(_3402_),
    .A1(_0753_),
    .Y(_0604_),
    .A2(_3378_));
 sg13g2_nand2_1 _7603_ (.Y(_3404_),
    .A(\led_controller.register_address[6] ),
    .B(_3397_));
 sg13g2_o21ai_1 _7604_ (.B1(net1134),
    .Y(_3405_),
    .A1(net1916),
    .A2(_0975_));
 sg13g2_mux2_1 _7605_ (.A0(_3269_),
    .A1(_3218_),
    .S(_3404_),
    .X(_3406_));
 sg13g2_a221oi_1 _7606_ (.B2(_3406_),
    .C1(net1104),
    .B1(_3405_),
    .A1(_0750_),
    .Y(_0605_),
    .A2(_3379_));
 sg13g2_nand2_2 _7607_ (.Y(_3407_),
    .A(_3217_),
    .B(_3263_));
 sg13g2_a21oi_1 _7608_ (.A1(net2345),
    .A2(_3407_),
    .Y(_3408_),
    .B1(net1106));
 sg13g2_o21ai_1 _7609_ (.B1(_3408_),
    .Y(_0606_),
    .A1(_0747_),
    .A2(_3407_));
 sg13g2_a21oi_1 _7610_ (.A1(net2264),
    .A2(_3407_),
    .Y(_3409_),
    .B1(net1107));
 sg13g2_o21ai_1 _7611_ (.B1(_3409_),
    .Y(_0607_),
    .A1(_0746_),
    .A2(_3407_));
 sg13g2_nand2_2 _7612_ (.Y(_3410_),
    .A(_3217_),
    .B(net969));
 sg13g2_nor2_2 _7613_ (.A(_3395_),
    .B(_3410_),
    .Y(_3411_));
 sg13g2_o21ai_1 _7614_ (.B1(net1155),
    .Y(_3412_),
    .A1(net2262),
    .A2(net890));
 sg13g2_a21oi_1 _7615_ (.A1(_0747_),
    .A2(net890),
    .Y(_0608_),
    .B1(_3412_));
 sg13g2_o21ai_1 _7616_ (.B1(net1146),
    .Y(_3413_),
    .A1(\led_controller.colors[1] ),
    .A2(net890));
 sg13g2_a21oi_1 _7617_ (.A1(_0746_),
    .A2(net890),
    .Y(_0609_),
    .B1(_3413_));
 sg13g2_o21ai_1 _7618_ (.B1(net1155),
    .Y(_3414_),
    .A1(net2122),
    .A2(net890));
 sg13g2_a21oi_1 _7619_ (.A1(_0745_),
    .A2(_3411_),
    .Y(_0610_),
    .B1(_3414_));
 sg13g2_o21ai_1 _7620_ (.B1(net1146),
    .Y(_3415_),
    .A1(\led_controller.colors[3] ),
    .A2(net890));
 sg13g2_a21oi_1 _7621_ (.A1(_0744_),
    .A2(net890),
    .Y(_0611_),
    .B1(_3415_));
 sg13g2_o21ai_1 _7622_ (.B1(net1156),
    .Y(_3416_),
    .A1(net2090),
    .A2(net890));
 sg13g2_a21oi_1 _7623_ (.A1(_0743_),
    .A2(net891),
    .Y(_0612_),
    .B1(_3416_));
 sg13g2_o21ai_1 _7624_ (.B1(net1155),
    .Y(_3417_),
    .A1(\led_controller.colors[5] ),
    .A2(net891));
 sg13g2_a21oi_1 _7625_ (.A1(_0742_),
    .A2(net891),
    .Y(_0613_),
    .B1(_3417_));
 sg13g2_o21ai_1 _7626_ (.B1(net1155),
    .Y(_3418_),
    .A1(\led_controller.colors[6] ),
    .A2(net891));
 sg13g2_a21oi_1 _7627_ (.A1(_0741_),
    .A2(net891),
    .Y(_0614_),
    .B1(_3418_));
 sg13g2_o21ai_1 _7628_ (.B1(net1151),
    .Y(_3419_),
    .A1(net2088),
    .A2(net891));
 sg13g2_a21oi_1 _7629_ (.A1(_0740_),
    .A2(net891),
    .Y(_0615_),
    .B1(_3419_));
 sg13g2_nor2_1 _7630_ (.A(_3390_),
    .B(_3410_),
    .Y(_3420_));
 sg13g2_nand3_1 _7631_ (.B(_3260_),
    .C(_3420_),
    .A(net1138),
    .Y(_3421_));
 sg13g2_nor3_2 _7632_ (.A(_0747_),
    .B(net1010),
    .C(net1062),
    .Y(_3422_));
 sg13g2_nor2_2 _7633_ (.A(_3386_),
    .B(_3410_),
    .Y(_3423_));
 sg13g2_nor3_1 _7634_ (.A(_3386_),
    .B(_3390_),
    .C(_3410_),
    .Y(_3424_));
 sg13g2_a22oi_1 _7635_ (.Y(_3425_),
    .B1(_3422_),
    .B2(net888),
    .A2(_3421_),
    .A1(net2302));
 sg13g2_nand2_1 _7636_ (.Y(_0616_),
    .A(net1160),
    .B(net2303));
 sg13g2_nor3_2 _7637_ (.A(_0746_),
    .B(net1010),
    .C(_3242_),
    .Y(_3426_));
 sg13g2_a22oi_1 _7638_ (.Y(_3427_),
    .B1(net887),
    .B2(_3426_),
    .A2(_3421_),
    .A1(net2297));
 sg13g2_nand2_1 _7639_ (.Y(_0617_),
    .A(net1158),
    .B(net2298));
 sg13g2_nor3_1 _7640_ (.A(_0745_),
    .B(net1010),
    .C(_3242_),
    .Y(_3428_));
 sg13g2_a22oi_1 _7641_ (.Y(_3429_),
    .B1(net887),
    .B2(_3428_),
    .A2(_3421_),
    .A1(net2279));
 sg13g2_nand2_1 _7642_ (.Y(_0618_),
    .A(net1155),
    .B(net2280));
 sg13g2_nor3_1 _7643_ (.A(_0744_),
    .B(net1010),
    .C(_3242_),
    .Y(_3430_));
 sg13g2_a22oi_1 _7644_ (.Y(_3431_),
    .B1(net887),
    .B2(_3430_),
    .A2(_3421_),
    .A1(net2254));
 sg13g2_nand2_1 _7645_ (.Y(_0619_),
    .A(net1146),
    .B(net2255));
 sg13g2_nor3_1 _7646_ (.A(_0743_),
    .B(net1010),
    .C(net1062),
    .Y(_3432_));
 sg13g2_a22oi_1 _7647_ (.Y(_3433_),
    .B1(net888),
    .B2(_3432_),
    .A2(_3421_),
    .A1(net2199));
 sg13g2_nand2_1 _7648_ (.Y(_0620_),
    .A(net1155),
    .B(_3433_));
 sg13g2_nor3_1 _7649_ (.A(_0742_),
    .B(net1010),
    .C(net1062),
    .Y(_3434_));
 sg13g2_a22oi_1 _7650_ (.Y(_3435_),
    .B1(net886),
    .B2(_3434_),
    .A2(_3421_),
    .A1(net2250));
 sg13g2_nand2_1 _7651_ (.Y(_0621_),
    .A(net1151),
    .B(_3435_));
 sg13g2_nor3_2 _7652_ (.A(_0741_),
    .B(_3235_),
    .C(net1062),
    .Y(_3436_));
 sg13g2_a22oi_1 _7653_ (.Y(_3437_),
    .B1(net886),
    .B2(_3436_),
    .A2(_3421_),
    .A1(net2180));
 sg13g2_nand2_1 _7654_ (.Y(_0622_),
    .A(net1155),
    .B(net2181));
 sg13g2_nor3_1 _7655_ (.A(_0740_),
    .B(net1010),
    .C(net1062),
    .Y(_3438_));
 sg13g2_a22oi_1 _7656_ (.Y(_3439_),
    .B1(net886),
    .B2(_3438_),
    .A2(_3421_),
    .A1(net2271));
 sg13g2_nand2_1 _7657_ (.Y(_0623_),
    .A(net1151),
    .B(_3439_));
 sg13g2_and2_1 _7658_ (.A(\led_controller.register_data[0] ),
    .B(net1004),
    .X(_3440_));
 sg13g2_nand3_1 _7659_ (.B(net1004),
    .C(_3420_),
    .A(net1139),
    .Y(_3441_));
 sg13g2_a22oi_1 _7660_ (.Y(_3442_),
    .B1(_3441_),
    .B2(net1967),
    .A2(_3440_),
    .A1(net888));
 sg13g2_nor2_1 _7661_ (.A(net1127),
    .B(net1968),
    .Y(_0624_));
 sg13g2_and2_1 _7662_ (.A(net2124),
    .B(net1005),
    .X(_3443_));
 sg13g2_a22oi_1 _7663_ (.Y(_3444_),
    .B1(_3443_),
    .B2(net887),
    .A2(_3441_),
    .A1(net2016));
 sg13g2_nor2_1 _7664_ (.A(net1119),
    .B(net2017),
    .Y(_0625_));
 sg13g2_and2_1 _7665_ (.A(net2091),
    .B(net1005),
    .X(_3445_));
 sg13g2_a22oi_1 _7666_ (.Y(_3446_),
    .B1(_3445_),
    .B2(net888),
    .A2(_3441_),
    .A1(net2269));
 sg13g2_nor2_1 _7667_ (.A(net1128),
    .B(_3446_),
    .Y(_0626_));
 sg13g2_and2_1 _7668_ (.A(net2000),
    .B(net1005),
    .X(_3447_));
 sg13g2_a22oi_1 _7669_ (.Y(_3448_),
    .B1(_3447_),
    .B2(net887),
    .A2(_3441_),
    .A1(net2150));
 sg13g2_nor2_1 _7670_ (.A(net1119),
    .B(_3448_),
    .Y(_0627_));
 sg13g2_and2_1 _7671_ (.A(net2047),
    .B(net1005),
    .X(_3449_));
 sg13g2_a22oi_1 _7672_ (.Y(_3450_),
    .B1(_3449_),
    .B2(net888),
    .A2(_3441_),
    .A1(net2021));
 sg13g2_nor2_1 _7673_ (.A(net1124),
    .B(net2022),
    .Y(_0628_));
 sg13g2_and2_1 _7674_ (.A(net1948),
    .B(net1004),
    .X(_3451_));
 sg13g2_a22oi_1 _7675_ (.Y(_3452_),
    .B1(_3451_),
    .B2(net886),
    .A2(_3441_),
    .A1(net2261));
 sg13g2_nor2_1 _7676_ (.A(net1110),
    .B(_3452_),
    .Y(_0629_));
 sg13g2_and2_1 _7677_ (.A(\led_controller.register_data[6] ),
    .B(net1004),
    .X(_3453_));
 sg13g2_a22oi_1 _7678_ (.Y(_3454_),
    .B1(_3453_),
    .B2(net886),
    .A2(_3441_),
    .A1(net2120));
 sg13g2_nor2_1 _7679_ (.A(net1112),
    .B(net2121),
    .Y(_0630_));
 sg13g2_and2_1 _7680_ (.A(net2042),
    .B(net1004),
    .X(_3455_));
 sg13g2_a22oi_1 _7681_ (.Y(_3456_),
    .B1(_3455_),
    .B2(net886),
    .A2(_3441_),
    .A1(net2178));
 sg13g2_nor2_1 _7682_ (.A(net1111),
    .B(_3456_),
    .Y(_0631_));
 sg13g2_and2_1 _7683_ (.A(net1068),
    .B(_3234_),
    .X(_3457_));
 sg13g2_and2_1 _7684_ (.A(\led_controller.register_data[0] ),
    .B(net1003),
    .X(_3458_));
 sg13g2_nand3_1 _7685_ (.B(_3420_),
    .C(net1003),
    .A(net1139),
    .Y(_3459_));
 sg13g2_a22oi_1 _7686_ (.Y(_3460_),
    .B1(_3459_),
    .B2(net1910),
    .A2(_3458_),
    .A1(net888));
 sg13g2_nor2_1 _7687_ (.A(net1123),
    .B(net1911),
    .Y(_0632_));
 sg13g2_and2_1 _7688_ (.A(net2124),
    .B(_3457_),
    .X(_3461_));
 sg13g2_a22oi_1 _7689_ (.Y(_3462_),
    .B1(_3461_),
    .B2(net887),
    .A2(_3459_),
    .A1(net2299));
 sg13g2_nor2_1 _7690_ (.A(net1122),
    .B(_3462_),
    .Y(_0633_));
 sg13g2_and2_1 _7691_ (.A(net2091),
    .B(_3457_),
    .X(_3463_));
 sg13g2_a22oi_1 _7692_ (.Y(_3464_),
    .B1(_3463_),
    .B2(net887),
    .A2(_3459_),
    .A1(net2057));
 sg13g2_nor2_1 _7693_ (.A(net1119),
    .B(net2058),
    .Y(_0634_));
 sg13g2_and2_1 _7694_ (.A(net2000),
    .B(_3457_),
    .X(_3465_));
 sg13g2_a22oi_1 _7695_ (.Y(_3466_),
    .B1(_3465_),
    .B2(net887),
    .A2(_3459_),
    .A1(net2098));
 sg13g2_nor2_1 _7696_ (.A(net1119),
    .B(_3466_),
    .Y(_0635_));
 sg13g2_and2_1 _7697_ (.A(net2047),
    .B(net1003),
    .X(_3467_));
 sg13g2_a22oi_1 _7698_ (.Y(_3468_),
    .B1(_3467_),
    .B2(net888),
    .A2(_3459_),
    .A1(net1998));
 sg13g2_nor2_1 _7699_ (.A(net1124),
    .B(net1999),
    .Y(_0636_));
 sg13g2_and2_1 _7700_ (.A(net1948),
    .B(net1003),
    .X(_3469_));
 sg13g2_a22oi_1 _7701_ (.Y(_3470_),
    .B1(_3469_),
    .B2(net886),
    .A2(_3459_),
    .A1(net2006));
 sg13g2_nor2_1 _7702_ (.A(net1112),
    .B(_3470_),
    .Y(_0637_));
 sg13g2_and2_1 _7703_ (.A(net2140),
    .B(net1003),
    .X(_3471_));
 sg13g2_a22oi_1 _7704_ (.Y(_3472_),
    .B1(_3471_),
    .B2(net889),
    .A2(_3459_),
    .A1(net2206));
 sg13g2_nor2_1 _7705_ (.A(net1112),
    .B(_3472_),
    .Y(_0638_));
 sg13g2_and2_1 _7706_ (.A(net2042),
    .B(net1003),
    .X(_3473_));
 sg13g2_a22oi_1 _7707_ (.Y(_3474_),
    .B1(_3473_),
    .B2(net886),
    .A2(_3459_),
    .A1(net2135));
 sg13g2_nor2_1 _7708_ (.A(net1114),
    .B(_3474_),
    .Y(_0639_));
 sg13g2_and3_2 _7709_ (.X(_3475_),
    .A(net1072),
    .B(_3234_),
    .C(net1061));
 sg13g2_nand2_2 _7710_ (.Y(_3476_),
    .A(net889),
    .B(net1002));
 sg13g2_and2_1 _7711_ (.A(\led_controller.register_data[0] ),
    .B(net1002),
    .X(_3477_));
 sg13g2_a22oi_1 _7712_ (.Y(_3478_),
    .B1(_3477_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net2068));
 sg13g2_nor2_1 _7713_ (.A(net1123),
    .B(net2069),
    .Y(_0640_));
 sg13g2_and2_1 _7714_ (.A(\led_controller.register_data[1] ),
    .B(net1002),
    .X(_3479_));
 sg13g2_a22oi_1 _7715_ (.Y(_3480_),
    .B1(_3479_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net2030));
 sg13g2_nor2_1 _7716_ (.A(net1118),
    .B(net2031),
    .Y(_0641_));
 sg13g2_and2_1 _7717_ (.A(\led_controller.register_data[2] ),
    .B(net1002),
    .X(_3481_));
 sg13g2_a22oi_1 _7718_ (.Y(_3482_),
    .B1(_3481_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net1985));
 sg13g2_nor2_1 _7719_ (.A(net1118),
    .B(net1986),
    .Y(_0642_));
 sg13g2_and2_1 _7720_ (.A(net2000),
    .B(_3475_),
    .X(_3483_));
 sg13g2_a22oi_1 _7721_ (.Y(_3484_),
    .B1(_3483_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net2061));
 sg13g2_nor2_1 _7722_ (.A(net1118),
    .B(_3484_),
    .Y(_0643_));
 sg13g2_and2_1 _7723_ (.A(\led_controller.register_data[4] ),
    .B(_3475_),
    .X(_3485_));
 sg13g2_a22oi_1 _7724_ (.Y(_3486_),
    .B1(_3485_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net1989));
 sg13g2_nor2_1 _7725_ (.A(net1124),
    .B(net1990),
    .Y(_0644_));
 sg13g2_and2_1 _7726_ (.A(net1948),
    .B(net1002),
    .X(_3487_));
 sg13g2_a22oi_1 _7727_ (.Y(_3488_),
    .B1(_3487_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net2062));
 sg13g2_nor2_1 _7728_ (.A(net1108),
    .B(_3488_),
    .Y(_0645_));
 sg13g2_and2_1 _7729_ (.A(\led_controller.register_data[6] ),
    .B(net1002),
    .X(_3489_));
 sg13g2_a22oi_1 _7730_ (.Y(_3490_),
    .B1(_3489_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net2036));
 sg13g2_nor2_1 _7731_ (.A(net1113),
    .B(net2037),
    .Y(_0646_));
 sg13g2_and2_1 _7732_ (.A(\led_controller.register_data[7] ),
    .B(net1002),
    .X(_3491_));
 sg13g2_a22oi_1 _7733_ (.Y(_3492_),
    .B1(_3491_),
    .B2(_3423_),
    .A2(_3476_),
    .A1(net1996));
 sg13g2_nor2_1 _7734_ (.A(net1112),
    .B(net1997),
    .Y(_0647_));
 sg13g2_nor2_1 _7735_ (.A(_3385_),
    .B(_3410_),
    .Y(_3493_));
 sg13g2_nand3_1 _7736_ (.B(_3389_),
    .C(net881),
    .A(_3260_),
    .Y(_3494_));
 sg13g2_a22oi_1 _7737_ (.Y(_3495_),
    .B1(_3494_),
    .B2(net1746),
    .A2(net884),
    .A1(_3422_));
 sg13g2_nor2_1 _7738_ (.A(net1123),
    .B(net1747),
    .Y(_0648_));
 sg13g2_a22oi_1 _7739_ (.Y(_3496_),
    .B1(_3494_),
    .B2(net1858),
    .A2(net883),
    .A1(_3426_));
 sg13g2_nor2_1 _7740_ (.A(net1119),
    .B(net1859),
    .Y(_0649_));
 sg13g2_a22oi_1 _7741_ (.Y(_3497_),
    .B1(_3494_),
    .B2(net1841),
    .A2(net882),
    .A1(_3428_));
 sg13g2_nor2_1 _7742_ (.A(net1108),
    .B(net1842),
    .Y(_0650_));
 sg13g2_a22oi_1 _7743_ (.Y(_3498_),
    .B1(_3494_),
    .B2(net1830),
    .A2(net882),
    .A1(_3430_));
 sg13g2_nor2_1 _7744_ (.A(net1118),
    .B(net1831),
    .Y(_0651_));
 sg13g2_a22oi_1 _7745_ (.Y(_3499_),
    .B1(_3494_),
    .B2(net1764),
    .A2(net885),
    .A1(_3432_));
 sg13g2_nor2_1 _7746_ (.A(net1124),
    .B(net1765),
    .Y(_0652_));
 sg13g2_a22oi_1 _7747_ (.Y(_3500_),
    .B1(_3494_),
    .B2(net2018),
    .A2(net880),
    .A1(_3434_));
 sg13g2_nor2_1 _7748_ (.A(net1110),
    .B(_3500_),
    .Y(_0653_));
 sg13g2_a22oi_1 _7749_ (.Y(_3501_),
    .B1(_3494_),
    .B2(net1679),
    .A2(net881),
    .A1(_3436_));
 sg13g2_nor2_1 _7750_ (.A(net1113),
    .B(net1680),
    .Y(_0654_));
 sg13g2_a22oi_1 _7751_ (.Y(_3502_),
    .B1(_3494_),
    .B2(net1862),
    .A2(net880),
    .A1(_3438_));
 sg13g2_nor2_1 _7752_ (.A(net1111),
    .B(net1863),
    .Y(_0655_));
 sg13g2_nand3_1 _7753_ (.B(_3389_),
    .C(net881),
    .A(net1004),
    .Y(_3503_));
 sg13g2_a22oi_1 _7754_ (.Y(_3504_),
    .B1(_3503_),
    .B2(net1819),
    .A2(net884),
    .A1(_3440_));
 sg13g2_nor2_1 _7755_ (.A(net1123),
    .B(net1820),
    .Y(_0656_));
 sg13g2_a22oi_1 _7756_ (.Y(_3505_),
    .B1(_3503_),
    .B2(net1762),
    .A2(net882),
    .A1(_3443_));
 sg13g2_nor2_1 _7757_ (.A(net1119),
    .B(net1763),
    .Y(_0657_));
 sg13g2_a22oi_1 _7758_ (.Y(_3506_),
    .B1(_3503_),
    .B2(net2233),
    .A2(net883),
    .A1(_3445_));
 sg13g2_nor2_1 _7759_ (.A(net1121),
    .B(_3506_),
    .Y(_0658_));
 sg13g2_a22oi_1 _7760_ (.Y(_3507_),
    .B1(_3503_),
    .B2(net2179),
    .A2(net882),
    .A1(_3447_));
 sg13g2_nor2_1 _7761_ (.A(net1122),
    .B(_3507_),
    .Y(_0659_));
 sg13g2_a22oi_1 _7762_ (.Y(_3508_),
    .B1(_3503_),
    .B2(net1752),
    .A2(net884),
    .A1(_3449_));
 sg13g2_nor2_1 _7763_ (.A(net1124),
    .B(net1753),
    .Y(_0660_));
 sg13g2_a22oi_1 _7764_ (.Y(_3509_),
    .B1(_3503_),
    .B2(net2046),
    .A2(net880),
    .A1(_3451_));
 sg13g2_nor2_1 _7765_ (.A(net1110),
    .B(_3509_),
    .Y(_0661_));
 sg13g2_a22oi_1 _7766_ (.Y(_3510_),
    .B1(_3503_),
    .B2(net1983),
    .A2(net881),
    .A1(_3453_));
 sg13g2_nor2_1 _7767_ (.A(net1113),
    .B(net1984),
    .Y(_0662_));
 sg13g2_a22oi_1 _7768_ (.Y(_3511_),
    .B1(_3503_),
    .B2(net2052),
    .A2(net880),
    .A1(_3455_));
 sg13g2_nor2_1 _7769_ (.A(net1110),
    .B(_3511_),
    .Y(_0663_));
 sg13g2_nand3b_1 _7770_ (.B(_3420_),
    .C(net1003),
    .Y(_3512_),
    .A_N(net1139));
 sg13g2_a22oi_1 _7771_ (.Y(_3513_),
    .B1(_3512_),
    .B2(net2070),
    .A2(net884),
    .A1(_3458_));
 sg13g2_nand2_1 _7772_ (.Y(_0664_),
    .A(net1160),
    .B(net2071));
 sg13g2_a22oi_1 _7773_ (.Y(_3514_),
    .B1(_3512_),
    .B2(net2296),
    .A2(net882),
    .A1(_3461_));
 sg13g2_nand2_1 _7774_ (.Y(_0665_),
    .A(net1157),
    .B(_3514_));
 sg13g2_a22oi_1 _7775_ (.Y(_3515_),
    .B1(_3512_),
    .B2(net2145),
    .A2(net883),
    .A1(_3463_));
 sg13g2_nand2_1 _7776_ (.Y(_0666_),
    .A(net1160),
    .B(_3515_));
 sg13g2_a22oi_1 _7777_ (.Y(_3516_),
    .B1(_3512_),
    .B2(net2245),
    .A2(net882),
    .A1(_3465_));
 sg13g2_nand2_1 _7778_ (.Y(_0667_),
    .A(net1160),
    .B(_3516_));
 sg13g2_a22oi_1 _7779_ (.Y(_3517_),
    .B1(_3512_),
    .B2(net2173),
    .A2(net884),
    .A1(_3467_));
 sg13g2_nand2_1 _7780_ (.Y(_0668_),
    .A(net1156),
    .B(_3517_));
 sg13g2_a22oi_1 _7781_ (.Y(_3518_),
    .B1(_3512_),
    .B2(net2274),
    .A2(net880),
    .A1(_3469_));
 sg13g2_nand2_1 _7782_ (.Y(_0669_),
    .A(net1152),
    .B(_3518_));
 sg13g2_a22oi_1 _7783_ (.Y(_3519_),
    .B1(_3512_),
    .B2(net2048),
    .A2(net881),
    .A1(_3471_));
 sg13g2_nand2_1 _7784_ (.Y(_0670_),
    .A(net1156),
    .B(net2049));
 sg13g2_a22oi_1 _7785_ (.Y(_3520_),
    .B1(_3512_),
    .B2(net2244),
    .A2(net880),
    .A1(_3473_));
 sg13g2_nand2_1 _7786_ (.Y(_0671_),
    .A(net1152),
    .B(_3520_));
 sg13g2_nand2_2 _7787_ (.Y(_3521_),
    .A(net1002),
    .B(net881));
 sg13g2_a22oi_1 _7788_ (.Y(_3522_),
    .B1(_3521_),
    .B2(net1750),
    .A2(net884),
    .A1(_3477_));
 sg13g2_nor2_1 _7789_ (.A(net1123),
    .B(net1751),
    .Y(_0672_));
 sg13g2_a22oi_1 _7790_ (.Y(_3523_),
    .B1(_3521_),
    .B2(net1832),
    .A2(net882),
    .A1(_3479_));
 sg13g2_nor2_1 _7791_ (.A(net1118),
    .B(net1833),
    .Y(_0673_));
 sg13g2_a22oi_1 _7792_ (.Y(_3524_),
    .B1(_3521_),
    .B2(net1693),
    .A2(net882),
    .A1(_3481_));
 sg13g2_nor2_1 _7793_ (.A(net1118),
    .B(net1694),
    .Y(_0674_));
 sg13g2_a22oi_1 _7794_ (.Y(_3525_),
    .B1(_3521_),
    .B2(net1885),
    .A2(net883),
    .A1(_3483_));
 sg13g2_nor2_1 _7795_ (.A(net1118),
    .B(net1886),
    .Y(_0675_));
 sg13g2_a22oi_1 _7796_ (.Y(_3526_),
    .B1(_3521_),
    .B2(net1814),
    .A2(net885),
    .A1(_3485_));
 sg13g2_nor2_1 _7797_ (.A(net1124),
    .B(net1815),
    .Y(_0676_));
 sg13g2_a22oi_1 _7798_ (.Y(_3527_),
    .B1(_3521_),
    .B2(net1914),
    .A2(net881),
    .A1(_3487_));
 sg13g2_nor2_1 _7799_ (.A(net1108),
    .B(net1915),
    .Y(_0677_));
 sg13g2_a22oi_1 _7800_ (.Y(_3528_),
    .B1(_3521_),
    .B2(net1773),
    .A2(net880),
    .A1(_3489_));
 sg13g2_nor2_1 _7801_ (.A(net1113),
    .B(net1774),
    .Y(_0678_));
 sg13g2_a22oi_1 _7802_ (.Y(_3529_),
    .B1(_3521_),
    .B2(net1866),
    .A2(net880),
    .A1(_3491_));
 sg13g2_nor2_1 _7803_ (.A(net1112),
    .B(net1867),
    .Y(_0679_));
 sg13g2_nor2_1 _7804_ (.A(_3389_),
    .B(_3410_),
    .Y(_3530_));
 sg13g2_nand3_1 _7805_ (.B(_3260_),
    .C(_3530_),
    .A(net1138),
    .Y(_3531_));
 sg13g2_nor3_2 _7806_ (.A(net1136),
    .B(_3386_),
    .C(_3410_),
    .Y(_3532_));
 sg13g2_a22oi_1 _7807_ (.Y(_3533_),
    .B1(net879),
    .B2(_3422_),
    .A2(_3531_),
    .A1(net1987));
 sg13g2_nor2_1 _7808_ (.A(net1123),
    .B(net1988),
    .Y(_0680_));
 sg13g2_a22oi_1 _7809_ (.Y(_3534_),
    .B1(net878),
    .B2(_3426_),
    .A2(_3531_),
    .A1(net2133));
 sg13g2_nor2_1 _7810_ (.A(net1119),
    .B(net2134),
    .Y(_0681_));
 sg13g2_a22oi_1 _7811_ (.Y(_3535_),
    .B1(net878),
    .B2(_3428_),
    .A2(_3531_),
    .A1(net2044));
 sg13g2_nor2_1 _7812_ (.A(net1108),
    .B(net2045),
    .Y(_0682_));
 sg13g2_a22oi_1 _7813_ (.Y(_3536_),
    .B1(net878),
    .B2(_3430_),
    .A2(_3531_),
    .A1(net2053));
 sg13g2_nor2_1 _7814_ (.A(net1118),
    .B(net2054),
    .Y(_0683_));
 sg13g2_a22oi_1 _7815_ (.Y(_3537_),
    .B1(net879),
    .B2(_3432_),
    .A2(_3531_),
    .A1(net1922));
 sg13g2_nor2_1 _7816_ (.A(net1124),
    .B(net1923),
    .Y(_0684_));
 sg13g2_a22oi_1 _7817_ (.Y(_3538_),
    .B1(net877),
    .B2(_3434_),
    .A2(_3531_),
    .A1(net2207));
 sg13g2_nor2_1 _7818_ (.A(net1110),
    .B(_3538_),
    .Y(_0685_));
 sg13g2_a22oi_1 _7819_ (.Y(_3539_),
    .B1(net877),
    .B2(_3436_),
    .A2(_3531_),
    .A1(net2007));
 sg13g2_nor2_1 _7820_ (.A(net1113),
    .B(net2008),
    .Y(_0686_));
 sg13g2_a22oi_1 _7821_ (.Y(_3540_),
    .B1(net877),
    .B2(_3438_),
    .A2(_3531_),
    .A1(net2251));
 sg13g2_nor2_1 _7822_ (.A(net1110),
    .B(_3540_),
    .Y(_0687_));
 sg13g2_nand3_1 _7823_ (.B(net1004),
    .C(_3530_),
    .A(net1139),
    .Y(_3541_));
 sg13g2_a22oi_1 _7824_ (.Y(_3542_),
    .B1(_3541_),
    .B2(net2032),
    .A2(net879),
    .A1(_3440_));
 sg13g2_nand2_1 _7825_ (.Y(_0688_),
    .A(net1160),
    .B(net2033));
 sg13g2_a22oi_1 _7826_ (.Y(_3543_),
    .B1(_3541_),
    .B2(net2249),
    .A2(net878),
    .A1(_3443_));
 sg13g2_nand2_1 _7827_ (.Y(_0689_),
    .A(net1158),
    .B(_3543_));
 sg13g2_a22oi_1 _7828_ (.Y(_3544_),
    .B1(_3541_),
    .B2(net2265),
    .A2(net878),
    .A1(_3445_));
 sg13g2_nand2_1 _7829_ (.Y(_0690_),
    .A(net1160),
    .B(_3544_));
 sg13g2_a22oi_1 _7830_ (.Y(_3545_),
    .B1(_3541_),
    .B2(net2215),
    .A2(net879),
    .A1(_3447_));
 sg13g2_nand2_1 _7831_ (.Y(_0691_),
    .A(net1157),
    .B(_3545_));
 sg13g2_a22oi_1 _7832_ (.Y(_3546_),
    .B1(_3541_),
    .B2(net2165),
    .A2(net879),
    .A1(_3449_));
 sg13g2_nand2_1 _7833_ (.Y(_0692_),
    .A(net1160),
    .B(_3546_));
 sg13g2_a22oi_1 _7834_ (.Y(_3547_),
    .B1(_3541_),
    .B2(net2166),
    .A2(net877),
    .A1(_3451_));
 sg13g2_nand2_1 _7835_ (.Y(_0693_),
    .A(net1150),
    .B(_3547_));
 sg13g2_a22oi_1 _7836_ (.Y(_3548_),
    .B1(_3541_),
    .B2(net2126),
    .A2(net877),
    .A1(_3453_));
 sg13g2_nand2_1 _7837_ (.Y(_0694_),
    .A(net1155),
    .B(net2127));
 sg13g2_a22oi_1 _7838_ (.Y(_3549_),
    .B1(_3541_),
    .B2(net2151),
    .A2(net877),
    .A1(_3455_));
 sg13g2_nand2_1 _7839_ (.Y(_0695_),
    .A(net1151),
    .B(_3549_));
 sg13g2_nand3_1 _7840_ (.B(net1003),
    .C(_3530_),
    .A(net1139),
    .Y(_3550_));
 sg13g2_a22oi_1 _7841_ (.Y(_3551_),
    .B1(_3550_),
    .B2(net1854),
    .A2(net879),
    .A1(_3458_));
 sg13g2_nor2_1 _7842_ (.A(net1123),
    .B(net1855),
    .Y(_0696_));
 sg13g2_a22oi_1 _7843_ (.Y(_3552_),
    .B1(_3550_),
    .B2(net1975),
    .A2(net878),
    .A1(_3461_));
 sg13g2_nor2_1 _7844_ (.A(net1122),
    .B(net1976),
    .Y(_0697_));
 sg13g2_a22oi_1 _7845_ (.Y(_3553_),
    .B1(_3550_),
    .B2(net2038),
    .A2(net878),
    .A1(_3463_));
 sg13g2_nor2_1 _7846_ (.A(net1123),
    .B(net2039),
    .Y(_0698_));
 sg13g2_a22oi_1 _7847_ (.Y(_3554_),
    .B1(_3550_),
    .B2(net2011),
    .A2(net878),
    .A1(_3465_));
 sg13g2_nor2_1 _7848_ (.A(net1119),
    .B(_3554_),
    .Y(_0699_));
 sg13g2_a22oi_1 _7849_ (.Y(_3555_),
    .B1(_3550_),
    .B2(net1788),
    .A2(net879),
    .A1(_3467_));
 sg13g2_nor2_1 _7850_ (.A(net1124),
    .B(net1789),
    .Y(_0700_));
 sg13g2_a22oi_1 _7851_ (.Y(_3556_),
    .B1(_3550_),
    .B2(net1919),
    .A2(net877),
    .A1(_3469_));
 sg13g2_nor2_1 _7852_ (.A(net1112),
    .B(net1920),
    .Y(_0701_));
 sg13g2_a22oi_1 _7853_ (.Y(_3557_),
    .B1(_3550_),
    .B2(net1868),
    .A2(_3532_),
    .A1(_3471_));
 sg13g2_nor2_1 _7854_ (.A(net1112),
    .B(net1869),
    .Y(_0702_));
 sg13g2_a22oi_1 _7855_ (.Y(_3558_),
    .B1(_3550_),
    .B2(net1848),
    .A2(net877),
    .A1(_3473_));
 sg13g2_nor2_1 _7856_ (.A(net1112),
    .B(net1849),
    .Y(_0703_));
 sg13g2_and2_1 _7857_ (.A(_3217_),
    .B(net954),
    .X(_3559_));
 sg13g2_nand2_2 _7858_ (.Y(_3560_),
    .A(_3217_),
    .B(_3264_));
 sg13g2_o21ai_1 _7859_ (.B1(net1147),
    .Y(_3561_),
    .A1(net2326),
    .A2(_3559_));
 sg13g2_a21oi_1 _7860_ (.A1(_0747_),
    .A2(_3559_),
    .Y(_0704_),
    .B1(_3561_));
 sg13g2_a21oi_1 _7861_ (.A1(net2252),
    .A2(_3560_),
    .Y(_3562_),
    .B1(net1106));
 sg13g2_o21ai_1 _7862_ (.B1(_3562_),
    .Y(_0705_),
    .A1(_0746_),
    .A2(_3560_));
 sg13g2_a21oi_1 _7863_ (.A1(net2300),
    .A2(_3560_),
    .Y(_3563_),
    .B1(net1107));
 sg13g2_o21ai_1 _7864_ (.B1(_3563_),
    .Y(_0706_),
    .A1(_0745_),
    .A2(_3560_));
 sg13g2_a21oi_1 _7865_ (.A1(net2208),
    .A2(_3560_),
    .Y(_3564_),
    .B1(net1107));
 sg13g2_o21ai_1 _7866_ (.B1(_3564_),
    .Y(_0707_),
    .A1(_0744_),
    .A2(_3560_));
 sg13g2_a21oi_1 _7867_ (.A1(net2201),
    .A2(_3560_),
    .Y(_3565_),
    .B1(net1107));
 sg13g2_o21ai_1 _7868_ (.B1(_3565_),
    .Y(_0708_),
    .A1(_0743_),
    .A2(_3560_));
 sg13g2_o21ai_1 _7869_ (.B1(net1147),
    .Y(_3566_),
    .A1(net2086),
    .A2(_3559_));
 sg13g2_a21oi_1 _7870_ (.A1(_0742_),
    .A2(_3559_),
    .Y(_0709_),
    .B1(_3566_));
 sg13g2_o21ai_1 _7871_ (.B1(net1147),
    .Y(_3567_),
    .A1(net2168),
    .A2(_3559_));
 sg13g2_a21oi_1 _7872_ (.A1(_0741_),
    .A2(_3559_),
    .Y(_0710_),
    .B1(_3567_));
 sg13g2_o21ai_1 _7873_ (.B1(net1147),
    .Y(_3568_),
    .A1(\led_controller.cpu.i_num_leds[7] ),
    .A2(_3559_));
 sg13g2_a21oi_1 _7874_ (.A1(_0740_),
    .A2(_3559_),
    .Y(_0711_),
    .B1(_3568_));
 sg13g2_and2_1 _7875_ (.A(_3217_),
    .B(_3256_),
    .X(_3569_));
 sg13g2_a21oi_1 _7876_ (.A1(\led_controller.register_data[0] ),
    .A2(_3569_),
    .Y(_3570_),
    .B1(net1120));
 sg13g2_o21ai_1 _7877_ (.B1(_3570_),
    .Y(_0712_),
    .A1(_0748_),
    .A2(_3569_));
 sg13g2_o21ai_1 _7878_ (.B1(net1148),
    .Y(_3571_),
    .A1(net2137),
    .A2(_3569_));
 sg13g2_a21oi_1 _7879_ (.A1(_0746_),
    .A2(_3569_),
    .Y(_0713_),
    .B1(_3571_));
 sg13g2_o21ai_1 _7880_ (.B1(net1148),
    .Y(_3572_),
    .A1(net2118),
    .A2(_3569_));
 sg13g2_a21oi_1 _7881_ (.A1(_0745_),
    .A2(_3569_),
    .Y(_0714_),
    .B1(_3572_));
 sg13g2_o21ai_1 _7882_ (.B1(net1148),
    .Y(_3573_),
    .A1(net2059),
    .A2(_3569_));
 sg13g2_a21oi_1 _7883_ (.A1(_0744_),
    .A2(_3569_),
    .Y(_0715_),
    .B1(_3573_));
 sg13g2_nor3_1 _7884_ (.A(_3218_),
    .B(net1062),
    .C(_3258_),
    .Y(_3574_));
 sg13g2_nand2_2 _7885_ (.Y(_3575_),
    .A(_3217_),
    .B(net955));
 sg13g2_a21oi_1 _7886_ (.A1(net2341),
    .A2(_3575_),
    .Y(_3576_),
    .B1(net1106));
 sg13g2_o21ai_1 _7887_ (.B1(_3576_),
    .Y(_0716_),
    .A1(_0747_),
    .A2(_3575_));
 sg13g2_o21ai_1 _7888_ (.B1(net1147),
    .Y(_3577_),
    .A1(net2195),
    .A2(net952));
 sg13g2_a21oi_1 _7889_ (.A1(_0746_),
    .A2(net952),
    .Y(_0717_),
    .B1(_3577_));
 sg13g2_a21oi_1 _7890_ (.A1(net2187),
    .A2(_3575_),
    .Y(_3578_),
    .B1(net1120));
 sg13g2_o21ai_1 _7891_ (.B1(_3578_),
    .Y(_0718_),
    .A1(_0745_),
    .A2(_3575_));
 sg13g2_o21ai_1 _7892_ (.B1(net1146),
    .Y(_3579_),
    .A1(net2144),
    .A2(net952));
 sg13g2_a21oi_1 _7893_ (.A1(_0744_),
    .A2(net953),
    .Y(_0719_),
    .B1(_3579_));
 sg13g2_o21ai_1 _7894_ (.B1(net1147),
    .Y(_3580_),
    .A1(net2132),
    .A2(net953));
 sg13g2_a21oi_1 _7895_ (.A1(_0743_),
    .A2(net953),
    .Y(_0720_),
    .B1(_3580_));
 sg13g2_o21ai_1 _7896_ (.B1(net1147),
    .Y(_3581_),
    .A1(net1995),
    .A2(net952));
 sg13g2_a21oi_1 _7897_ (.A1(_0742_),
    .A2(net952),
    .Y(_0721_),
    .B1(_3581_));
 sg13g2_o21ai_1 _7898_ (.B1(net1147),
    .Y(_3582_),
    .A1(net2185),
    .A2(net953));
 sg13g2_a21oi_1 _7899_ (.A1(_0741_),
    .A2(net952),
    .Y(_0722_),
    .B1(_3582_));
 sg13g2_o21ai_1 _7900_ (.B1(net1144),
    .Y(_3583_),
    .A1(net2111),
    .A2(net952));
 sg13g2_a21oi_1 _7901_ (.A1(_0740_),
    .A2(net952),
    .Y(_0723_),
    .B1(_3583_));
 sg13g2_nand3_1 _7902_ (.B(_1054_),
    .C(_1096_),
    .A(_1052_),
    .Y(_3584_));
 sg13g2_a21oi_2 _7903_ (.B1(net1033),
    .Y(_3585_),
    .A2(_1205_),
    .A1(_1052_));
 sg13g2_nand2_1 _7904_ (.Y(_3586_),
    .A(net820),
    .B(_3585_));
 sg13g2_o21ai_1 _7905_ (.B1(_3586_),
    .Y(_0724_),
    .A1(net936),
    .A2(_3584_));
 sg13g2_nand2_1 _7906_ (.Y(_3587_),
    .A(net1286),
    .B(_3585_));
 sg13g2_o21ai_1 _7907_ (.B1(_3587_),
    .Y(_0725_),
    .A1(net931),
    .A2(_3584_));
 sg13g2_nand2_1 _7908_ (.Y(_3588_),
    .A(net799),
    .B(_3585_));
 sg13g2_o21ai_1 _7909_ (.B1(_3588_),
    .Y(_0726_),
    .A1(net930),
    .A2(_3584_));
 sg13g2_nand2_1 _7910_ (.Y(_3589_),
    .A(net1225),
    .B(_3585_));
 sg13g2_o21ai_1 _7911_ (.B1(_3589_),
    .Y(_0727_),
    .A1(net928),
    .A2(_3584_));
 sg13g2_nand2_1 _7912_ (.Y(_3590_),
    .A(net1342),
    .B(_3585_));
 sg13g2_o21ai_1 _7913_ (.B1(_3590_),
    .Y(_0728_),
    .A1(net924),
    .A2(_3584_));
 sg13g2_nand2_1 _7914_ (.Y(_3591_),
    .A(net1261),
    .B(_3585_));
 sg13g2_o21ai_1 _7915_ (.B1(_3591_),
    .Y(_0729_),
    .A1(net923),
    .A2(_3584_));
 sg13g2_nand2_1 _7916_ (.Y(_3592_),
    .A(net1229),
    .B(_3585_));
 sg13g2_o21ai_1 _7917_ (.B1(_3592_),
    .Y(_0730_),
    .A1(net920),
    .A2(_3584_));
 sg13g2_nand2_1 _7918_ (.Y(_3593_),
    .A(net817),
    .B(_3585_));
 sg13g2_o21ai_1 _7919_ (.B1(_3593_),
    .Y(_0731_),
    .A1(net916),
    .A2(_3584_));
 sg13g2_nand2_2 _7920_ (.Y(_3594_),
    .A(_1052_),
    .B(_1127_));
 sg13g2_a21oi_2 _7921_ (.B1(net1031),
    .Y(_3595_),
    .A2(_1127_),
    .A1(_1052_));
 sg13g2_nand2_1 _7922_ (.Y(_3596_),
    .A(net1303),
    .B(_3595_));
 sg13g2_o21ai_1 _7923_ (.B1(_3596_),
    .Y(_0732_),
    .A1(net935),
    .A2(_3594_));
 sg13g2_nand2_1 _7924_ (.Y(_3597_),
    .A(net1243),
    .B(_3595_));
 sg13g2_o21ai_1 _7925_ (.B1(_3597_),
    .Y(_0733_),
    .A1(net932),
    .A2(_3594_));
 sg13g2_nand2_1 _7926_ (.Y(_3598_),
    .A(net1268),
    .B(_3595_));
 sg13g2_o21ai_1 _7927_ (.B1(_3598_),
    .Y(_0734_),
    .A1(net929),
    .A2(_3594_));
 sg13g2_nand2_1 _7928_ (.Y(_3599_),
    .A(net1277),
    .B(_3595_));
 sg13g2_o21ai_1 _7929_ (.B1(_3599_),
    .Y(_0735_),
    .A1(net926),
    .A2(_3594_));
 sg13g2_nand2_1 _7930_ (.Y(_3600_),
    .A(net1258),
    .B(_3595_));
 sg13g2_o21ai_1 _7931_ (.B1(_3600_),
    .Y(_0736_),
    .A1(net924),
    .A2(_3594_));
 sg13g2_nand2_1 _7932_ (.Y(_3601_),
    .A(net1256),
    .B(_3595_));
 sg13g2_o21ai_1 _7933_ (.B1(_3601_),
    .Y(_0737_),
    .A1(net921),
    .A2(_3594_));
 sg13g2_nand2_1 _7934_ (.Y(_3602_),
    .A(net1315),
    .B(_3595_));
 sg13g2_o21ai_1 _7935_ (.B1(_3602_),
    .Y(_0738_),
    .A1(net918),
    .A2(_3594_));
 sg13g2_nand2_1 _7936_ (.Y(_3603_),
    .A(net1231),
    .B(_3595_));
 sg13g2_o21ai_1 _7937_ (.B1(_3603_),
    .Y(_0739_),
    .A1(net917),
    .A2(_3594_));
 sg13g2_a21oi_1 _7938_ (.A1(_0855_),
    .A2(net947),
    .Y(_0351_),
    .B1(_1046_));
 sg13g2_a21oi_1 _7939_ (.A1(_0854_),
    .A2(net946),
    .Y(_0352_),
    .B1(_1047_));
 sg13g2_a21oi_1 _7940_ (.A1(_0853_),
    .A2(net946),
    .Y(_0353_),
    .B1(_1048_));
 sg13g2_a21oi_1 _7941_ (.A1(_0852_),
    .A2(net946),
    .Y(_0354_),
    .B1(_1049_));
 sg13g2_dfrbpq_2 _7942_ (.RESET_B(net24),
    .D(_0019_),
    .Q(\led_controller.led_effect_pulse.fade_out ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _7943_ (.RESET_B(net69),
    .D(net1710),
    .Q(\led_controller.led_effect_pulse.state[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _7944_ (.RESET_B(net759),
    .D(net1381),
    .Q(\led_controller.led_effect_pulse.state[1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _7945_ (.RESET_B(net647),
    .D(_0020_),
    .Q(_0000_),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _7946_ (.RESET_B(net646),
    .D(_0021_),
    .Q(_0001_),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _7947_ (.RESET_B(net645),
    .D(_0022_),
    .Q(_0002_),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _7948_ (.RESET_B(net644),
    .D(_0023_),
    .Q(_0003_),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _7949_ (.RESET_B(net643),
    .D(_0024_),
    .Q(\led_controller.cpu.scratch_memory[14][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7950_ (.RESET_B(net641),
    .D(_0025_),
    .Q(\led_controller.cpu.scratch_memory[14][1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7951_ (.RESET_B(net639),
    .D(_0026_),
    .Q(\led_controller.cpu.scratch_memory[14][2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _7952_ (.RESET_B(net637),
    .D(_0027_),
    .Q(\led_controller.cpu.scratch_memory[14][3] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7953_ (.RESET_B(net635),
    .D(_0028_),
    .Q(\led_controller.cpu.scratch_memory[14][4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7954_ (.RESET_B(net633),
    .D(net1534),
    .Q(\led_controller.cpu.scratch_memory[14][5] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _7955_ (.RESET_B(net631),
    .D(_0030_),
    .Q(\led_controller.cpu.scratch_memory[14][6] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7956_ (.RESET_B(net629),
    .D(_0031_),
    .Q(\led_controller.cpu.scratch_memory[14][7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7957_ (.RESET_B(net627),
    .D(net1311),
    .Q(\led_controller.cpu.scratch_memory[9][0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7958_ (.RESET_B(net625),
    .D(net1240),
    .Q(\led_controller.cpu.scratch_memory[9][1] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _7959_ (.RESET_B(net623),
    .D(net801),
    .Q(\led_controller.cpu.scratch_memory[9][2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7960_ (.RESET_B(net621),
    .D(net1242),
    .Q(\led_controller.cpu.scratch_memory[9][3] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7961_ (.RESET_B(net619),
    .D(net1285),
    .Q(\led_controller.cpu.scratch_memory[9][4] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7962_ (.RESET_B(net617),
    .D(net1251),
    .Q(\led_controller.cpu.scratch_memory[9][5] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7963_ (.RESET_B(net615),
    .D(net1291),
    .Q(\led_controller.cpu.scratch_memory[9][6] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7964_ (.RESET_B(net613),
    .D(net794),
    .Q(\led_controller.cpu.scratch_memory[9][7] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7965_ (.RESET_B(net611),
    .D(net1298),
    .Q(\led_controller.cpu.scratch_memory[11][0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7966_ (.RESET_B(net609),
    .D(net1227),
    .Q(\led_controller.cpu.scratch_memory[11][1] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7967_ (.RESET_B(net607),
    .D(net804),
    .Q(\led_controller.cpu.scratch_memory[11][2] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _7968_ (.RESET_B(net605),
    .D(net1264),
    .Q(\led_controller.cpu.scratch_memory[11][3] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7969_ (.RESET_B(net603),
    .D(net813),
    .Q(\led_controller.cpu.scratch_memory[11][4] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7970_ (.RESET_B(net601),
    .D(net1362),
    .Q(\led_controller.cpu.scratch_memory[11][5] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7971_ (.RESET_B(net599),
    .D(net1365),
    .Q(\led_controller.cpu.scratch_memory[11][6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7972_ (.RESET_B(net597),
    .D(net1302),
    .Q(\led_controller.cpu.scratch_memory[11][7] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7973_ (.RESET_B(net595),
    .D(net807),
    .Q(\led_controller.cpu.scratch_memory[10][0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7974_ (.RESET_B(net591),
    .D(net1328),
    .Q(\led_controller.cpu.scratch_memory[10][1] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _7975_ (.RESET_B(net589),
    .D(net768),
    .Q(\led_controller.cpu.scratch_memory[10][2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7976_ (.RESET_B(net587),
    .D(net778),
    .Q(\led_controller.cpu.scratch_memory[10][3] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7977_ (.RESET_B(net585),
    .D(net1332),
    .Q(\led_controller.cpu.scratch_memory[10][4] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7978_ (.RESET_B(net583),
    .D(net1388),
    .Q(\led_controller.cpu.scratch_memory[10][5] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7979_ (.RESET_B(net581),
    .D(net797),
    .Q(\led_controller.cpu.scratch_memory[10][6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7980_ (.RESET_B(net579),
    .D(net774),
    .Q(\led_controller.cpu.scratch_memory[10][7] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _7981_ (.RESET_B(net577),
    .D(_0056_),
    .Q(\led_controller.cpu.scratch_memory[5][0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _7982_ (.RESET_B(net575),
    .D(_0057_),
    .Q(\led_controller.cpu.scratch_memory[5][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _7983_ (.RESET_B(net573),
    .D(_0058_),
    .Q(\led_controller.cpu.scratch_memory[5][2] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7984_ (.RESET_B(net571),
    .D(_0059_),
    .Q(\led_controller.cpu.scratch_memory[5][3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _7985_ (.RESET_B(net569),
    .D(_0060_),
    .Q(\led_controller.cpu.scratch_memory[5][4] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7986_ (.RESET_B(net567),
    .D(_0061_),
    .Q(\led_controller.cpu.scratch_memory[5][5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7987_ (.RESET_B(net565),
    .D(_0062_),
    .Q(\led_controller.cpu.scratch_memory[5][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _7988_ (.RESET_B(net70),
    .D(_0063_),
    .Q(\led_controller.cpu.scratch_memory[5][7] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _7989_ (.RESET_B(net71),
    .D(net1827),
    .Q(\led_controller.spi_state[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _7990_ (.RESET_B(net96),
    .D(_0017_),
    .Q(\led_controller.spi_state[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _7991_ (.RESET_B(net563),
    .D(_0018_),
    .Q(\led_controller.spi_state[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _7992_ (.RESET_B(net561),
    .D(_0064_),
    .Q(\led_controller.timer_100hz.div_counter[0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _7993_ (.RESET_B(net560),
    .D(_0065_),
    .Q(\led_controller.timer_100hz.div_counter[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _7994_ (.RESET_B(net559),
    .D(net1516),
    .Q(\led_controller.timer_100hz.div_counter[2] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _7995_ (.RESET_B(net558),
    .D(_0067_),
    .Q(\led_controller.timer_100hz.div_counter[3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7996_ (.RESET_B(net557),
    .D(net1795),
    .Q(\led_controller.timer_100hz.div_counter[4] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7997_ (.RESET_B(net556),
    .D(_0069_),
    .Q(\led_controller.timer_100hz.div_counter[5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _7998_ (.RESET_B(net555),
    .D(_0070_),
    .Q(\led_controller.timer_100hz.div_counter[6] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7999_ (.RESET_B(net554),
    .D(_0071_),
    .Q(\led_controller.timer_100hz.div_counter[7] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _8000_ (.RESET_B(net553),
    .D(_0072_),
    .Q(\led_controller.cpu.scratch_memory[4][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _8001_ (.RESET_B(net551),
    .D(_0073_),
    .Q(\led_controller.cpu.scratch_memory[4][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _8002_ (.RESET_B(net549),
    .D(_0074_),
    .Q(\led_controller.cpu.scratch_memory[4][2] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _8003_ (.RESET_B(net547),
    .D(_0075_),
    .Q(\led_controller.cpu.scratch_memory[4][3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _8004_ (.RESET_B(net545),
    .D(_0076_),
    .Q(\led_controller.cpu.scratch_memory[4][4] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _8005_ (.RESET_B(net543),
    .D(_0077_),
    .Q(\led_controller.cpu.scratch_memory[4][5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _8006_ (.RESET_B(net541),
    .D(_0078_),
    .Q(\led_controller.cpu.scratch_memory[4][6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _8007_ (.RESET_B(net539),
    .D(_0079_),
    .Q(\led_controller.cpu.scratch_memory[4][7] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8008_ (.RESET_B(net537),
    .D(net1348),
    .Q(\led_controller.cpu.scratch_memory[3][0] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8009_ (.RESET_B(net535),
    .D(_0081_),
    .Q(\led_controller.cpu.scratch_memory[3][1] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8010_ (.RESET_B(net533),
    .D(_0082_),
    .Q(\led_controller.cpu.scratch_memory[3][2] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8011_ (.RESET_B(net531),
    .D(_0083_),
    .Q(\led_controller.cpu.scratch_memory[3][3] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _8012_ (.RESET_B(net529),
    .D(_0084_),
    .Q(\led_controller.cpu.scratch_memory[3][4] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8013_ (.RESET_B(net527),
    .D(_0085_),
    .Q(\led_controller.cpu.scratch_memory[3][5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8014_ (.RESET_B(net526),
    .D(_0086_),
    .Q(\led_controller.cpu.scratch_memory[3][6] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8015_ (.RESET_B(net97),
    .D(_0087_),
    .Q(\led_controller.cpu.scratch_memory[3][7] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8016_ (.RESET_B(net98),
    .D(net1577),
    .Q(\led_controller.flash.state[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _8017_ (.RESET_B(net99),
    .D(_0005_),
    .Q(\led_controller.flash.state[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8018_ (.RESET_B(net100),
    .D(net1502),
    .Q(\led_controller.flash.state[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8019_ (.RESET_B(net101),
    .D(net1530),
    .Q(\led_controller.flash.state[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8020_ (.RESET_B(net102),
    .D(_0008_),
    .Q(\led_controller.flash.state[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8021_ (.RESET_B(net103),
    .D(_0009_),
    .Q(\led_controller.flash.state[5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _8022_ (.RESET_B(net104),
    .D(net2078),
    .Q(\led_controller.flash.state[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _8023_ (.RESET_B(net105),
    .D(net1877),
    .Q(\led_controller.rgbw.state[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _8024_ (.RESET_B(net593),
    .D(_0014_),
    .Q(\led_controller.rgbw.state[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _8025_ (.RESET_B(net524),
    .D(net2354),
    .Q(\led_controller.rgbw.state[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _8026_ (.RESET_B(net522),
    .D(_0088_),
    .Q(\led_controller.cpu.scratch_memory[12][0] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _8027_ (.RESET_B(net520),
    .D(_0089_),
    .Q(\led_controller.cpu.scratch_memory[12][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8028_ (.RESET_B(net518),
    .D(_0090_),
    .Q(\led_controller.cpu.scratch_memory[12][2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8029_ (.RESET_B(net516),
    .D(_0091_),
    .Q(\led_controller.cpu.scratch_memory[12][3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _8030_ (.RESET_B(net514),
    .D(_0092_),
    .Q(\led_controller.cpu.scratch_memory[12][4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8031_ (.RESET_B(net512),
    .D(_0093_),
    .Q(\led_controller.cpu.scratch_memory[12][5] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _8032_ (.RESET_B(net510),
    .D(_0094_),
    .Q(\led_controller.cpu.scratch_memory[12][6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8033_ (.RESET_B(net508),
    .D(_0095_),
    .Q(\led_controller.cpu.scratch_memory[12][7] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _8034_ (.RESET_B(net506),
    .D(net2340),
    .Q(\led_controller.cpu.fetch_pc[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _8035_ (.RESET_B(net504),
    .D(net2217),
    .Q(\led_controller.cpu.fetch_pc[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _8036_ (.RESET_B(net502),
    .D(net2010),
    .Q(\led_controller.cpu.fetch_pc[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _8037_ (.RESET_B(net500),
    .D(net2156),
    .Q(\led_controller.cpu.fetch_pc[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _8038_ (.RESET_B(net498),
    .D(net2227),
    .Q(\led_controller.cpu.fetch_pc[5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8039_ (.RESET_B(net496),
    .D(net1925),
    .Q(\led_controller.cpu.fetch_pc[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _8040_ (.RESET_B(net494),
    .D(net1835),
    .Q(\led_controller.cpu.fetch_pc[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _8041_ (.RESET_B(net492),
    .D(net1905),
    .Q(\led_controller.cpu.fetch_pc[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _8042_ (.RESET_B(net490),
    .D(net1875),
    .Q(\led_controller.cpu.fetch_pc[9] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _8043_ (.RESET_B(net488),
    .D(_0105_),
    .Q(\led_controller.cpu.fetch_pc[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8044_ (.RESET_B(net486),
    .D(net1839),
    .Q(\led_controller.cpu.fetch_pc[11] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _8045_ (.RESET_B(net484),
    .D(net2273),
    .Q(\led_controller.cpu.fetch_pc[12] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _8046_ (.RESET_B(net482),
    .D(net2225),
    .Q(\led_controller.cpu.fetch_pc[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8047_ (.RESET_B(net480),
    .D(net1918),
    .Q(\led_controller.cpu.fetch_pc[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8048_ (.RESET_B(net478),
    .D(_0110_),
    .Q(\led_controller.cpu.fetch_pc[15] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _8049_ (.RESET_B(net476),
    .D(_0111_),
    .Q(\led_controller.cpu.scratch_memory[6][0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8050_ (.RESET_B(net474),
    .D(_0112_),
    .Q(\led_controller.cpu.scratch_memory[6][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _8051_ (.RESET_B(net472),
    .D(_0113_),
    .Q(\led_controller.cpu.scratch_memory[6][2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8052_ (.RESET_B(net470),
    .D(_0114_),
    .Q(\led_controller.cpu.scratch_memory[6][3] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _8053_ (.RESET_B(net468),
    .D(_0115_),
    .Q(\led_controller.cpu.scratch_memory[6][4] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8054_ (.RESET_B(net466),
    .D(_0116_),
    .Q(\led_controller.cpu.scratch_memory[6][5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _8055_ (.RESET_B(net464),
    .D(_0117_),
    .Q(\led_controller.cpu.scratch_memory[6][6] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8056_ (.RESET_B(net462),
    .D(_0118_),
    .Q(\led_controller.cpu.scratch_memory[6][7] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _8057_ (.RESET_B(net460),
    .D(_0119_),
    .Q(\led_controller.cpu.scratch_memory[1][0] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8058_ (.RESET_B(net458),
    .D(_0120_),
    .Q(\led_controller.cpu.scratch_memory[1][1] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8059_ (.RESET_B(net456),
    .D(_0121_),
    .Q(\led_controller.cpu.scratch_memory[1][2] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8060_ (.RESET_B(net454),
    .D(_0122_),
    .Q(\led_controller.cpu.scratch_memory[1][3] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8061_ (.RESET_B(net452),
    .D(_0123_),
    .Q(\led_controller.cpu.scratch_memory[1][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8062_ (.RESET_B(net450),
    .D(_0124_),
    .Q(\led_controller.cpu.scratch_memory[1][5] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _8063_ (.RESET_B(net448),
    .D(_0125_),
    .Q(\led_controller.cpu.scratch_memory[1][6] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8064_ (.RESET_B(net446),
    .D(_0126_),
    .Q(\led_controller.cpu.scratch_memory[1][7] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _8065_ (.RESET_B(net444),
    .D(net786),
    .Q(\led_controller.rgbw.counter[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _8066_ (.RESET_B(net443),
    .D(net1873),
    .Q(\led_controller.rgbw.counter[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _8067_ (.RESET_B(net442),
    .D(net1590),
    .Q(\led_controller.rgbw.counter[2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _8068_ (.RESET_B(net441),
    .D(net1725),
    .Q(\led_controller.rgbw.counter[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _8069_ (.RESET_B(net440),
    .D(net1802),
    .Q(\led_controller.rgbw.counter[4] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _8070_ (.RESET_B(net439),
    .D(net1829),
    .Q(\led_controller.rgbw.counter[5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _8071_ (.RESET_B(net438),
    .D(net1929),
    .Q(\led_controller.rgbw.counter[6] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _8072_ (.RESET_B(net437),
    .D(_0134_),
    .Q(\led_controller.rgbw.counter[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _8073_ (.RESET_B(net436),
    .D(_0135_),
    .Q(\led_controller.spi_slave.o_tx_start_strb ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _8074_ (.RESET_B(net435),
    .D(net1490),
    .Q(\led_controller.o_spi_miso ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8075_ (.RESET_B(net434),
    .D(net1495),
    .Q(\led_controller.spi_slave.data_bits[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8076_ (.RESET_B(net433),
    .D(_0138_),
    .Q(\led_controller.spi_slave.data_bits[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _8077_ (.RESET_B(net432),
    .D(net1889),
    .Q(\led_controller.spi_slave.data_bits[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _8078_ (.RESET_B(net431),
    .D(net1666),
    .Q(\led_controller.spi_slave.data_bits[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _8079_ (.RESET_B(net430),
    .D(_0141_),
    .Q(\led_controller.spi_data[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8080_ (.RESET_B(net429),
    .D(_0142_),
    .Q(\led_controller.spi_data[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8081_ (.RESET_B(net428),
    .D(_0143_),
    .Q(\led_controller.spi_data[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8082_ (.RESET_B(net427),
    .D(_0144_),
    .Q(\led_controller.spi_data[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8083_ (.RESET_B(net426),
    .D(_0145_),
    .Q(\led_controller.spi_data[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8084_ (.RESET_B(net425),
    .D(_0146_),
    .Q(\led_controller.spi_data[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8085_ (.RESET_B(net424),
    .D(_0147_),
    .Q(\led_controller.spi_data[6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8086_ (.RESET_B(net423),
    .D(_0148_),
    .Q(\led_controller.spi_data[7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _8087_ (.RESET_B(net422),
    .D(_0149_),
    .Q(\led_controller.spi_slave.output_register[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _8088_ (.RESET_B(net421),
    .D(net1429),
    .Q(\led_controller.spi_slave.output_register[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8089_ (.RESET_B(net420),
    .D(net1234),
    .Q(\led_controller.spi_slave.output_register[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _8090_ (.RESET_B(net419),
    .D(net1352),
    .Q(\led_controller.spi_slave.output_register[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _8091_ (.RESET_B(net418),
    .D(net1313),
    .Q(\led_controller.spi_slave.output_register[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _8092_ (.RESET_B(net417),
    .D(net782),
    .Q(\led_controller.spi_slave.output_register[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _8093_ (.RESET_B(net416),
    .D(net1394),
    .Q(\led_controller.spi_slave.output_register[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _8094_ (.RESET_B(net415),
    .D(net1336),
    .Q(\led_controller.spi_slave.output_register[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _8095_ (.RESET_B(net414),
    .D(_0157_),
    .Q(\led_controller.spi_slave.last_sck ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _8096_ (.RESET_B(net413),
    .D(_0158_),
    .Q(\led_controller.spi_slave.sck ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _8097_ (.RESET_B(net412),
    .D(_0159_),
    .Q(\led_controller.spi_slave.sync_mosi.data ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _8098_ (.RESET_B(net411),
    .D(_0160_),
    .Q(\led_controller.spi_slave.mosi ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8099_ (.RESET_B(net410),
    .D(_0161_),
    .Q(\led_controller.spi_slave.last_ss ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _8100_ (.RESET_B(net409),
    .D(_0162_),
    .Q(\led_controller.spi_slave.ss_n ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _8101_ (.RESET_B(net408),
    .D(_0163_),
    .Q(\led_controller.spi_slave.sync_sck.data ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8102_ (.RESET_B(net407),
    .D(net1715),
    .Q(\led_controller.timer_2hz.counter[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _8103_ (.RESET_B(net405),
    .D(net1407),
    .Q(\led_controller.timer_2hz.counter[1] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _8104_ (.RESET_B(net403),
    .D(net1632),
    .Q(\led_controller.timer_2hz.counter[2] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _8105_ (.RESET_B(net401),
    .D(_0167_),
    .Q(\led_controller.timer_2hz.counter[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _8106_ (.RESET_B(net399),
    .D(_0168_),
    .Q(\led_controller.timer_2hz.counter[4] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _8107_ (.RESET_B(net397),
    .D(_0169_),
    .Q(\led_controller.timer_2hz.counter[5] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _8108_ (.RESET_B(net395),
    .D(net1699),
    .Q(\led_controller.timer_10hz.counter[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _8109_ (.RESET_B(net393),
    .D(net1963),
    .Q(\led_controller.timer_10hz.counter[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _8110_ (.RESET_B(net391),
    .D(net1560),
    .Q(\led_controller.timer_10hz.counter[2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _8111_ (.RESET_B(net389),
    .D(_0173_),
    .Q(\led_controller.timer_10hz.counter[3] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _8112_ (.RESET_B(net387),
    .D(_0174_),
    .Q(\led_controller.spi_slave.sync_ss_n.data ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8113_ (.RESET_B(net386),
    .D(_0175_),
    .Q(\led_controller.timer_100hz.counter[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _8114_ (.RESET_B(net384),
    .D(net1772),
    .Q(\led_controller.timer_100hz.counter[1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _8115_ (.RESET_B(net382),
    .D(_0177_),
    .Q(\led_controller.timer_100hz.counter[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _8116_ (.RESET_B(net380),
    .D(_0178_),
    .Q(\led_controller.timer_100hz.counter[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _8117_ (.RESET_B(net378),
    .D(_0179_),
    .Q(\led_controller.timer_100hz.counter[4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _8118_ (.RESET_B(net376),
    .D(net2065),
    .Q(\led_controller.timer_100hz.counter[5] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _8119_ (.RESET_B(net374),
    .D(net2106),
    .Q(\led_controller.timer_100hz.counter[6] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _8120_ (.RESET_B(net372),
    .D(net2171),
    .Q(\led_controller.timer_100hz.counter[7] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _8121_ (.RESET_B(net370),
    .D(net2025),
    .Q(\led_controller.timer_100hz.counter[8] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _8122_ (.RESET_B(net368),
    .D(net1456),
    .Q(\led_controller.timer_100hz.counter[9] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _8123_ (.RESET_B(net366),
    .D(_0185_),
    .Q(\led_controller.timer_100hz.counter[10] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _8124_ (.RESET_B(net364),
    .D(_0186_),
    .Q(\led_controller.timer_100hz.counter[11] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _8125_ (.RESET_B(net362),
    .D(_0187_),
    .Q(\led_controller.timer_100hz.counter[12] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _8126_ (.RESET_B(net360),
    .D(net1897),
    .Q(\led_controller.timer_100hz.counter[13] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8127_ (.RESET_B(net358),
    .D(_0189_),
    .Q(\led_controller.timer_100hz.counter[14] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _8128_ (.RESET_B(net356),
    .D(_0190_),
    .Q(\led_controller.timer_100hz.counter[15] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8129_ (.RESET_B(net354),
    .D(net1935),
    .Q(\led_controller.timer_100hz.counter[16] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8130_ (.RESET_B(net352),
    .D(_0192_),
    .Q(\led_controller.timer_100hz.counter[17] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8131_ (.RESET_B(net350),
    .D(net2184),
    .Q(\led_controller.timer_100hz.counter[18] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8132_ (.RESET_B(net348),
    .D(net1902),
    .Q(\led_controller.timer_100hz.counter[19] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _8133_ (.RESET_B(net346),
    .D(_0195_),
    .Q(\led_controller.timer_100hz.counter[20] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _8134_ (.RESET_B(net344),
    .D(_0196_),
    .Q(\led_controller.timer_100hz.counter[21] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8135_ (.RESET_B(net342),
    .D(net1960),
    .Q(\led_controller.timer_100hz.counter[22] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8136_ (.RESET_B(net340),
    .D(net2260),
    .Q(\led_controller.timer_100hz.counter[23] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8137_ (.RESET_B(net338),
    .D(_0199_),
    .Q(\led_controller.timer_100hz.counter[24] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8138_ (.RESET_B(net336),
    .D(_0200_),
    .Q(\led_controller.timer_100hz.counter[25] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _8139_ (.RESET_B(net334),
    .D(net2176),
    .Q(\led_controller.timer_100hz.counter[26] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _8140_ (.RESET_B(net332),
    .D(_0202_),
    .Q(\led_controller.timer_100hz.counter[27] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _8141_ (.RESET_B(net330),
    .D(net1813),
    .Q(\led_controller.timer_100hz.counter[28] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _8142_ (.RESET_B(net328),
    .D(net2074),
    .Q(\led_controller.timer_100hz.counter[29] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _8143_ (.RESET_B(net326),
    .D(net1307),
    .Q(\led_controller.timer_100hz.counter[30] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _8144_ (.RESET_B(net324),
    .D(net1548),
    .Q(\led_controller.timer_100hz.counter[31] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _8145_ (.RESET_B(net322),
    .D(_0207_),
    .Q(\led_controller.cpu.i_timer_100hz ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _8146_ (.RESET_B(net321),
    .D(_0208_),
    .Q(\led_controller.cpu.scratch_memory[2][0] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8147_ (.RESET_B(net319),
    .D(_0209_),
    .Q(\led_controller.cpu.scratch_memory[2][1] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8148_ (.RESET_B(net317),
    .D(_0210_),
    .Q(\led_controller.cpu.scratch_memory[2][2] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8149_ (.RESET_B(net315),
    .D(_0211_),
    .Q(\led_controller.cpu.scratch_memory[2][3] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _8150_ (.RESET_B(net313),
    .D(_0212_),
    .Q(\led_controller.cpu.scratch_memory[2][4] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _8151_ (.RESET_B(net311),
    .D(_0213_),
    .Q(\led_controller.cpu.scratch_memory[2][5] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _8152_ (.RESET_B(net309),
    .D(_0214_),
    .Q(\led_controller.cpu.scratch_memory[2][6] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _8153_ (.RESET_B(net307),
    .D(_0215_),
    .Q(\led_controller.cpu.scratch_memory[2][7] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8154_ (.RESET_B(net305),
    .D(net1410),
    .Q(\led_controller.o_data ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _8155_ (.RESET_B(net303),
    .D(net2334),
    .Q(\led_controller.rgbw.pixel_counter[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _8156_ (.RESET_B(net301),
    .D(_0218_),
    .Q(\led_controller.rgbw.pixel_counter[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _8157_ (.RESET_B(net299),
    .D(_0219_),
    .Q(\led_controller.rgbw.pixel_counter[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _8158_ (.RESET_B(net297),
    .D(_0220_),
    .Q(\led_controller.rgbw.pixel_counter[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8159_ (.RESET_B(net295),
    .D(_0221_),
    .Q(\led_controller.rgbw.pixel_counter[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8160_ (.RESET_B(net293),
    .D(net1733),
    .Q(\led_controller.rgbw.pixel_counter[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8161_ (.RESET_B(net291),
    .D(_0223_),
    .Q(\led_controller.led_effect_pulse.color_1.active ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8162_ (.RESET_B(net290),
    .D(_0224_),
    .Q(\led_controller.rgbw.color[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8163_ (.RESET_B(net288),
    .D(_0225_),
    .Q(\led_controller.rgbw.color[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _8164_ (.RESET_B(net286),
    .D(_0226_),
    .Q(\led_controller.rgbw.color[2] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _8165_ (.RESET_B(net284),
    .D(_0227_),
    .Q(\led_controller.rgbw.color[3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _8166_ (.RESET_B(net282),
    .D(_0228_),
    .Q(\led_controller.rgbw.color[4] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _8167_ (.RESET_B(net280),
    .D(_0229_),
    .Q(\led_controller.rgbw.color[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8168_ (.RESET_B(net278),
    .D(_0230_),
    .Q(\led_controller.rgbw.color[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8169_ (.RESET_B(net276),
    .D(_0231_),
    .Q(\led_controller.rgbw.color[7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8170_ (.RESET_B(net274),
    .D(_0232_),
    .Q(\led_controller.rgbw.color[8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _8171_ (.RESET_B(net272),
    .D(_0233_),
    .Q(\led_controller.rgbw.color[9] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _8172_ (.RESET_B(net270),
    .D(_0234_),
    .Q(\led_controller.rgbw.color[10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8173_ (.RESET_B(net268),
    .D(_0235_),
    .Q(\led_controller.rgbw.color[11] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8174_ (.RESET_B(net266),
    .D(_0236_),
    .Q(\led_controller.rgbw.color[12] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8175_ (.RESET_B(net264),
    .D(_0237_),
    .Q(\led_controller.rgbw.color[13] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8176_ (.RESET_B(net262),
    .D(_0238_),
    .Q(\led_controller.rgbw.color[14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8177_ (.RESET_B(net260),
    .D(_0239_),
    .Q(\led_controller.rgbw.color[15] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _8178_ (.RESET_B(net258),
    .D(_0240_),
    .Q(\led_controller.rgbw.color[16] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8179_ (.RESET_B(net256),
    .D(_0241_),
    .Q(\led_controller.rgbw.color[17] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8180_ (.RESET_B(net254),
    .D(_0242_),
    .Q(\led_controller.rgbw.color[18] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8181_ (.RESET_B(net252),
    .D(_0243_),
    .Q(\led_controller.rgbw.color[19] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8182_ (.RESET_B(net250),
    .D(_0244_),
    .Q(\led_controller.rgbw.color[20] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8183_ (.RESET_B(net248),
    .D(_0245_),
    .Q(\led_controller.rgbw.color[21] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _8184_ (.RESET_B(net246),
    .D(_0246_),
    .Q(\led_controller.rgbw.color[22] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8185_ (.RESET_B(net244),
    .D(_0247_),
    .Q(\led_controller.rgbw.color[23] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _8186_ (.RESET_B(net242),
    .D(_0248_),
    .Q(\led_controller.rgbw.color[24] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8187_ (.RESET_B(net240),
    .D(_0249_),
    .Q(\led_controller.rgbw.color[25] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8188_ (.RESET_B(net238),
    .D(_0250_),
    .Q(\led_controller.rgbw.color[26] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8189_ (.RESET_B(net236),
    .D(_0251_),
    .Q(\led_controller.rgbw.color[27] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8190_ (.RESET_B(net234),
    .D(_0252_),
    .Q(\led_controller.rgbw.color[28] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _8191_ (.RESET_B(net232),
    .D(_0253_),
    .Q(\led_controller.rgbw.color[29] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _8192_ (.RESET_B(net230),
    .D(_0254_),
    .Q(\led_controller.rgbw.color[30] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _8193_ (.RESET_B(net228),
    .D(_0255_),
    .Q(\led_controller.rgbw.color[31] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _8194_ (.RESET_B(net226),
    .D(_0256_),
    .Q(\led_controller.rgbw.low_cycles[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _8195_ (.RESET_B(net224),
    .D(_0257_),
    .Q(\led_controller.rgbw.low_cycles[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _8196_ (.RESET_B(net222),
    .D(net2113),
    .Q(\led_controller.rgbw.low_cycles[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _8197_ (.RESET_B(net220),
    .D(net2029),
    .Q(\led_controller.rgbw.low_cycles[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _8198_ (.RESET_B(net218),
    .D(_0260_),
    .Q(\led_controller.rgbw.low_cycles[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _8199_ (.RESET_B(net216),
    .D(_0261_),
    .Q(\led_controller.rgbw.low_cycles[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _8200_ (.RESET_B(net214),
    .D(_0262_),
    .Q(\led_controller.rgbw.low_cycles[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _8201_ (.RESET_B(net212),
    .D(_0263_),
    .Q(\led_controller.rgbw.low_cycles[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _8202_ (.RESET_B(net210),
    .D(_0264_),
    .Q(\led_controller.rgbw.low_cycles[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _8203_ (.RESET_B(net208),
    .D(net1891),
    .Q(\led_controller.rgbw.low_cycles[9] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8204_ (.RESET_B(net206),
    .D(_0266_),
    .Q(\led_controller.rgbw.high_cycles[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _8205_ (.RESET_B(net204),
    .D(net2189),
    .Q(\led_controller.rgbw.high_cycles[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _8206_ (.RESET_B(net202),
    .D(net2110),
    .Q(\led_controller.rgbw.high_cycles[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _8207_ (.RESET_B(net200),
    .D(_0269_),
    .Q(\led_controller.flash.master.bit_counter[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8208_ (.RESET_B(net198),
    .D(net1524),
    .Q(\led_controller.flash.master.tx_data[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8209_ (.RESET_B(net196),
    .D(net1947),
    .Q(\led_controller.flash.master.tx_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8210_ (.RESET_B(net194),
    .D(net1611),
    .Q(\led_controller.flash.master.tx_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8211_ (.RESET_B(net192),
    .D(net1894),
    .Q(\led_controller.flash.master.tx_data[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8212_ (.RESET_B(net190),
    .D(_0274_),
    .Q(\led_controller.flash.master.tx_data[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8213_ (.RESET_B(net188),
    .D(net1586),
    .Q(\led_controller.flash.master.tx_data[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8214_ (.RESET_B(net186),
    .D(net1940),
    .Q(\led_controller.flash.master.tx_data[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8215_ (.RESET_B(net184),
    .D(_0277_),
    .Q(\led_controller.cpu.o_led_strb ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _8216_ (.RESET_B(net182),
    .D(net1479),
    .Q(\led_controller.cpu.o_led_color[0] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _8217_ (.RESET_B(net180),
    .D(net1436),
    .Q(\led_controller.cpu.o_led_color[1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _8218_ (.RESET_B(net178),
    .D(net1636),
    .Q(\led_controller.cpu.led_writing ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8219_ (.RESET_B(net176),
    .D(_0281_),
    .Q(\led_controller.cpu.led_write_pending ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8220_ (.RESET_B(net174),
    .D(_0282_),
    .Q(\led_controller.cpu.pc[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _8221_ (.RESET_B(net172),
    .D(_0283_),
    .Q(\led_controller.cpu.pc[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _8222_ (.RESET_B(net170),
    .D(_0284_),
    .Q(\led_controller.cpu.pc[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _8223_ (.RESET_B(net168),
    .D(_0285_),
    .Q(\led_controller.cpu.pc[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _8224_ (.RESET_B(net166),
    .D(net2323),
    .Q(\led_controller.cpu.pc[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _8225_ (.RESET_B(net164),
    .D(net2360),
    .Q(\led_controller.cpu.pc[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8226_ (.RESET_B(net162),
    .D(net2350),
    .Q(\led_controller.cpu.pc[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _8227_ (.RESET_B(net160),
    .D(_0289_),
    .Q(\led_controller.cpu.pc[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8228_ (.RESET_B(net158),
    .D(_0290_),
    .Q(\led_controller.cpu.pc[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8229_ (.RESET_B(net156),
    .D(_0291_),
    .Q(\led_controller.cpu.pc[9] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8230_ (.RESET_B(net154),
    .D(_0292_),
    .Q(\led_controller.cpu.pc[10] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _8231_ (.RESET_B(net152),
    .D(_0293_),
    .Q(\led_controller.cpu.pc[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _8232_ (.RESET_B(net150),
    .D(_0294_),
    .Q(\led_controller.cpu.pc[12] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8233_ (.RESET_B(net148),
    .D(_0295_),
    .Q(\led_controller.cpu.pc[13] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _8234_ (.RESET_B(net146),
    .D(_0296_),
    .Q(\led_controller.cpu.pc[14] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _8235_ (.RESET_B(net144),
    .D(_0297_),
    .Q(\led_controller.cpu.pc[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _8236_ (.RESET_B(net142),
    .D(_0298_),
    .Q(\led_controller.cpu.register_x[0] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _8237_ (.RESET_B(net140),
    .D(_0299_),
    .Q(\led_controller.cpu.register_x[1] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8238_ (.RESET_B(net138),
    .D(_0300_),
    .Q(\led_controller.cpu.register_x[2] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _8239_ (.RESET_B(net136),
    .D(_0301_),
    .Q(\led_controller.cpu.register_x[3] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _8240_ (.RESET_B(net134),
    .D(_0302_),
    .Q(\led_controller.cpu.register_x[4] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _8241_ (.RESET_B(net132),
    .D(_0303_),
    .Q(\led_controller.cpu.register_x[5] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _8242_ (.RESET_B(net130),
    .D(net2257),
    .Q(\led_controller.cpu.register_x[6] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8243_ (.RESET_B(net128),
    .D(net2338),
    .Q(\led_controller.cpu.register_x[7] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _8244_ (.RESET_B(net126),
    .D(_0306_),
    .Q(\led_controller.cpu.register_y[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8245_ (.RESET_B(net124),
    .D(_0307_),
    .Q(\led_controller.cpu.register_y[1] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8246_ (.RESET_B(net122),
    .D(_0308_),
    .Q(\led_controller.cpu.register_y[2] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8247_ (.RESET_B(net120),
    .D(_0309_),
    .Q(\led_controller.cpu.register_y[3] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _8248_ (.RESET_B(net118),
    .D(_0310_),
    .Q(\led_controller.cpu.register_y[4] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _8249_ (.RESET_B(net116),
    .D(_0311_),
    .Q(\led_controller.cpu.register_y[5] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _8250_ (.RESET_B(net114),
    .D(_0312_),
    .Q(\led_controller.cpu.register_y[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _8251_ (.RESET_B(net112),
    .D(_0313_),
    .Q(\led_controller.cpu.register_y[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _8252_ (.RESET_B(net110),
    .D(_0314_),
    .Q(\led_controller.cpu.status_zero ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _8253_ (.RESET_B(net108),
    .D(_0315_),
    .Q(\led_controller.cpu.status_negative ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _8254_ (.RESET_B(net106),
    .D(_0316_),
    .Q(\led_controller.cpu.stall_counter[0] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _8255_ (.RESET_B(net94),
    .D(_0317_),
    .Q(\led_controller.cpu.stall_counter[1] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _8256_ (.RESET_B(net92),
    .D(net2143),
    .Q(\led_controller.cpu.stall_counter[2] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _8257_ (.RESET_B(net90),
    .D(net1627),
    .Q(\led_controller.cpu.stall_counter[3] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _8258_ (.RESET_B(net88),
    .D(_0320_),
    .Q(\led_controller.cpu.stall_counter[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _8259_ (.RESET_B(net86),
    .D(_0321_),
    .Q(\led_controller.cpu.stall_counter[5] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _8260_ (.RESET_B(net84),
    .D(_0322_),
    .Q(\led_controller.cpu.stall_counter[6] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _8261_ (.RESET_B(net82),
    .D(net1532),
    .Q(\led_controller.cpu.stall_counter[7] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _8262_ (.RESET_B(net80),
    .D(_0324_),
    .Q(\led_controller.cpu.led_write_color[0] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _8263_ (.RESET_B(net78),
    .D(_0325_),
    .Q(\led_controller.cpu.led_write_color[1] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _8264_ (.RESET_B(net76),
    .D(_0326_),
    .Q(\led_controller.cpu.o_bus_addr[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _8265_ (.RESET_B(net74),
    .D(_0327_),
    .Q(\led_controller.cpu.o_bus_addr[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _8266_ (.RESET_B(net72),
    .D(net1729),
    .Q(\led_controller.cpu.o_bus_addr[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8267_ (.RESET_B(net67),
    .D(net2103),
    .Q(\led_controller.cpu.o_bus_addr[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _8268_ (.RESET_B(net65),
    .D(net1857),
    .Q(\led_controller.cpu.o_bus_addr[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _8269_ (.RESET_B(net63),
    .D(net1818),
    .Q(\led_controller.cpu.o_bus_addr[5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8270_ (.RESET_B(net61),
    .D(_0332_),
    .Q(\led_controller.cpu.o_bus_addr[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _8271_ (.RESET_B(net59),
    .D(_0333_),
    .Q(\led_controller.cpu.o_bus_addr[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8272_ (.RESET_B(net57),
    .D(_0334_),
    .Q(\led_controller.cpu.o_bus_addr[8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _8273_ (.RESET_B(net55),
    .D(_0335_),
    .Q(\led_controller.cpu.o_bus_addr[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8274_ (.RESET_B(net53),
    .D(net1603),
    .Q(\led_controller.cpu.o_bus_addr[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8275_ (.RESET_B(net51),
    .D(net2191),
    .Q(\led_controller.cpu.o_bus_addr[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8276_ (.RESET_B(net49),
    .D(_0338_),
    .Q(\led_controller.cpu.o_bus_addr[12] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _8277_ (.RESET_B(net47),
    .D(net1539),
    .Q(\led_controller.cpu.o_bus_addr[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8278_ (.RESET_B(net45),
    .D(net2219),
    .Q(\led_controller.cpu.o_bus_addr[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8279_ (.RESET_B(net43),
    .D(net1623),
    .Q(\led_controller.cpu.o_bus_addr[15] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8280_ (.RESET_B(net41),
    .D(net2316),
    .Q(\led_controller.cpu.o_bus_addr_valid ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _8281_ (.RESET_B(net39),
    .D(net1574),
    .Q(\led_controller.cpu.fetch_instruction[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _8282_ (.RESET_B(net37),
    .D(net1454),
    .Q(\led_controller.cpu.fetch_instruction[9] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _8283_ (.RESET_B(net35),
    .D(net1460),
    .Q(\led_controller.cpu.fetch_instruction[10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _8284_ (.RESET_B(net33),
    .D(net1441),
    .Q(\led_controller.cpu.fetch_instruction[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _8285_ (.RESET_B(net31),
    .D(net1542),
    .Q(\led_controller.cpu.fetch_instruction[12] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _8286_ (.RESET_B(net29),
    .D(net1374),
    .Q(\led_controller.cpu.fetch_instruction[13] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _8287_ (.RESET_B(net27),
    .D(net1417),
    .Q(\led_controller.cpu.fetch_instruction[14] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _8288_ (.RESET_B(net25),
    .D(net1419),
    .Q(\led_controller.cpu.fetch_instruction[15] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _8289_ (.RESET_B(net757),
    .D(_0351_),
    .Q(\led_controller.cpu.current_instruction[0] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _8290_ (.RESET_B(net755),
    .D(_0352_),
    .Q(\led_controller.cpu.current_instruction[1] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8291_ (.RESET_B(net753),
    .D(_0353_),
    .Q(\led_controller.cpu.current_instruction[2] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8292_ (.RESET_B(net751),
    .D(_0354_),
    .Q(\led_controller.cpu.current_instruction[3] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _8293_ (.RESET_B(net749),
    .D(net1625),
    .Q(\led_controller.cpu.current_instruction[4] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _8294_ (.RESET_B(net747),
    .D(net1598),
    .Q(\led_controller.cpu.current_instruction[5] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _8295_ (.RESET_B(net745),
    .D(net1444),
    .Q(\led_controller.cpu.current_instruction[6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _8296_ (.RESET_B(net743),
    .D(net1508),
    .Q(\led_controller.cpu.current_instruction[7] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _8297_ (.RESET_B(net741),
    .D(_0359_),
    .Q(\led_controller.cpu.current_instruction[8] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _8298_ (.RESET_B(net739),
    .D(_0360_),
    .Q(\led_controller.cpu.current_instruction[9] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _8299_ (.RESET_B(net737),
    .D(_0361_),
    .Q(\led_controller.cpu.current_instruction[10] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _8300_ (.RESET_B(net736),
    .D(_0362_),
    .Q(\led_controller.cpu.current_instruction[11] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _8301_ (.RESET_B(net734),
    .D(_0363_),
    .Q(\led_controller.cpu.current_instruction[12] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _8302_ (.RESET_B(net732),
    .D(net1340),
    .Q(\led_controller.cpu.current_instruction[13] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _8303_ (.RESET_B(net730),
    .D(net1360),
    .Q(\led_controller.cpu.current_instruction[14] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _8304_ (.RESET_B(net728),
    .D(net1346),
    .Q(\led_controller.cpu.current_instruction[15] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _8305_ (.RESET_B(net726),
    .D(net1552),
    .Q(\led_controller.cpu.current_instruction_pc[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _8306_ (.RESET_B(net724),
    .D(net1652),
    .Q(\led_controller.cpu.current_instruction_pc[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _8307_ (.RESET_B(net722),
    .D(net1484),
    .Q(\led_controller.cpu.current_instruction_pc[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _8308_ (.RESET_B(net720),
    .D(net1452),
    .Q(\led_controller.cpu.current_instruction_pc[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _8309_ (.RESET_B(net718),
    .D(net1562),
    .Q(\led_controller.cpu.current_instruction_pc[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _8310_ (.RESET_B(net716),
    .D(net1497),
    .Q(\led_controller.cpu.current_instruction_pc[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8311_ (.RESET_B(net714),
    .D(net1554),
    .Q(\led_controller.cpu.current_instruction_pc[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _8312_ (.RESET_B(net712),
    .D(_0374_),
    .Q(\led_controller.cpu.current_instruction_pc[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _8313_ (.RESET_B(net710),
    .D(net1506),
    .Q(\led_controller.cpu.current_instruction_pc[8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _8314_ (.RESET_B(net708),
    .D(net1504),
    .Q(\led_controller.cpu.current_instruction_pc[9] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8315_ (.RESET_B(net706),
    .D(net1462),
    .Q(\led_controller.cpu.current_instruction_pc[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8316_ (.RESET_B(net704),
    .D(net1518),
    .Q(\led_controller.cpu.current_instruction_pc[11] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8317_ (.RESET_B(net702),
    .D(net1477),
    .Q(\led_controller.cpu.current_instruction_pc[12] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8318_ (.RESET_B(net700),
    .D(net1450),
    .Q(\led_controller.cpu.current_instruction_pc[13] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8319_ (.RESET_B(net698),
    .D(net1486),
    .Q(\led_controller.cpu.current_instruction_pc[14] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _8320_ (.RESET_B(net696),
    .D(net1446),
    .Q(\led_controller.cpu.current_instruction_pc[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _8321_ (.RESET_B(net694),
    .D(_0383_),
    .Q(\led_controller.cpu.current_instruction_valid ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _8322_ (.RESET_B(net692),
    .D(_0384_),
    .Q(\led_controller.cpu.bus_hi_valid ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _8323_ (.RESET_B(net690),
    .D(_0385_),
    .Q(\led_controller.cpu.fetch_pc_valid ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _8324_ (.RESET_B(net688),
    .D(net1973),
    .Q(\led_controller.cpu.fetch_pc[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _8325_ (.RESET_B(net686),
    .D(_0387_),
    .Q(\led_controller.cpu.led_write_strb ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _8326_ (.RESET_B(net685),
    .D(net1943),
    .Q(\led_controller.flash.o_cs_n ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8327_ (.RESET_B(net683),
    .D(net1438),
    .Q(\led_controller.flash.addr[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8328_ (.RESET_B(net681),
    .D(net1401),
    .Q(\led_controller.flash.addr[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8329_ (.RESET_B(net679),
    .D(net1475),
    .Q(\led_controller.flash.addr[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8330_ (.RESET_B(net677),
    .D(net1493),
    .Q(\led_controller.flash.addr[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8331_ (.RESET_B(net675),
    .D(net1431),
    .Q(\led_controller.flash.addr[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8332_ (.RESET_B(net673),
    .D(net1383),
    .Q(\led_controller.flash.addr[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8333_ (.RESET_B(net671),
    .D(net1399),
    .Q(\led_controller.flash.addr[6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8334_ (.RESET_B(net669),
    .D(net1371),
    .Q(\led_controller.flash.addr[7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8335_ (.RESET_B(net667),
    .D(net1344),
    .Q(\led_controller.flash.addr[8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8336_ (.RESET_B(net665),
    .D(net1385),
    .Q(\led_controller.flash.addr[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8337_ (.RESET_B(net663),
    .D(net1379),
    .Q(\led_controller.flash.addr[10] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8338_ (.RESET_B(net661),
    .D(net1326),
    .Q(\led_controller.flash.addr[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8339_ (.RESET_B(net659),
    .D(net1330),
    .Q(\led_controller.flash.addr[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8340_ (.RESET_B(net657),
    .D(net1357),
    .Q(\led_controller.flash.addr[13] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8341_ (.RESET_B(net655),
    .D(net1322),
    .Q(\led_controller.flash.addr[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8342_ (.RESET_B(net653),
    .D(net1390),
    .Q(\led_controller.flash.addr[15] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _8343_ (.RESET_B(net651),
    .D(_0405_),
    .Q(\led_controller.flash.master.i_tx_data[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _8344_ (.RESET_B(net649),
    .D(_0406_),
    .Q(\led_controller.flash.master.i_tx_data[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _8345_ (.RESET_B(net642),
    .D(_0407_),
    .Q(\led_controller.flash.master.i_tx_data[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _8346_ (.RESET_B(net638),
    .D(_0408_),
    .Q(\led_controller.flash.master.i_tx_data[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _8347_ (.RESET_B(net634),
    .D(_0409_),
    .Q(\led_controller.flash.master.i_tx_data[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _8348_ (.RESET_B(net630),
    .D(_0410_),
    .Q(\led_controller.flash.master.i_tx_data[5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _8349_ (.RESET_B(net626),
    .D(_0411_),
    .Q(\led_controller.flash.master.i_tx_data[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8350_ (.RESET_B(net622),
    .D(_0412_),
    .Q(\led_controller.flash.master.i_tx_data[7] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _8351_ (.RESET_B(net618),
    .D(net1354),
    .Q(\led_controller.cpu.i_bus_data_valid ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8352_ (.RESET_B(net616),
    .D(net1805),
    .Q(\led_controller.flash.master.bit_counter[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _8353_ (.RESET_B(net612),
    .D(_0415_),
    .Q(\led_controller.flash.master.bit_counter[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8354_ (.RESET_B(net608),
    .D(net1685),
    .Q(\led_controller.flash.master.bit_counter[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _8355_ (.RESET_B(net604),
    .D(net1565),
    .Q(\led_controller.flash.master.sck_counter[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _8356_ (.RESET_B(net600),
    .D(_0418_),
    .Q(\led_controller.flash.master.sck_counter[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _8357_ (.RESET_B(net596),
    .D(net1527),
    .Q(\led_controller.flash.master.sck_counter[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _8358_ (.RESET_B(net590),
    .D(_0420_),
    .Q(\led_controller.flash.master.sck_counter[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _8359_ (.RESET_B(net586),
    .D(_0421_),
    .Q(\led_controller.flash.master.sck_counter[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _8360_ (.RESET_B(net582),
    .D(net1521),
    .Q(\led_controller.flash.master.sck_counter[5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8361_ (.RESET_B(net578),
    .D(_0423_),
    .Q(\led_controller.flash.master.sck_counter[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8362_ (.RESET_B(net574),
    .D(_0424_),
    .Q(\led_controller.flash.master.sck_counter[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _8363_ (.RESET_B(net570),
    .D(net1609),
    .Q(\led_controller.flash.master.active ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _8364_ (.RESET_B(net566),
    .D(_0426_),
    .Q(\led_controller.flash.master.o_busy ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _8365_ (.RESET_B(net564),
    .D(_0427_),
    .Q(\led_controller.cpu.i_bus_data[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _8366_ (.RESET_B(net552),
    .D(net1707),
    .Q(\led_controller.cpu.i_bus_data[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _8367_ (.RESET_B(net548),
    .D(_0429_),
    .Q(\led_controller.cpu.i_bus_data[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _8368_ (.RESET_B(net544),
    .D(net1629),
    .Q(\led_controller.cpu.i_bus_data[3] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _8369_ (.RESET_B(net540),
    .D(_0431_),
    .Q(\led_controller.cpu.i_bus_data[4] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _8370_ (.RESET_B(net536),
    .D(_0432_),
    .Q(\led_controller.cpu.i_bus_data[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _8371_ (.RESET_B(net532),
    .D(net1735),
    .Q(\led_controller.cpu.i_bus_data[6] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _8372_ (.RESET_B(net528),
    .D(_0434_),
    .Q(\led_controller.cpu.i_bus_data[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _8373_ (.RESET_B(net525),
    .D(_0435_),
    .Q(\led_controller.flash.master.sck ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _8374_ (.RESET_B(net521),
    .D(net765),
    .Q(\led_controller.flash.cs_delay_counter[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8375_ (.RESET_B(net519),
    .D(net2344),
    .Q(\led_controller.flash.cs_delay_counter[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8376_ (.RESET_B(net517),
    .D(net1557),
    .Q(\led_controller.flash.cs_delay_counter[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _8377_ (.RESET_B(net515),
    .D(_0439_),
    .Q(\led_controller.flash.cs_delay_counter[3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8378_ (.RESET_B(net513),
    .D(_0440_),
    .Q(\led_controller.flash.cs_delay_counter[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _8379_ (.RESET_B(net511),
    .D(net1720),
    .Q(\led_controller.flash.cs_delay_counter[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _8380_ (.RESET_B(net509),
    .D(net1607),
    .Q(\led_controller.flash.cs_delay_counter[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _8381_ (.RESET_B(net507),
    .D(net1567),
    .Q(\led_controller.flash.cs_delay_counter[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8382_ (.RESET_B(net505),
    .D(net1266),
    .Q(\led_controller.flash.master.o_mosi ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _8383_ (.RESET_B(net501),
    .D(_0445_),
    .Q(\led_controller.flash.master.tx_data[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _8384_ (.RESET_B(net497),
    .D(_0446_),
    .Q(\led_controller.cpu.scratch_memory[13][0] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _8385_ (.RESET_B(net493),
    .D(net1296),
    .Q(\led_controller.cpu.scratch_memory[13][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8386_ (.RESET_B(net489),
    .D(_0448_),
    .Q(\led_controller.cpu.scratch_memory[13][2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8387_ (.RESET_B(net485),
    .D(_0449_),
    .Q(\led_controller.cpu.scratch_memory[13][3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _8388_ (.RESET_B(net481),
    .D(_0450_),
    .Q(\led_controller.cpu.scratch_memory[13][4] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _8389_ (.RESET_B(net477),
    .D(_0451_),
    .Q(\led_controller.cpu.scratch_memory[13][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8390_ (.RESET_B(net473),
    .D(_0452_),
    .Q(\led_controller.cpu.scratch_memory[13][6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8391_ (.RESET_B(net469),
    .D(_0453_),
    .Q(\led_controller.cpu.scratch_memory[13][7] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _8392_ (.RESET_B(net465),
    .D(net1601),
    .Q(\led_controller.effect_chase_led_strb ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8393_ (.RESET_B(net461),
    .D(_0455_),
    .Q(\led_controller.effect_chase_led_color[0] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _8394_ (.RESET_B(net457),
    .D(net2291),
    .Q(\led_controller.effect_chase_led_color[1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _8395_ (.RESET_B(net453),
    .D(net1334),
    .Q(\led_controller.flash.master.o_rx_data_valid ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _8396_ (.RESET_B(net451),
    .D(_0458_),
    .Q(\led_controller.led_effect_chase.current_led[0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _8397_ (.RESET_B(net447),
    .D(net2331),
    .Q(\led_controller.led_effect_chase.current_led[1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _8398_ (.RESET_B(net406),
    .D(_0460_),
    .Q(\led_controller.led_effect_chase.current_led[2] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _8399_ (.RESET_B(net402),
    .D(_0461_),
    .Q(\led_controller.led_effect_chase.current_led[3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _8400_ (.RESET_B(net398),
    .D(_0462_),
    .Q(\led_controller.led_effect_chase.current_led[4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _8401_ (.RESET_B(net394),
    .D(net2116),
    .Q(\led_controller.led_effect_chase.current_led[5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _8402_ (.RESET_B(net390),
    .D(net1545),
    .Q(\led_controller.led_effect_chase.current_led[6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _8403_ (.RESET_B(net385),
    .D(net1654),
    .Q(\led_controller.led_effect_chase.current_led[7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _8404_ (.RESET_B(net381),
    .D(_0466_),
    .Q(\led_controller.cpu.scratch_memory[15][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _8405_ (.RESET_B(net377),
    .D(_0467_),
    .Q(\led_controller.cpu.scratch_memory[15][1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _8406_ (.RESET_B(net373),
    .D(_0468_),
    .Q(\led_controller.cpu.scratch_memory[15][2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _8407_ (.RESET_B(net369),
    .D(net1572),
    .Q(\led_controller.cpu.scratch_memory[15][3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _8408_ (.RESET_B(net365),
    .D(_0470_),
    .Q(\led_controller.cpu.scratch_memory[15][4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _8409_ (.RESET_B(net361),
    .D(_0471_),
    .Q(\led_controller.cpu.scratch_memory[15][5] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8410_ (.RESET_B(net357),
    .D(_0472_),
    .Q(\led_controller.cpu.scratch_memory[15][6] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _8411_ (.RESET_B(net353),
    .D(_0473_),
    .Q(\led_controller.cpu.scratch_memory[15][7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _8412_ (.RESET_B(net349),
    .D(_0474_),
    .Q(\led_controller.cpu.scratch_memory[7][0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8413_ (.RESET_B(net345),
    .D(_0475_),
    .Q(\led_controller.cpu.scratch_memory[7][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _8414_ (.RESET_B(net341),
    .D(_0476_),
    .Q(\led_controller.cpu.scratch_memory[7][2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _8415_ (.RESET_B(net337),
    .D(_0477_),
    .Q(\led_controller.cpu.scratch_memory[7][3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _8416_ (.RESET_B(net333),
    .D(_0478_),
    .Q(\led_controller.cpu.scratch_memory[7][4] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8417_ (.RESET_B(net329),
    .D(_0479_),
    .Q(\led_controller.cpu.scratch_memory[7][5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8418_ (.RESET_B(net325),
    .D(net809),
    .Q(\led_controller.cpu.scratch_memory[7][6] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8419_ (.RESET_B(net320),
    .D(_0481_),
    .Q(\led_controller.cpu.scratch_memory[7][7] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _8420_ (.RESET_B(net316),
    .D(net1846),
    .Q(\led_controller.effect_pulse_led_strb ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _8421_ (.RESET_B(net312),
    .D(net1427),
    .Q(\led_controller.effect_pulse_led_color[0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8422_ (.RESET_B(net308),
    .D(net1510),
    .Q(\led_controller.effect_pulse_led_color[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8423_ (.RESET_B(net304),
    .D(net1397),
    .Q(\led_controller.effect_pulse_led_color[2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _8424_ (.RESET_B(net300),
    .D(net1413),
    .Q(\led_controller.effect_pulse_led_color[3] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _8425_ (.RESET_B(net296),
    .D(net1423),
    .Q(\led_controller.effect_pulse_led_color[4] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8426_ (.RESET_B(net292),
    .D(net1425),
    .Q(\led_controller.effect_pulse_led_color[5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8427_ (.RESET_B(net287),
    .D(net1433),
    .Q(\led_controller.effect_pulse_led_color[6] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8428_ (.RESET_B(net283),
    .D(net1369),
    .Q(\led_controller.effect_pulse_led_color[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8429_ (.RESET_B(net279),
    .D(_0491_),
    .Q(\led_controller.effect_pulse_led_color[8] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8430_ (.RESET_B(net275),
    .D(net1421),
    .Q(\led_controller.effect_pulse_led_color[9] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _8431_ (.RESET_B(net271),
    .D(net1448),
    .Q(\led_controller.effect_pulse_led_color[10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8432_ (.RESET_B(net267),
    .D(_0494_),
    .Q(\led_controller.effect_pulse_led_color[11] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8433_ (.RESET_B(net263),
    .D(_0495_),
    .Q(\led_controller.effect_pulse_led_color[12] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8434_ (.RESET_B(net259),
    .D(_0496_),
    .Q(\led_controller.effect_pulse_led_color[13] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8435_ (.RESET_B(net255),
    .D(_0497_),
    .Q(\led_controller.effect_pulse_led_color[14] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8436_ (.RESET_B(net251),
    .D(_0498_),
    .Q(\led_controller.effect_pulse_led_color[15] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8437_ (.RESET_B(net247),
    .D(net1488),
    .Q(\led_controller.effect_pulse_led_color[16] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8438_ (.RESET_B(net243),
    .D(net1467),
    .Q(\led_controller.effect_pulse_led_color[17] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8439_ (.RESET_B(net239),
    .D(_0501_),
    .Q(\led_controller.effect_pulse_led_color[18] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8440_ (.RESET_B(net235),
    .D(net1469),
    .Q(\led_controller.effect_pulse_led_color[19] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _8441_ (.RESET_B(net231),
    .D(net1376),
    .Q(\led_controller.effect_pulse_led_color[20] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8442_ (.RESET_B(net227),
    .D(net1367),
    .Q(\led_controller.effect_pulse_led_color[21] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8443_ (.RESET_B(net223),
    .D(net1392),
    .Q(\led_controller.effect_pulse_led_color[22] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8444_ (.RESET_B(net219),
    .D(net1403),
    .Q(\led_controller.effect_pulse_led_color[23] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8445_ (.RESET_B(net215),
    .D(net1550),
    .Q(\led_controller.effect_pulse_led_color[24] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8446_ (.RESET_B(net211),
    .D(net1513),
    .Q(\led_controller.effect_pulse_led_color[25] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8447_ (.RESET_B(net207),
    .D(net1458),
    .Q(\led_controller.effect_pulse_led_color[26] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8448_ (.RESET_B(net203),
    .D(net1482),
    .Q(\led_controller.effect_pulse_led_color[27] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8449_ (.RESET_B(net199),
    .D(net1620),
    .Q(\led_controller.effect_pulse_led_color[28] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8450_ (.RESET_B(net195),
    .D(net1473),
    .Q(\led_controller.effect_pulse_led_color[29] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8451_ (.RESET_B(net191),
    .D(net1415),
    .Q(\led_controller.effect_pulse_led_color[30] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8452_ (.RESET_B(net187),
    .D(net1536),
    .Q(\led_controller.effect_pulse_led_color[31] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _8453_ (.RESET_B(net183),
    .D(net2239),
    .Q(\led_controller.led_effect_pulse.finished ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _8454_ (.RESET_B(net179),
    .D(_0516_),
    .Q(\led_controller.led_effect_pulse.current_led[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _8455_ (.RESET_B(net175),
    .D(net1777),
    .Q(\led_controller.led_effect_pulse.current_led[1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _8456_ (.RESET_B(net171),
    .D(_0518_),
    .Q(\led_controller.led_effect_pulse.current_led[2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8457_ (.RESET_B(net167),
    .D(net1594),
    .Q(\led_controller.led_effect_pulse.current_led[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _8458_ (.RESET_B(net163),
    .D(net1582),
    .Q(\led_controller.led_effect_pulse.current_led[4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _8459_ (.RESET_B(net159),
    .D(net2149),
    .Q(\led_controller.led_effect_pulse.current_led[5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _8460_ (.RESET_B(net155),
    .D(net1884),
    .Q(\led_controller.led_effect_pulse.current_led[6] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _8461_ (.RESET_B(net151),
    .D(net1739),
    .Q(\led_controller.led_effect_pulse.current_led[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _8462_ (.RESET_B(net147),
    .D(net1737),
    .Q(\led_controller.led_effect_pulse.color_index[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8463_ (.RESET_B(net143),
    .D(net2003),
    .Q(\led_controller.led_effect_pulse.color_index[1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8464_ (.RESET_B(net139),
    .D(_0526_),
    .Q(\led_controller.led_effect_pulse.brightness[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _8465_ (.RESET_B(net135),
    .D(_0527_),
    .Q(\led_controller.led_effect_pulse.brightness[1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _8466_ (.RESET_B(net131),
    .D(net2282),
    .Q(\led_controller.led_effect_pulse.brightness[2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _8467_ (.RESET_B(net127),
    .D(_0529_),
    .Q(\led_controller.led_effect_pulse.brightness[3] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _8468_ (.RESET_B(net123),
    .D(net2278),
    .Q(\led_controller.led_effect_pulse.brightness[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _8469_ (.RESET_B(net119),
    .D(net2230),
    .Q(\led_controller.led_effect_pulse.color_1.i_strb ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _8470_ (.RESET_B(net115),
    .D(_0532_),
    .Q(\led_controller.led_effect_pulse.calc_color_valid ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _8471_ (.RESET_B(net113),
    .D(_0533_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8472_ (.RESET_B(net111),
    .D(_0534_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8473_ (.RESET_B(net109),
    .D(net1881),
    .Q(\led_controller.led_effect_pulse.calc_color_out[2] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _8474_ (.RESET_B(net107),
    .D(_0536_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[3] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _8475_ (.RESET_B(net95),
    .D(_0537_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[4] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8476_ (.RESET_B(net93),
    .D(_0538_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[5] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8477_ (.RESET_B(net91),
    .D(_0539_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8478_ (.RESET_B(net89),
    .D(_0540_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[7] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8479_ (.RESET_B(net87),
    .D(_0541_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[8] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8480_ (.RESET_B(net85),
    .D(net1810),
    .Q(\led_controller.led_effect_pulse.calc_color_out[9] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _8481_ (.RESET_B(net83),
    .D(_0543_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8482_ (.RESET_B(net81),
    .D(_0544_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[11] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8483_ (.RESET_B(net79),
    .D(_0545_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[12] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8484_ (.RESET_B(net77),
    .D(_0546_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[13] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8485_ (.RESET_B(net75),
    .D(_0547_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[14] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8486_ (.RESET_B(net73),
    .D(_0548_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[15] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8487_ (.RESET_B(net68),
    .D(_0549_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[16] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8488_ (.RESET_B(net66),
    .D(_0550_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[17] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8489_ (.RESET_B(net64),
    .D(net1465),
    .Q(\led_controller.led_effect_pulse.calc_color_out[18] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8490_ (.RESET_B(net62),
    .D(_0552_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[19] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _8491_ (.RESET_B(net60),
    .D(_0553_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[20] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8492_ (.RESET_B(net58),
    .D(_0554_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[21] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8493_ (.RESET_B(net56),
    .D(_0555_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[22] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8494_ (.RESET_B(net54),
    .D(net1692),
    .Q(\led_controller.led_effect_pulse.calc_color_out[23] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8495_ (.RESET_B(net52),
    .D(_0557_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[24] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8496_ (.RESET_B(net50),
    .D(net1871),
    .Q(\led_controller.led_effect_pulse.calc_color_out[25] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8497_ (.RESET_B(net48),
    .D(_0559_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[26] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8498_ (.RESET_B(net46),
    .D(_0560_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[27] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8499_ (.RESET_B(net44),
    .D(net1932),
    .Q(\led_controller.led_effect_pulse.calc_color_out[28] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _8500_ (.RESET_B(net42),
    .D(_0562_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[29] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8501_ (.RESET_B(net40),
    .D(_0563_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[30] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8502_ (.RESET_B(net38),
    .D(_0564_),
    .Q(\led_controller.led_effect_pulse.calc_color_out[31] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _8503_ (.RESET_B(net36),
    .D(_0565_),
    .Q(\led_controller.led_effect_pulse.color_1.counter[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _8504_ (.RESET_B(net34),
    .D(_0566_),
    .Q(\led_controller.led_effect_pulse.color_1.counter[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _8505_ (.RESET_B(net32),
    .D(_0567_),
    .Q(\led_controller.led_effect_chase.finished ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _8506_ (.RESET_B(net30),
    .D(_0568_),
    .Q(\led_controller.cpu.fetch_instruction[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _8507_ (.RESET_B(net26),
    .D(_0569_),
    .Q(\led_controller.cpu.fetch_instruction[1] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _8508_ (.RESET_B(net756),
    .D(_0570_),
    .Q(\led_controller.cpu.fetch_instruction[2] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _8509_ (.RESET_B(net752),
    .D(_0571_),
    .Q(\led_controller.cpu.fetch_instruction[3] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _8510_ (.RESET_B(net748),
    .D(_0572_),
    .Q(\led_controller.cpu.fetch_instruction[4] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _8511_ (.RESET_B(net744),
    .D(_0573_),
    .Q(\led_controller.cpu.fetch_instruction[5] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _8512_ (.RESET_B(net740),
    .D(_0574_),
    .Q(\led_controller.cpu.fetch_instruction[6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _8513_ (.RESET_B(net594),
    .D(_0575_),
    .Q(\led_controller.cpu.fetch_instruction[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _8514_ (.RESET_B(net1),
    .D(net760),
    .Q(\led_controller.led_effect_chase.i_reset_n ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _8515_ (.RESET_B(net1),
    .D(net1),
    .Q(\led_controller.reset.reset1 ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _8516_ (.RESET_B(net733),
    .D(_0576_),
    .Q(\led_controller.cpu_reset_counter[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8517_ (.RESET_B(net731),
    .D(_0577_),
    .Q(\led_controller.cpu_reset_counter[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8518_ (.RESET_B(net729),
    .D(_0578_),
    .Q(\led_controller.cpu_reset_counter[2] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _8519_ (.RESET_B(net727),
    .D(_0579_),
    .Q(\led_controller.cpu_reset_counter[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8520_ (.RESET_B(net725),
    .D(_0580_),
    .Q(\led_controller.spi_data_write_strb ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8521_ (.RESET_B(net723),
    .D(net2309),
    .Q(\led_controller.flash.i_addr_width_24 ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _8522_ (.RESET_B(net719),
    .D(net1499),
    .Q(\led_controller.spi_data_write[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _8523_ (.RESET_B(net715),
    .D(_0583_),
    .Q(\led_controller.spi_data_write[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8524_ (.RESET_B(net711),
    .D(_0584_),
    .Q(\led_controller.spi_data_write[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _8525_ (.RESET_B(net707),
    .D(_0585_),
    .Q(\led_controller.spi_data_write[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8526_ (.RESET_B(net703),
    .D(_0586_),
    .Q(\led_controller.spi_data_write[4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _8527_ (.RESET_B(net699),
    .D(_0587_),
    .Q(\led_controller.spi_data_write[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8528_ (.RESET_B(net695),
    .D(_0588_),
    .Q(\led_controller.spi_data_write[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _8529_ (.RESET_B(net691),
    .D(_0589_),
    .Q(\led_controller.spi_data_write[7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8530_ (.RESET_B(net687),
    .D(_0590_),
    .Q(\led_controller.register_data[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8531_ (.RESET_B(net682),
    .D(_0591_),
    .Q(\led_controller.register_data[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8532_ (.RESET_B(net678),
    .D(_0592_),
    .Q(\led_controller.register_data[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8533_ (.RESET_B(net674),
    .D(_0593_),
    .Q(\led_controller.register_data[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8534_ (.RESET_B(net670),
    .D(_0594_),
    .Q(\led_controller.register_data[4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8535_ (.RESET_B(net666),
    .D(_0595_),
    .Q(\led_controller.register_data[5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _8536_ (.RESET_B(net662),
    .D(_0596_),
    .Q(\led_controller.register_data[6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8537_ (.RESET_B(net658),
    .D(_0597_),
    .Q(\led_controller.register_data[7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _8538_ (.RESET_B(net654),
    .D(_0598_),
    .Q(\led_controller.register_address[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _8539_ (.RESET_B(net650),
    .D(net1953),
    .Q(\led_controller.register_address[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _8540_ (.RESET_B(net640),
    .D(net1787),
    .Q(\led_controller.register_address[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8541_ (.RESET_B(net632),
    .D(net1799),
    .Q(\led_controller.register_address[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8542_ (.RESET_B(net624),
    .D(_0602_),
    .Q(\led_controller.register_address[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _8543_ (.RESET_B(net614),
    .D(_0603_),
    .Q(\led_controller.register_address[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _8544_ (.RESET_B(net606),
    .D(net1634),
    .Q(\led_controller.register_address[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _8545_ (.RESET_B(net598),
    .D(net2129),
    .Q(\led_controller.register_address[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _8546_ (.RESET_B(net588),
    .D(_0606_),
    .Q(\led_controller.cpu.i_num_colors[0] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8547_ (.RESET_B(net580),
    .D(_0607_),
    .Q(\led_controller.cpu.i_num_colors[1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8548_ (.RESET_B(net572),
    .D(net2263),
    .Q(\led_controller.colors[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8549_ (.RESET_B(net562),
    .D(net2125),
    .Q(\led_controller.colors[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8550_ (.RESET_B(net546),
    .D(net2123),
    .Q(\led_controller.colors[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8551_ (.RESET_B(net538),
    .D(net2001),
    .Q(\led_controller.colors[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8552_ (.RESET_B(net530),
    .D(_0612_),
    .Q(\led_controller.colors[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8553_ (.RESET_B(net523),
    .D(net1949),
    .Q(\led_controller.colors[5] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8554_ (.RESET_B(net499),
    .D(net2141),
    .Q(\led_controller.colors[6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8555_ (.RESET_B(net491),
    .D(_0615_),
    .Q(\led_controller.colors[7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _8556_ (.RESET_B(net483),
    .D(_0616_),
    .Q(\led_controller.colors[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _8557_ (.RESET_B(net475),
    .D(_0617_),
    .Q(\led_controller.colors[9] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8558_ (.RESET_B(net467),
    .D(_0618_),
    .Q(\led_controller.colors[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8559_ (.RESET_B(net459),
    .D(_0619_),
    .Q(\led_controller.colors[11] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8560_ (.RESET_B(net449),
    .D(_0620_),
    .Q(\led_controller.colors[12] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8561_ (.RESET_B(net404),
    .D(_0621_),
    .Q(\led_controller.colors[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8562_ (.RESET_B(net396),
    .D(_0622_),
    .Q(\led_controller.colors[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8563_ (.RESET_B(net388),
    .D(_0623_),
    .Q(\led_controller.colors[15] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8564_ (.RESET_B(net379),
    .D(_0624_),
    .Q(\led_controller.colors[16] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8565_ (.RESET_B(net371),
    .D(_0625_),
    .Q(\led_controller.colors[17] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8566_ (.RESET_B(net363),
    .D(_0626_),
    .Q(\led_controller.colors[18] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _8567_ (.RESET_B(net355),
    .D(_0627_),
    .Q(\led_controller.colors[19] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8568_ (.RESET_B(net347),
    .D(_0628_),
    .Q(\led_controller.colors[20] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8569_ (.RESET_B(net339),
    .D(_0629_),
    .Q(\led_controller.colors[21] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _8570_ (.RESET_B(net331),
    .D(_0630_),
    .Q(\led_controller.colors[22] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8571_ (.RESET_B(net323),
    .D(_0631_),
    .Q(\led_controller.colors[23] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8572_ (.RESET_B(net314),
    .D(_0632_),
    .Q(\led_controller.colors[24] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8573_ (.RESET_B(net306),
    .D(_0633_),
    .Q(\led_controller.colors[25] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8574_ (.RESET_B(net298),
    .D(_0634_),
    .Q(\led_controller.colors[26] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8575_ (.RESET_B(net289),
    .D(_0635_),
    .Q(\led_controller.colors[27] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8576_ (.RESET_B(net281),
    .D(_0636_),
    .Q(\led_controller.colors[28] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8577_ (.RESET_B(net273),
    .D(_0637_),
    .Q(\led_controller.colors[29] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8578_ (.RESET_B(net265),
    .D(_0638_),
    .Q(\led_controller.colors[30] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8579_ (.RESET_B(net257),
    .D(_0639_),
    .Q(\led_controller.colors[31] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8580_ (.RESET_B(net249),
    .D(_0640_),
    .Q(\led_controller.colors[32] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8581_ (.RESET_B(net241),
    .D(_0641_),
    .Q(\led_controller.colors[33] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8582_ (.RESET_B(net233),
    .D(_0642_),
    .Q(\led_controller.colors[34] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8583_ (.RESET_B(net225),
    .D(_0643_),
    .Q(\led_controller.colors[35] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8584_ (.RESET_B(net217),
    .D(_0644_),
    .Q(\led_controller.colors[36] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8585_ (.RESET_B(net209),
    .D(_0645_),
    .Q(\led_controller.colors[37] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8586_ (.RESET_B(net201),
    .D(_0646_),
    .Q(\led_controller.colors[38] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8587_ (.RESET_B(net193),
    .D(_0647_),
    .Q(\led_controller.colors[39] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8588_ (.RESET_B(net185),
    .D(_0648_),
    .Q(\led_controller.colors[40] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8589_ (.RESET_B(net177),
    .D(_0649_),
    .Q(\led_controller.colors[41] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8590_ (.RESET_B(net169),
    .D(_0650_),
    .Q(\led_controller.colors[42] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8591_ (.RESET_B(net161),
    .D(_0651_),
    .Q(\led_controller.colors[43] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8592_ (.RESET_B(net153),
    .D(_0652_),
    .Q(\led_controller.colors[44] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8593_ (.RESET_B(net145),
    .D(_0653_),
    .Q(\led_controller.colors[45] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8594_ (.RESET_B(net137),
    .D(_0654_),
    .Q(\led_controller.colors[46] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8595_ (.RESET_B(net129),
    .D(_0655_),
    .Q(\led_controller.colors[47] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8596_ (.RESET_B(net121),
    .D(_0656_),
    .Q(\led_controller.colors[48] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _8597_ (.RESET_B(net28),
    .D(_0657_),
    .Q(\led_controller.colors[49] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8598_ (.RESET_B(net754),
    .D(_0658_),
    .Q(\led_controller.colors[50] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8599_ (.RESET_B(net746),
    .D(_0659_),
    .Q(\led_controller.colors[51] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8600_ (.RESET_B(net738),
    .D(_0660_),
    .Q(\led_controller.colors[52] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _8601_ (.RESET_B(net721),
    .D(_0661_),
    .Q(\led_controller.colors[53] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8602_ (.RESET_B(net713),
    .D(_0662_),
    .Q(\led_controller.colors[54] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8603_ (.RESET_B(net705),
    .D(_0663_),
    .Q(\led_controller.colors[55] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8604_ (.RESET_B(net697),
    .D(_0664_),
    .Q(\led_controller.colors[56] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _8605_ (.RESET_B(net689),
    .D(_0665_),
    .Q(\led_controller.colors[57] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8606_ (.RESET_B(net680),
    .D(_0666_),
    .Q(\led_controller.colors[58] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8607_ (.RESET_B(net672),
    .D(_0667_),
    .Q(\led_controller.colors[59] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8608_ (.RESET_B(net664),
    .D(_0668_),
    .Q(\led_controller.colors[60] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8609_ (.RESET_B(net656),
    .D(_0669_),
    .Q(\led_controller.colors[61] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _8610_ (.RESET_B(net648),
    .D(_0670_),
    .Q(\led_controller.colors[62] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8611_ (.RESET_B(net628),
    .D(_0671_),
    .Q(\led_controller.colors[63] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8612_ (.RESET_B(net610),
    .D(_0672_),
    .Q(\led_controller.colors[64] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8613_ (.RESET_B(net592),
    .D(_0673_),
    .Q(\led_controller.colors[65] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8614_ (.RESET_B(net576),
    .D(_0674_),
    .Q(\led_controller.colors[66] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8615_ (.RESET_B(net550),
    .D(_0675_),
    .Q(\led_controller.colors[67] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8616_ (.RESET_B(net534),
    .D(_0676_),
    .Q(\led_controller.colors[68] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8617_ (.RESET_B(net503),
    .D(_0677_),
    .Q(\led_controller.colors[69] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8618_ (.RESET_B(net487),
    .D(_0678_),
    .Q(\led_controller.colors[70] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8619_ (.RESET_B(net471),
    .D(_0679_),
    .Q(\led_controller.colors[71] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8620_ (.RESET_B(net455),
    .D(_0680_),
    .Q(\led_controller.colors[72] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8621_ (.RESET_B(net400),
    .D(_0681_),
    .Q(\led_controller.colors[73] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8622_ (.RESET_B(net383),
    .D(_0682_),
    .Q(\led_controller.colors[74] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8623_ (.RESET_B(net367),
    .D(_0683_),
    .Q(\led_controller.colors[75] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8624_ (.RESET_B(net351),
    .D(_0684_),
    .Q(\led_controller.colors[76] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8625_ (.RESET_B(net335),
    .D(_0685_),
    .Q(\led_controller.colors[77] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _8626_ (.RESET_B(net318),
    .D(_0686_),
    .Q(\led_controller.colors[78] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8627_ (.RESET_B(net302),
    .D(_0687_),
    .Q(\led_controller.colors[79] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8628_ (.RESET_B(net285),
    .D(_0688_),
    .Q(\led_controller.colors[80] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _8629_ (.RESET_B(net269),
    .D(_0689_),
    .Q(\led_controller.colors[81] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8630_ (.RESET_B(net253),
    .D(_0690_),
    .Q(\led_controller.colors[82] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8631_ (.RESET_B(net237),
    .D(_0691_),
    .Q(\led_controller.colors[83] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8632_ (.RESET_B(net221),
    .D(_0692_),
    .Q(\led_controller.colors[84] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _8633_ (.RESET_B(net205),
    .D(_0693_),
    .Q(\led_controller.colors[85] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _8634_ (.RESET_B(net189),
    .D(_0694_),
    .Q(\led_controller.colors[86] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8635_ (.RESET_B(net173),
    .D(_0695_),
    .Q(\led_controller.colors[87] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8636_ (.RESET_B(net157),
    .D(_0696_),
    .Q(\led_controller.colors[88] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _8637_ (.RESET_B(net141),
    .D(_0697_),
    .Q(\led_controller.colors[89] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8638_ (.RESET_B(net125),
    .D(_0698_),
    .Q(\led_controller.colors[90] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _8639_ (.RESET_B(net758),
    .D(_0699_),
    .Q(\led_controller.colors[91] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8640_ (.RESET_B(net742),
    .D(_0700_),
    .Q(\led_controller.colors[92] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _8641_ (.RESET_B(net717),
    .D(_0701_),
    .Q(\led_controller.colors[93] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8642_ (.RESET_B(net701),
    .D(_0702_),
    .Q(\led_controller.colors[94] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _8643_ (.RESET_B(net684),
    .D(_0703_),
    .Q(\led_controller.colors[95] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _8644_ (.RESET_B(net668),
    .D(_0704_),
    .Q(\led_controller.cpu.i_num_leds[0] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8645_ (.RESET_B(net652),
    .D(net2253),
    .Q(\led_controller.cpu.i_num_leds[1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8646_ (.RESET_B(net620),
    .D(net2301),
    .Q(\led_controller.cpu.i_num_leds[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8647_ (.RESET_B(net584),
    .D(net2209),
    .Q(\led_controller.cpu.i_num_leds[3] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8648_ (.RESET_B(net542),
    .D(net2202),
    .Q(\led_controller.cpu.i_num_leds[4] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8649_ (.RESET_B(net495),
    .D(_0709_),
    .Q(\led_controller.cpu.i_num_leds[5] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8650_ (.RESET_B(net463),
    .D(_0710_),
    .Q(\led_controller.cpu.i_num_leds[6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8651_ (.RESET_B(net392),
    .D(net2043),
    .Q(\led_controller.cpu.i_num_leds[7] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8652_ (.RESET_B(net359),
    .D(net2163),
    .Q(\led_controller.effect[0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8653_ (.RESET_B(net327),
    .D(_0713_),
    .Q(\led_controller.effect[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8654_ (.RESET_B(net294),
    .D(_0714_),
    .Q(\led_controller.effect[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8655_ (.RESET_B(net261),
    .D(_0715_),
    .Q(\led_controller.effect[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8656_ (.RESET_B(net229),
    .D(_0716_),
    .Q(\led_controller.clock_divider[0] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8657_ (.RESET_B(net197),
    .D(_0717_),
    .Q(\led_controller.clock_divider[1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8658_ (.RESET_B(net165),
    .D(_0718_),
    .Q(\led_controller.clock_divider[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _8659_ (.RESET_B(net133),
    .D(_0719_),
    .Q(\led_controller.clock_divider[3] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8660_ (.RESET_B(net750),
    .D(_0720_),
    .Q(\led_controller.clock_divider[4] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8661_ (.RESET_B(net709),
    .D(_0721_),
    .Q(\led_controller.clock_divider[5] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8662_ (.RESET_B(net676),
    .D(_0722_),
    .Q(\led_controller.clock_divider[6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8663_ (.RESET_B(net636),
    .D(_0723_),
    .Q(\led_controller.clock_divider[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _8664_ (.RESET_B(net568),
    .D(_0724_),
    .Q(\led_controller.cpu.scratch_memory[0][0] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _8665_ (.RESET_B(net479),
    .D(_0725_),
    .Q(\led_controller.cpu.scratch_memory[0][1] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8666_ (.RESET_B(net375),
    .D(_0726_),
    .Q(\led_controller.cpu.scratch_memory[0][2] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _8667_ (.RESET_B(net310),
    .D(_0727_),
    .Q(\led_controller.cpu.scratch_memory[0][3] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8668_ (.RESET_B(net245),
    .D(_0728_),
    .Q(\led_controller.cpu.scratch_memory[0][4] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8669_ (.RESET_B(net181),
    .D(_0729_),
    .Q(\led_controller.cpu.scratch_memory[0][5] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8670_ (.RESET_B(net117),
    .D(_0730_),
    .Q(\led_controller.cpu.scratch_memory[0][6] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8671_ (.RESET_B(net693),
    .D(_0731_),
    .Q(\led_controller.cpu.scratch_memory[0][7] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8672_ (.RESET_B(net602),
    .D(net1304),
    .Q(\led_controller.cpu.scratch_memory[8][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _8673_ (.RESET_B(net445),
    .D(net1244),
    .Q(\led_controller.cpu.scratch_memory[8][1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _8674_ (.RESET_B(net277),
    .D(net1269),
    .Q(\led_controller.cpu.scratch_memory[8][2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _8675_ (.RESET_B(net149),
    .D(net1278),
    .Q(\led_controller.cpu.scratch_memory[8][3] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8676_ (.RESET_B(net660),
    .D(net1259),
    .Q(\led_controller.cpu.scratch_memory[8][4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8677_ (.RESET_B(net343),
    .D(net1257),
    .Q(\led_controller.cpu.scratch_memory[8][5] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _8678_ (.RESET_B(net735),
    .D(net1316),
    .Q(\led_controller.cpu.scratch_memory[8][6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _8679_ (.RESET_B(net213),
    .D(net1232),
    .Q(\led_controller.cpu.scratch_memory[8][7] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_tiehi _8288__25 (.L_HI(net25));
 sg13g2_tiehi _8507__26 (.L_HI(net26));
 sg13g2_tiehi _8287__27 (.L_HI(net27));
 sg13g2_tiehi _8597__28 (.L_HI(net28));
 sg13g2_tiehi _8286__29 (.L_HI(net29));
 sg13g2_tiehi _8506__30 (.L_HI(net30));
 sg13g2_tiehi _8285__31 (.L_HI(net31));
 sg13g2_tiehi _8505__32 (.L_HI(net32));
 sg13g2_tiehi _8284__33 (.L_HI(net33));
 sg13g2_tiehi _8504__34 (.L_HI(net34));
 sg13g2_tiehi _8283__35 (.L_HI(net35));
 sg13g2_tiehi _8503__36 (.L_HI(net36));
 sg13g2_tiehi _8282__37 (.L_HI(net37));
 sg13g2_tiehi _8502__38 (.L_HI(net38));
 sg13g2_tiehi _8281__39 (.L_HI(net39));
 sg13g2_tiehi _8501__40 (.L_HI(net40));
 sg13g2_tiehi _8280__41 (.L_HI(net41));
 sg13g2_tiehi _8500__42 (.L_HI(net42));
 sg13g2_tiehi _8279__43 (.L_HI(net43));
 sg13g2_tiehi _8499__44 (.L_HI(net44));
 sg13g2_tiehi _8278__45 (.L_HI(net45));
 sg13g2_tiehi _8498__46 (.L_HI(net46));
 sg13g2_tiehi _8277__47 (.L_HI(net47));
 sg13g2_tiehi _8497__48 (.L_HI(net48));
 sg13g2_tiehi _8276__49 (.L_HI(net49));
 sg13g2_tiehi _8496__50 (.L_HI(net50));
 sg13g2_tiehi _8275__51 (.L_HI(net51));
 sg13g2_tiehi _8495__52 (.L_HI(net52));
 sg13g2_tiehi _8274__53 (.L_HI(net53));
 sg13g2_tiehi _8494__54 (.L_HI(net54));
 sg13g2_tiehi _8273__55 (.L_HI(net55));
 sg13g2_tiehi _8493__56 (.L_HI(net56));
 sg13g2_tiehi _8272__57 (.L_HI(net57));
 sg13g2_tiehi _8492__58 (.L_HI(net58));
 sg13g2_tiehi _8271__59 (.L_HI(net59));
 sg13g2_tiehi _8491__60 (.L_HI(net60));
 sg13g2_tiehi _8270__61 (.L_HI(net61));
 sg13g2_tiehi _8490__62 (.L_HI(net62));
 sg13g2_tiehi _8269__63 (.L_HI(net63));
 sg13g2_tiehi _8489__64 (.L_HI(net64));
 sg13g2_tiehi _8268__65 (.L_HI(net65));
 sg13g2_tiehi _8488__66 (.L_HI(net66));
 sg13g2_tiehi _8267__67 (.L_HI(net67));
 sg13g2_tiehi _8487__68 (.L_HI(net68));
 sg13g2_tiehi _7943__69 (.L_HI(net69));
 sg13g2_tiehi _7988__70 (.L_HI(net70));
 sg13g2_tiehi _7989__71 (.L_HI(net71));
 sg13g2_tiehi _8266__72 (.L_HI(net72));
 sg13g2_tiehi _8486__73 (.L_HI(net73));
 sg13g2_tiehi _8265__74 (.L_HI(net74));
 sg13g2_tiehi _8485__75 (.L_HI(net75));
 sg13g2_tiehi _8264__76 (.L_HI(net76));
 sg13g2_tiehi _8484__77 (.L_HI(net77));
 sg13g2_tiehi _8263__78 (.L_HI(net78));
 sg13g2_tiehi _8483__79 (.L_HI(net79));
 sg13g2_tiehi _8262__80 (.L_HI(net80));
 sg13g2_tiehi _8482__81 (.L_HI(net81));
 sg13g2_tiehi _8261__82 (.L_HI(net82));
 sg13g2_tiehi _8481__83 (.L_HI(net83));
 sg13g2_tiehi _8260__84 (.L_HI(net84));
 sg13g2_tiehi _8480__85 (.L_HI(net85));
 sg13g2_tiehi _8259__86 (.L_HI(net86));
 sg13g2_tiehi _8479__87 (.L_HI(net87));
 sg13g2_tiehi _8258__88 (.L_HI(net88));
 sg13g2_tiehi _8478__89 (.L_HI(net89));
 sg13g2_tiehi _8257__90 (.L_HI(net90));
 sg13g2_tiehi _8477__91 (.L_HI(net91));
 sg13g2_tiehi _8256__92 (.L_HI(net92));
 sg13g2_tiehi _8476__93 (.L_HI(net93));
 sg13g2_tiehi _8255__94 (.L_HI(net94));
 sg13g2_tiehi _8475__95 (.L_HI(net95));
 sg13g2_tiehi _7990__96 (.L_HI(net96));
 sg13g2_tiehi _8015__97 (.L_HI(net97));
 sg13g2_tiehi _8016__98 (.L_HI(net98));
 sg13g2_tiehi _8017__99 (.L_HI(net99));
 sg13g2_tiehi _8018__100 (.L_HI(net100));
 sg13g2_tiehi _8019__101 (.L_HI(net101));
 sg13g2_tiehi _8020__102 (.L_HI(net102));
 sg13g2_tiehi _8021__103 (.L_HI(net103));
 sg13g2_tiehi _8022__104 (.L_HI(net104));
 sg13g2_tiehi _8023__105 (.L_HI(net105));
 sg13g2_tiehi _8254__106 (.L_HI(net106));
 sg13g2_tiehi _8474__107 (.L_HI(net107));
 sg13g2_tiehi _8253__108 (.L_HI(net108));
 sg13g2_tiehi _8473__109 (.L_HI(net109));
 sg13g2_tiehi _8252__110 (.L_HI(net110));
 sg13g2_tiehi _8472__111 (.L_HI(net111));
 sg13g2_tiehi _8251__112 (.L_HI(net112));
 sg13g2_tiehi _8471__113 (.L_HI(net113));
 sg13g2_tiehi _8250__114 (.L_HI(net114));
 sg13g2_tiehi _8470__115 (.L_HI(net115));
 sg13g2_tiehi _8249__116 (.L_HI(net116));
 sg13g2_tiehi _8670__117 (.L_HI(net117));
 sg13g2_tiehi _8248__118 (.L_HI(net118));
 sg13g2_tiehi _8469__119 (.L_HI(net119));
 sg13g2_tiehi _8247__120 (.L_HI(net120));
 sg13g2_tiehi _8596__121 (.L_HI(net121));
 sg13g2_tiehi _8246__122 (.L_HI(net122));
 sg13g2_tiehi _8468__123 (.L_HI(net123));
 sg13g2_tiehi _8245__124 (.L_HI(net124));
 sg13g2_tiehi _8638__125 (.L_HI(net125));
 sg13g2_tiehi _8244__126 (.L_HI(net126));
 sg13g2_tiehi _8467__127 (.L_HI(net127));
 sg13g2_tiehi _8243__128 (.L_HI(net128));
 sg13g2_tiehi _8595__129 (.L_HI(net129));
 sg13g2_tiehi _8242__130 (.L_HI(net130));
 sg13g2_tiehi _8466__131 (.L_HI(net131));
 sg13g2_tiehi _8241__132 (.L_HI(net132));
 sg13g2_tiehi _8659__133 (.L_HI(net133));
 sg13g2_tiehi _8240__134 (.L_HI(net134));
 sg13g2_tiehi _8465__135 (.L_HI(net135));
 sg13g2_tiehi _8239__136 (.L_HI(net136));
 sg13g2_tiehi _8594__137 (.L_HI(net137));
 sg13g2_tiehi _8238__138 (.L_HI(net138));
 sg13g2_tiehi _8464__139 (.L_HI(net139));
 sg13g2_tiehi _8237__140 (.L_HI(net140));
 sg13g2_tiehi _8637__141 (.L_HI(net141));
 sg13g2_tiehi _8236__142 (.L_HI(net142));
 sg13g2_tiehi _8463__143 (.L_HI(net143));
 sg13g2_tiehi _8235__144 (.L_HI(net144));
 sg13g2_tiehi _8593__145 (.L_HI(net145));
 sg13g2_tiehi _8234__146 (.L_HI(net146));
 sg13g2_tiehi _8462__147 (.L_HI(net147));
 sg13g2_tiehi _8233__148 (.L_HI(net148));
 sg13g2_tiehi _8675__149 (.L_HI(net149));
 sg13g2_tiehi _8232__150 (.L_HI(net150));
 sg13g2_tiehi _8461__151 (.L_HI(net151));
 sg13g2_tiehi _8231__152 (.L_HI(net152));
 sg13g2_tiehi _8592__153 (.L_HI(net153));
 sg13g2_tiehi _8230__154 (.L_HI(net154));
 sg13g2_tiehi _8460__155 (.L_HI(net155));
 sg13g2_tiehi _8229__156 (.L_HI(net156));
 sg13g2_tiehi _8636__157 (.L_HI(net157));
 sg13g2_tiehi _8228__158 (.L_HI(net158));
 sg13g2_tiehi _8459__159 (.L_HI(net159));
 sg13g2_tiehi _8227__160 (.L_HI(net160));
 sg13g2_tiehi _8591__161 (.L_HI(net161));
 sg13g2_tiehi _8226__162 (.L_HI(net162));
 sg13g2_tiehi _8458__163 (.L_HI(net163));
 sg13g2_tiehi _8225__164 (.L_HI(net164));
 sg13g2_tiehi _8658__165 (.L_HI(net165));
 sg13g2_tiehi _8224__166 (.L_HI(net166));
 sg13g2_tiehi _8457__167 (.L_HI(net167));
 sg13g2_tiehi _8223__168 (.L_HI(net168));
 sg13g2_tiehi _8590__169 (.L_HI(net169));
 sg13g2_tiehi _8222__170 (.L_HI(net170));
 sg13g2_tiehi _8456__171 (.L_HI(net171));
 sg13g2_tiehi _8221__172 (.L_HI(net172));
 sg13g2_tiehi _8635__173 (.L_HI(net173));
 sg13g2_tiehi _8220__174 (.L_HI(net174));
 sg13g2_tiehi _8455__175 (.L_HI(net175));
 sg13g2_tiehi _8219__176 (.L_HI(net176));
 sg13g2_tiehi _8589__177 (.L_HI(net177));
 sg13g2_tiehi _8218__178 (.L_HI(net178));
 sg13g2_tiehi _8454__179 (.L_HI(net179));
 sg13g2_tiehi _8217__180 (.L_HI(net180));
 sg13g2_tiehi _8669__181 (.L_HI(net181));
 sg13g2_tiehi _8216__182 (.L_HI(net182));
 sg13g2_tiehi _8453__183 (.L_HI(net183));
 sg13g2_tiehi _8215__184 (.L_HI(net184));
 sg13g2_tiehi _8588__185 (.L_HI(net185));
 sg13g2_tiehi _8214__186 (.L_HI(net186));
 sg13g2_tiehi _8452__187 (.L_HI(net187));
 sg13g2_tiehi _8213__188 (.L_HI(net188));
 sg13g2_tiehi _8634__189 (.L_HI(net189));
 sg13g2_tiehi _8212__190 (.L_HI(net190));
 sg13g2_tiehi _8451__191 (.L_HI(net191));
 sg13g2_tiehi _8211__192 (.L_HI(net192));
 sg13g2_tiehi _8587__193 (.L_HI(net193));
 sg13g2_tiehi _8210__194 (.L_HI(net194));
 sg13g2_tiehi _8450__195 (.L_HI(net195));
 sg13g2_tiehi _8209__196 (.L_HI(net196));
 sg13g2_tiehi _8657__197 (.L_HI(net197));
 sg13g2_tiehi _8208__198 (.L_HI(net198));
 sg13g2_tiehi _8449__199 (.L_HI(net199));
 sg13g2_tiehi _8207__200 (.L_HI(net200));
 sg13g2_tiehi _8586__201 (.L_HI(net201));
 sg13g2_tiehi _8206__202 (.L_HI(net202));
 sg13g2_tiehi _8448__203 (.L_HI(net203));
 sg13g2_tiehi _8205__204 (.L_HI(net204));
 sg13g2_tiehi _8633__205 (.L_HI(net205));
 sg13g2_tiehi _8204__206 (.L_HI(net206));
 sg13g2_tiehi _8447__207 (.L_HI(net207));
 sg13g2_tiehi _8203__208 (.L_HI(net208));
 sg13g2_tiehi _8585__209 (.L_HI(net209));
 sg13g2_tiehi _8202__210 (.L_HI(net210));
 sg13g2_tiehi _8446__211 (.L_HI(net211));
 sg13g2_tiehi _8201__212 (.L_HI(net212));
 sg13g2_tiehi _8679__213 (.L_HI(net213));
 sg13g2_tiehi _8200__214 (.L_HI(net214));
 sg13g2_tiehi _8445__215 (.L_HI(net215));
 sg13g2_tiehi _8199__216 (.L_HI(net216));
 sg13g2_tiehi _8584__217 (.L_HI(net217));
 sg13g2_tiehi _8198__218 (.L_HI(net218));
 sg13g2_tiehi _8444__219 (.L_HI(net219));
 sg13g2_tiehi _8197__220 (.L_HI(net220));
 sg13g2_tiehi _8632__221 (.L_HI(net221));
 sg13g2_tiehi _8196__222 (.L_HI(net222));
 sg13g2_tiehi _8443__223 (.L_HI(net223));
 sg13g2_tiehi _8195__224 (.L_HI(net224));
 sg13g2_tiehi _8583__225 (.L_HI(net225));
 sg13g2_tiehi _8194__226 (.L_HI(net226));
 sg13g2_tiehi _8442__227 (.L_HI(net227));
 sg13g2_tiehi _8193__228 (.L_HI(net228));
 sg13g2_tiehi _8656__229 (.L_HI(net229));
 sg13g2_tiehi _8192__230 (.L_HI(net230));
 sg13g2_tiehi _8441__231 (.L_HI(net231));
 sg13g2_tiehi _8191__232 (.L_HI(net232));
 sg13g2_tiehi _8582__233 (.L_HI(net233));
 sg13g2_tiehi _8190__234 (.L_HI(net234));
 sg13g2_tiehi _8440__235 (.L_HI(net235));
 sg13g2_tiehi _8189__236 (.L_HI(net236));
 sg13g2_tiehi _8631__237 (.L_HI(net237));
 sg13g2_tiehi _8188__238 (.L_HI(net238));
 sg13g2_tiehi _8439__239 (.L_HI(net239));
 sg13g2_tiehi _8187__240 (.L_HI(net240));
 sg13g2_tiehi _8581__241 (.L_HI(net241));
 sg13g2_tiehi _8186__242 (.L_HI(net242));
 sg13g2_tiehi _8438__243 (.L_HI(net243));
 sg13g2_tiehi _8185__244 (.L_HI(net244));
 sg13g2_tiehi _8668__245 (.L_HI(net245));
 sg13g2_tiehi _8184__246 (.L_HI(net246));
 sg13g2_tiehi _8437__247 (.L_HI(net247));
 sg13g2_tiehi _8183__248 (.L_HI(net248));
 sg13g2_tiehi _8580__249 (.L_HI(net249));
 sg13g2_tiehi _8182__250 (.L_HI(net250));
 sg13g2_tiehi _8436__251 (.L_HI(net251));
 sg13g2_tiehi _8181__252 (.L_HI(net252));
 sg13g2_tiehi _8630__253 (.L_HI(net253));
 sg13g2_tiehi _8180__254 (.L_HI(net254));
 sg13g2_tiehi _8435__255 (.L_HI(net255));
 sg13g2_tiehi _8179__256 (.L_HI(net256));
 sg13g2_tiehi _8579__257 (.L_HI(net257));
 sg13g2_tiehi _8178__258 (.L_HI(net258));
 sg13g2_tiehi _8434__259 (.L_HI(net259));
 sg13g2_tiehi _8177__260 (.L_HI(net260));
 sg13g2_tiehi _8655__261 (.L_HI(net261));
 sg13g2_tiehi _8176__262 (.L_HI(net262));
 sg13g2_tiehi _8433__263 (.L_HI(net263));
 sg13g2_tiehi _8175__264 (.L_HI(net264));
 sg13g2_tiehi _8578__265 (.L_HI(net265));
 sg13g2_tiehi _8174__266 (.L_HI(net266));
 sg13g2_tiehi _8432__267 (.L_HI(net267));
 sg13g2_tiehi _8173__268 (.L_HI(net268));
 sg13g2_tiehi _8629__269 (.L_HI(net269));
 sg13g2_tiehi _8172__270 (.L_HI(net270));
 sg13g2_tiehi _8431__271 (.L_HI(net271));
 sg13g2_tiehi _8171__272 (.L_HI(net272));
 sg13g2_tiehi _8577__273 (.L_HI(net273));
 sg13g2_tiehi _8170__274 (.L_HI(net274));
 sg13g2_tiehi _8430__275 (.L_HI(net275));
 sg13g2_tiehi _8169__276 (.L_HI(net276));
 sg13g2_tiehi _8674__277 (.L_HI(net277));
 sg13g2_tiehi _8168__278 (.L_HI(net278));
 sg13g2_tiehi _8429__279 (.L_HI(net279));
 sg13g2_tiehi _8167__280 (.L_HI(net280));
 sg13g2_tiehi _8576__281 (.L_HI(net281));
 sg13g2_tiehi _8166__282 (.L_HI(net282));
 sg13g2_tiehi _8428__283 (.L_HI(net283));
 sg13g2_tiehi _8165__284 (.L_HI(net284));
 sg13g2_tiehi _8628__285 (.L_HI(net285));
 sg13g2_tiehi _8164__286 (.L_HI(net286));
 sg13g2_tiehi _8427__287 (.L_HI(net287));
 sg13g2_tiehi _8163__288 (.L_HI(net288));
 sg13g2_tiehi _8575__289 (.L_HI(net289));
 sg13g2_tiehi _8162__290 (.L_HI(net290));
 sg13g2_tiehi _8161__291 (.L_HI(net291));
 sg13g2_tiehi _8426__292 (.L_HI(net292));
 sg13g2_tiehi _8160__293 (.L_HI(net293));
 sg13g2_tiehi _8654__294 (.L_HI(net294));
 sg13g2_tiehi _8159__295 (.L_HI(net295));
 sg13g2_tiehi _8425__296 (.L_HI(net296));
 sg13g2_tiehi _8158__297 (.L_HI(net297));
 sg13g2_tiehi _8574__298 (.L_HI(net298));
 sg13g2_tiehi _8157__299 (.L_HI(net299));
 sg13g2_tiehi _8424__300 (.L_HI(net300));
 sg13g2_tiehi _8156__301 (.L_HI(net301));
 sg13g2_tiehi _8627__302 (.L_HI(net302));
 sg13g2_tiehi _8155__303 (.L_HI(net303));
 sg13g2_tiehi _8423__304 (.L_HI(net304));
 sg13g2_tiehi _8154__305 (.L_HI(net305));
 sg13g2_tiehi _8573__306 (.L_HI(net306));
 sg13g2_tiehi _8153__307 (.L_HI(net307));
 sg13g2_tiehi _8422__308 (.L_HI(net308));
 sg13g2_tiehi _8152__309 (.L_HI(net309));
 sg13g2_tiehi _8667__310 (.L_HI(net310));
 sg13g2_tiehi _8151__311 (.L_HI(net311));
 sg13g2_tiehi _8421__312 (.L_HI(net312));
 sg13g2_tiehi _8150__313 (.L_HI(net313));
 sg13g2_tiehi _8572__314 (.L_HI(net314));
 sg13g2_tiehi _8149__315 (.L_HI(net315));
 sg13g2_tiehi _8420__316 (.L_HI(net316));
 sg13g2_tiehi _8148__317 (.L_HI(net317));
 sg13g2_tiehi _8626__318 (.L_HI(net318));
 sg13g2_tiehi _8147__319 (.L_HI(net319));
 sg13g2_tiehi _8419__320 (.L_HI(net320));
 sg13g2_tiehi _8146__321 (.L_HI(net321));
 sg13g2_tiehi _8145__322 (.L_HI(net322));
 sg13g2_tiehi _8571__323 (.L_HI(net323));
 sg13g2_tiehi _8144__324 (.L_HI(net324));
 sg13g2_tiehi _8418__325 (.L_HI(net325));
 sg13g2_tiehi _8143__326 (.L_HI(net326));
 sg13g2_tiehi _8653__327 (.L_HI(net327));
 sg13g2_tiehi _8142__328 (.L_HI(net328));
 sg13g2_tiehi _8417__329 (.L_HI(net329));
 sg13g2_tiehi _8141__330 (.L_HI(net330));
 sg13g2_tiehi _8570__331 (.L_HI(net331));
 sg13g2_tiehi _8140__332 (.L_HI(net332));
 sg13g2_tiehi _8416__333 (.L_HI(net333));
 sg13g2_tiehi _8139__334 (.L_HI(net334));
 sg13g2_tiehi _8625__335 (.L_HI(net335));
 sg13g2_tiehi _8138__336 (.L_HI(net336));
 sg13g2_tiehi _8415__337 (.L_HI(net337));
 sg13g2_tiehi _8137__338 (.L_HI(net338));
 sg13g2_tiehi _8569__339 (.L_HI(net339));
 sg13g2_tiehi _8136__340 (.L_HI(net340));
 sg13g2_tiehi _8414__341 (.L_HI(net341));
 sg13g2_tiehi _8135__342 (.L_HI(net342));
 sg13g2_tiehi _8677__343 (.L_HI(net343));
 sg13g2_tiehi _8134__344 (.L_HI(net344));
 sg13g2_tiehi _8413__345 (.L_HI(net345));
 sg13g2_tiehi _8133__346 (.L_HI(net346));
 sg13g2_tiehi _8568__347 (.L_HI(net347));
 sg13g2_tiehi _8132__348 (.L_HI(net348));
 sg13g2_tiehi _8412__349 (.L_HI(net349));
 sg13g2_tiehi _8131__350 (.L_HI(net350));
 sg13g2_tiehi _8624__351 (.L_HI(net351));
 sg13g2_tiehi _8130__352 (.L_HI(net352));
 sg13g2_tiehi _8411__353 (.L_HI(net353));
 sg13g2_tiehi _8129__354 (.L_HI(net354));
 sg13g2_tiehi _8567__355 (.L_HI(net355));
 sg13g2_tiehi _8128__356 (.L_HI(net356));
 sg13g2_tiehi _8410__357 (.L_HI(net357));
 sg13g2_tiehi _8127__358 (.L_HI(net358));
 sg13g2_tiehi _8652__359 (.L_HI(net359));
 sg13g2_tiehi _8126__360 (.L_HI(net360));
 sg13g2_tiehi _8409__361 (.L_HI(net361));
 sg13g2_tiehi _8125__362 (.L_HI(net362));
 sg13g2_tiehi _8566__363 (.L_HI(net363));
 sg13g2_tiehi _8124__364 (.L_HI(net364));
 sg13g2_tiehi _8408__365 (.L_HI(net365));
 sg13g2_tiehi _8123__366 (.L_HI(net366));
 sg13g2_tiehi _8623__367 (.L_HI(net367));
 sg13g2_tiehi _8122__368 (.L_HI(net368));
 sg13g2_tiehi _8407__369 (.L_HI(net369));
 sg13g2_tiehi _8121__370 (.L_HI(net370));
 sg13g2_tiehi _8565__371 (.L_HI(net371));
 sg13g2_tiehi _8120__372 (.L_HI(net372));
 sg13g2_tiehi _8406__373 (.L_HI(net373));
 sg13g2_tiehi _8119__374 (.L_HI(net374));
 sg13g2_tiehi _8666__375 (.L_HI(net375));
 sg13g2_tiehi _8118__376 (.L_HI(net376));
 sg13g2_tiehi _8405__377 (.L_HI(net377));
 sg13g2_tiehi _8117__378 (.L_HI(net378));
 sg13g2_tiehi _8564__379 (.L_HI(net379));
 sg13g2_tiehi _8116__380 (.L_HI(net380));
 sg13g2_tiehi _8404__381 (.L_HI(net381));
 sg13g2_tiehi _8115__382 (.L_HI(net382));
 sg13g2_tiehi _8622__383 (.L_HI(net383));
 sg13g2_tiehi _8114__384 (.L_HI(net384));
 sg13g2_tiehi _8403__385 (.L_HI(net385));
 sg13g2_tiehi _8113__386 (.L_HI(net386));
 sg13g2_tiehi _8112__387 (.L_HI(net387));
 sg13g2_tiehi _8563__388 (.L_HI(net388));
 sg13g2_tiehi _8111__389 (.L_HI(net389));
 sg13g2_tiehi _8402__390 (.L_HI(net390));
 sg13g2_tiehi _8110__391 (.L_HI(net391));
 sg13g2_tiehi _8651__392 (.L_HI(net392));
 sg13g2_tiehi _8109__393 (.L_HI(net393));
 sg13g2_tiehi _8401__394 (.L_HI(net394));
 sg13g2_tiehi _8108__395 (.L_HI(net395));
 sg13g2_tiehi _8562__396 (.L_HI(net396));
 sg13g2_tiehi _8107__397 (.L_HI(net397));
 sg13g2_tiehi _8400__398 (.L_HI(net398));
 sg13g2_tiehi _8106__399 (.L_HI(net399));
 sg13g2_tiehi _8621__400 (.L_HI(net400));
 sg13g2_tiehi _8105__401 (.L_HI(net401));
 sg13g2_tiehi _8399__402 (.L_HI(net402));
 sg13g2_tiehi _8104__403 (.L_HI(net403));
 sg13g2_tiehi _8561__404 (.L_HI(net404));
 sg13g2_tiehi _8103__405 (.L_HI(net405));
 sg13g2_tiehi _8398__406 (.L_HI(net406));
 sg13g2_tiehi _8102__407 (.L_HI(net407));
 sg13g2_tiehi _8101__408 (.L_HI(net408));
 sg13g2_tiehi _8100__409 (.L_HI(net409));
 sg13g2_tiehi _8099__410 (.L_HI(net410));
 sg13g2_tiehi _8098__411 (.L_HI(net411));
 sg13g2_tiehi _8097__412 (.L_HI(net412));
 sg13g2_tiehi _8096__413 (.L_HI(net413));
 sg13g2_tiehi _8095__414 (.L_HI(net414));
 sg13g2_tiehi _8094__415 (.L_HI(net415));
 sg13g2_tiehi _8093__416 (.L_HI(net416));
 sg13g2_tiehi _8092__417 (.L_HI(net417));
 sg13g2_tiehi _8091__418 (.L_HI(net418));
 sg13g2_tiehi _8090__419 (.L_HI(net419));
 sg13g2_tiehi _8089__420 (.L_HI(net420));
 sg13g2_tiehi _8088__421 (.L_HI(net421));
 sg13g2_tiehi _8087__422 (.L_HI(net422));
 sg13g2_tiehi _8086__423 (.L_HI(net423));
 sg13g2_tiehi _8085__424 (.L_HI(net424));
 sg13g2_tiehi _8084__425 (.L_HI(net425));
 sg13g2_tiehi _8083__426 (.L_HI(net426));
 sg13g2_tiehi _8082__427 (.L_HI(net427));
 sg13g2_tiehi _8081__428 (.L_HI(net428));
 sg13g2_tiehi _8080__429 (.L_HI(net429));
 sg13g2_tiehi _8079__430 (.L_HI(net430));
 sg13g2_tiehi _8078__431 (.L_HI(net431));
 sg13g2_tiehi _8077__432 (.L_HI(net432));
 sg13g2_tiehi _8076__433 (.L_HI(net433));
 sg13g2_tiehi _8075__434 (.L_HI(net434));
 sg13g2_tiehi _8074__435 (.L_HI(net435));
 sg13g2_tiehi _8073__436 (.L_HI(net436));
 sg13g2_tiehi _8072__437 (.L_HI(net437));
 sg13g2_tiehi _8071__438 (.L_HI(net438));
 sg13g2_tiehi _8070__439 (.L_HI(net439));
 sg13g2_tiehi _8069__440 (.L_HI(net440));
 sg13g2_tiehi _8068__441 (.L_HI(net441));
 sg13g2_tiehi _8067__442 (.L_HI(net442));
 sg13g2_tiehi _8066__443 (.L_HI(net443));
 sg13g2_tiehi _8065__444 (.L_HI(net444));
 sg13g2_tiehi _8673__445 (.L_HI(net445));
 sg13g2_tiehi _8064__446 (.L_HI(net446));
 sg13g2_tiehi _8397__447 (.L_HI(net447));
 sg13g2_tiehi _8063__448 (.L_HI(net448));
 sg13g2_tiehi _8560__449 (.L_HI(net449));
 sg13g2_tiehi _8062__450 (.L_HI(net450));
 sg13g2_tiehi _8396__451 (.L_HI(net451));
 sg13g2_tiehi _8061__452 (.L_HI(net452));
 sg13g2_tiehi _8395__453 (.L_HI(net453));
 sg13g2_tiehi _8060__454 (.L_HI(net454));
 sg13g2_tiehi _8620__455 (.L_HI(net455));
 sg13g2_tiehi _8059__456 (.L_HI(net456));
 sg13g2_tiehi _8394__457 (.L_HI(net457));
 sg13g2_tiehi _8058__458 (.L_HI(net458));
 sg13g2_tiehi _8559__459 (.L_HI(net459));
 sg13g2_tiehi _8057__460 (.L_HI(net460));
 sg13g2_tiehi _8393__461 (.L_HI(net461));
 sg13g2_tiehi _8056__462 (.L_HI(net462));
 sg13g2_tiehi _8650__463 (.L_HI(net463));
 sg13g2_tiehi _8055__464 (.L_HI(net464));
 sg13g2_tiehi _8392__465 (.L_HI(net465));
 sg13g2_tiehi _8054__466 (.L_HI(net466));
 sg13g2_tiehi _8558__467 (.L_HI(net467));
 sg13g2_tiehi _8053__468 (.L_HI(net468));
 sg13g2_tiehi _8391__469 (.L_HI(net469));
 sg13g2_tiehi _8052__470 (.L_HI(net470));
 sg13g2_tiehi _8619__471 (.L_HI(net471));
 sg13g2_tiehi _8051__472 (.L_HI(net472));
 sg13g2_tiehi _8390__473 (.L_HI(net473));
 sg13g2_tiehi _8050__474 (.L_HI(net474));
 sg13g2_tiehi _8557__475 (.L_HI(net475));
 sg13g2_tiehi _8049__476 (.L_HI(net476));
 sg13g2_tiehi _8389__477 (.L_HI(net477));
 sg13g2_tiehi _8048__478 (.L_HI(net478));
 sg13g2_tiehi _8665__479 (.L_HI(net479));
 sg13g2_tiehi _8047__480 (.L_HI(net480));
 sg13g2_tiehi _8388__481 (.L_HI(net481));
 sg13g2_tiehi _8046__482 (.L_HI(net482));
 sg13g2_tiehi _8556__483 (.L_HI(net483));
 sg13g2_tiehi _8045__484 (.L_HI(net484));
 sg13g2_tiehi _8387__485 (.L_HI(net485));
 sg13g2_tiehi _8044__486 (.L_HI(net486));
 sg13g2_tiehi _8618__487 (.L_HI(net487));
 sg13g2_tiehi _8043__488 (.L_HI(net488));
 sg13g2_tiehi _8386__489 (.L_HI(net489));
 sg13g2_tiehi _8042__490 (.L_HI(net490));
 sg13g2_tiehi _8555__491 (.L_HI(net491));
 sg13g2_tiehi _8041__492 (.L_HI(net492));
 sg13g2_tiehi _8385__493 (.L_HI(net493));
 sg13g2_tiehi _8040__494 (.L_HI(net494));
 sg13g2_tiehi _8649__495 (.L_HI(net495));
 sg13g2_tiehi _8039__496 (.L_HI(net496));
 sg13g2_tiehi _8384__497 (.L_HI(net497));
 sg13g2_tiehi _8038__498 (.L_HI(net498));
 sg13g2_tiehi _8554__499 (.L_HI(net499));
 sg13g2_tiehi _8037__500 (.L_HI(net500));
 sg13g2_tiehi _8383__501 (.L_HI(net501));
 sg13g2_tiehi _8036__502 (.L_HI(net502));
 sg13g2_tiehi _8617__503 (.L_HI(net503));
 sg13g2_tiehi _8035__504 (.L_HI(net504));
 sg13g2_tiehi _8382__505 (.L_HI(net505));
 sg13g2_tiehi _8034__506 (.L_HI(net506));
 sg13g2_tiehi _8381__507 (.L_HI(net507));
 sg13g2_tiehi _8033__508 (.L_HI(net508));
 sg13g2_tiehi _8380__509 (.L_HI(net509));
 sg13g2_tiehi _8032__510 (.L_HI(net510));
 sg13g2_tiehi _8379__511 (.L_HI(net511));
 sg13g2_tiehi _8031__512 (.L_HI(net512));
 sg13g2_tiehi _8378__513 (.L_HI(net513));
 sg13g2_tiehi _8030__514 (.L_HI(net514));
 sg13g2_tiehi _8377__515 (.L_HI(net515));
 sg13g2_tiehi _8029__516 (.L_HI(net516));
 sg13g2_tiehi _8376__517 (.L_HI(net517));
 sg13g2_tiehi _8028__518 (.L_HI(net518));
 sg13g2_tiehi _8375__519 (.L_HI(net519));
 sg13g2_tiehi _8027__520 (.L_HI(net520));
 sg13g2_tiehi _8374__521 (.L_HI(net521));
 sg13g2_tiehi _8026__522 (.L_HI(net522));
 sg13g2_tiehi _8553__523 (.L_HI(net523));
 sg13g2_tiehi _8025__524 (.L_HI(net524));
 sg13g2_tiehi _8373__525 (.L_HI(net525));
 sg13g2_tiehi _8014__526 (.L_HI(net526));
 sg13g2_tiehi _8013__527 (.L_HI(net527));
 sg13g2_tiehi _8372__528 (.L_HI(net528));
 sg13g2_tiehi _8012__529 (.L_HI(net529));
 sg13g2_tiehi _8552__530 (.L_HI(net530));
 sg13g2_tiehi _8011__531 (.L_HI(net531));
 sg13g2_tiehi _8371__532 (.L_HI(net532));
 sg13g2_tiehi _8010__533 (.L_HI(net533));
 sg13g2_tiehi _8616__534 (.L_HI(net534));
 sg13g2_tiehi _8009__535 (.L_HI(net535));
 sg13g2_tiehi _8370__536 (.L_HI(net536));
 sg13g2_tiehi _8008__537 (.L_HI(net537));
 sg13g2_tiehi _8551__538 (.L_HI(net538));
 sg13g2_tiehi _8007__539 (.L_HI(net539));
 sg13g2_tiehi _8369__540 (.L_HI(net540));
 sg13g2_tiehi _8006__541 (.L_HI(net541));
 sg13g2_tiehi _8648__542 (.L_HI(net542));
 sg13g2_tiehi _8005__543 (.L_HI(net543));
 sg13g2_tiehi _8368__544 (.L_HI(net544));
 sg13g2_tiehi _8004__545 (.L_HI(net545));
 sg13g2_tiehi _8550__546 (.L_HI(net546));
 sg13g2_tiehi _8003__547 (.L_HI(net547));
 sg13g2_tiehi _8367__548 (.L_HI(net548));
 sg13g2_tiehi _8002__549 (.L_HI(net549));
 sg13g2_tiehi _8615__550 (.L_HI(net550));
 sg13g2_tiehi _8001__551 (.L_HI(net551));
 sg13g2_tiehi _8366__552 (.L_HI(net552));
 sg13g2_tiehi _8000__553 (.L_HI(net553));
 sg13g2_tiehi _7999__554 (.L_HI(net554));
 sg13g2_tiehi _7998__555 (.L_HI(net555));
 sg13g2_tiehi _7997__556 (.L_HI(net556));
 sg13g2_tiehi _7996__557 (.L_HI(net557));
 sg13g2_tiehi _7995__558 (.L_HI(net558));
 sg13g2_tiehi _7994__559 (.L_HI(net559));
 sg13g2_tiehi _7993__560 (.L_HI(net560));
 sg13g2_tiehi _7992__561 (.L_HI(net561));
 sg13g2_tiehi _8549__562 (.L_HI(net562));
 sg13g2_tiehi _7991__563 (.L_HI(net563));
 sg13g2_tiehi _8365__564 (.L_HI(net564));
 sg13g2_tiehi _7987__565 (.L_HI(net565));
 sg13g2_tiehi _8364__566 (.L_HI(net566));
 sg13g2_tiehi _7986__567 (.L_HI(net567));
 sg13g2_tiehi _8664__568 (.L_HI(net568));
 sg13g2_tiehi _7985__569 (.L_HI(net569));
 sg13g2_tiehi _8363__570 (.L_HI(net570));
 sg13g2_tiehi _7984__571 (.L_HI(net571));
 sg13g2_tiehi _8548__572 (.L_HI(net572));
 sg13g2_tiehi _7983__573 (.L_HI(net573));
 sg13g2_tiehi _8362__574 (.L_HI(net574));
 sg13g2_tiehi _7982__575 (.L_HI(net575));
 sg13g2_tiehi _8614__576 (.L_HI(net576));
 sg13g2_tiehi _7981__577 (.L_HI(net577));
 sg13g2_tiehi _8361__578 (.L_HI(net578));
 sg13g2_tiehi _7980__579 (.L_HI(net579));
 sg13g2_tiehi _8547__580 (.L_HI(net580));
 sg13g2_tiehi _7979__581 (.L_HI(net581));
 sg13g2_tiehi _8360__582 (.L_HI(net582));
 sg13g2_tiehi _7978__583 (.L_HI(net583));
 sg13g2_tiehi _8647__584 (.L_HI(net584));
 sg13g2_tiehi _7977__585 (.L_HI(net585));
 sg13g2_tiehi _8359__586 (.L_HI(net586));
 sg13g2_tiehi _7976__587 (.L_HI(net587));
 sg13g2_tiehi _8546__588 (.L_HI(net588));
 sg13g2_tiehi _7975__589 (.L_HI(net589));
 sg13g2_tiehi _8358__590 (.L_HI(net590));
 sg13g2_tiehi _7974__591 (.L_HI(net591));
 sg13g2_tiehi _8613__592 (.L_HI(net592));
 sg13g2_tiehi _8024__593 (.L_HI(net593));
 sg13g2_tiehi _8513__594 (.L_HI(net594));
 sg13g2_tiehi _7973__595 (.L_HI(net595));
 sg13g2_tiehi _8357__596 (.L_HI(net596));
 sg13g2_tiehi _7972__597 (.L_HI(net597));
 sg13g2_tiehi _8545__598 (.L_HI(net598));
 sg13g2_tiehi _7971__599 (.L_HI(net599));
 sg13g2_tiehi _8356__600 (.L_HI(net600));
 sg13g2_tiehi _7970__601 (.L_HI(net601));
 sg13g2_tiehi _8672__602 (.L_HI(net602));
 sg13g2_tiehi _7969__603 (.L_HI(net603));
 sg13g2_tiehi _8355__604 (.L_HI(net604));
 sg13g2_tiehi _7968__605 (.L_HI(net605));
 sg13g2_tiehi _8544__606 (.L_HI(net606));
 sg13g2_tiehi _7967__607 (.L_HI(net607));
 sg13g2_tiehi _8354__608 (.L_HI(net608));
 sg13g2_tiehi _7966__609 (.L_HI(net609));
 sg13g2_tiehi _8612__610 (.L_HI(net610));
 sg13g2_tiehi _7965__611 (.L_HI(net611));
 sg13g2_tiehi _8353__612 (.L_HI(net612));
 sg13g2_tiehi _7964__613 (.L_HI(net613));
 sg13g2_tiehi _8543__614 (.L_HI(net614));
 sg13g2_tiehi _7963__615 (.L_HI(net615));
 sg13g2_tiehi _8352__616 (.L_HI(net616));
 sg13g2_tiehi _7962__617 (.L_HI(net617));
 sg13g2_tiehi _8351__618 (.L_HI(net618));
 sg13g2_tiehi _7961__619 (.L_HI(net619));
 sg13g2_tiehi _8646__620 (.L_HI(net620));
 sg13g2_tiehi _7960__621 (.L_HI(net621));
 sg13g2_tiehi _8350__622 (.L_HI(net622));
 sg13g2_tiehi _7959__623 (.L_HI(net623));
 sg13g2_tiehi _8542__624 (.L_HI(net624));
 sg13g2_tiehi _7958__625 (.L_HI(net625));
 sg13g2_tiehi _8349__626 (.L_HI(net626));
 sg13g2_tiehi _7957__627 (.L_HI(net627));
 sg13g2_tiehi _8611__628 (.L_HI(net628));
 sg13g2_tiehi _7956__629 (.L_HI(net629));
 sg13g2_tiehi _8348__630 (.L_HI(net630));
 sg13g2_tiehi _7955__631 (.L_HI(net631));
 sg13g2_tiehi _8541__632 (.L_HI(net632));
 sg13g2_tiehi _7954__633 (.L_HI(net633));
 sg13g2_tiehi _8347__634 (.L_HI(net634));
 sg13g2_tiehi _7953__635 (.L_HI(net635));
 sg13g2_tiehi _8663__636 (.L_HI(net636));
 sg13g2_tiehi _7952__637 (.L_HI(net637));
 sg13g2_tiehi _8346__638 (.L_HI(net638));
 sg13g2_tiehi _7951__639 (.L_HI(net639));
 sg13g2_tiehi _8540__640 (.L_HI(net640));
 sg13g2_tiehi _7950__641 (.L_HI(net641));
 sg13g2_tiehi _8345__642 (.L_HI(net642));
 sg13g2_tiehi _7949__643 (.L_HI(net643));
 sg13g2_tiehi _7948__644 (.L_HI(net644));
 sg13g2_tiehi _7947__645 (.L_HI(net645));
 sg13g2_tiehi _7946__646 (.L_HI(net646));
 sg13g2_tiehi _7945__647 (.L_HI(net647));
 sg13g2_tiehi _8610__648 (.L_HI(net648));
 sg13g2_tiehi _8344__649 (.L_HI(net649));
 sg13g2_tiehi _8539__650 (.L_HI(net650));
 sg13g2_tiehi _8343__651 (.L_HI(net651));
 sg13g2_tiehi _8645__652 (.L_HI(net652));
 sg13g2_tiehi _8342__653 (.L_HI(net653));
 sg13g2_tiehi _8538__654 (.L_HI(net654));
 sg13g2_tiehi _8341__655 (.L_HI(net655));
 sg13g2_tiehi _8609__656 (.L_HI(net656));
 sg13g2_tiehi _8340__657 (.L_HI(net657));
 sg13g2_tiehi _8537__658 (.L_HI(net658));
 sg13g2_tiehi _8339__659 (.L_HI(net659));
 sg13g2_tiehi _8676__660 (.L_HI(net660));
 sg13g2_tiehi _8338__661 (.L_HI(net661));
 sg13g2_tiehi _8536__662 (.L_HI(net662));
 sg13g2_tiehi _8337__663 (.L_HI(net663));
 sg13g2_tiehi _8608__664 (.L_HI(net664));
 sg13g2_tiehi _8336__665 (.L_HI(net665));
 sg13g2_tiehi _8535__666 (.L_HI(net666));
 sg13g2_tiehi _8335__667 (.L_HI(net667));
 sg13g2_tiehi _8644__668 (.L_HI(net668));
 sg13g2_tiehi _8334__669 (.L_HI(net669));
 sg13g2_tiehi _8534__670 (.L_HI(net670));
 sg13g2_tiehi _8333__671 (.L_HI(net671));
 sg13g2_tiehi _8607__672 (.L_HI(net672));
 sg13g2_tiehi _8332__673 (.L_HI(net673));
 sg13g2_tiehi _8533__674 (.L_HI(net674));
 sg13g2_tiehi _8331__675 (.L_HI(net675));
 sg13g2_tiehi _8662__676 (.L_HI(net676));
 sg13g2_tiehi _8330__677 (.L_HI(net677));
 sg13g2_tiehi _8532__678 (.L_HI(net678));
 sg13g2_tiehi _8329__679 (.L_HI(net679));
 sg13g2_tiehi _8606__680 (.L_HI(net680));
 sg13g2_tiehi _8328__681 (.L_HI(net681));
 sg13g2_tiehi _8531__682 (.L_HI(net682));
 sg13g2_tiehi _8327__683 (.L_HI(net683));
 sg13g2_tiehi _8643__684 (.L_HI(net684));
 sg13g2_tiehi _8326__685 (.L_HI(net685));
 sg13g2_tiehi _8325__686 (.L_HI(net686));
 sg13g2_tiehi _8530__687 (.L_HI(net687));
 sg13g2_tiehi _8324__688 (.L_HI(net688));
 sg13g2_tiehi _8605__689 (.L_HI(net689));
 sg13g2_tiehi _8323__690 (.L_HI(net690));
 sg13g2_tiehi _8529__691 (.L_HI(net691));
 sg13g2_tiehi _8322__692 (.L_HI(net692));
 sg13g2_tiehi _8671__693 (.L_HI(net693));
 sg13g2_tiehi _8321__694 (.L_HI(net694));
 sg13g2_tiehi _8528__695 (.L_HI(net695));
 sg13g2_tiehi _8320__696 (.L_HI(net696));
 sg13g2_tiehi _8604__697 (.L_HI(net697));
 sg13g2_tiehi _8319__698 (.L_HI(net698));
 sg13g2_tiehi _8527__699 (.L_HI(net699));
 sg13g2_tiehi _8318__700 (.L_HI(net700));
 sg13g2_tiehi _8642__701 (.L_HI(net701));
 sg13g2_tiehi _8317__702 (.L_HI(net702));
 sg13g2_tiehi _8526__703 (.L_HI(net703));
 sg13g2_tiehi _8316__704 (.L_HI(net704));
 sg13g2_tiehi _8603__705 (.L_HI(net705));
 sg13g2_tiehi _8315__706 (.L_HI(net706));
 sg13g2_tiehi _8525__707 (.L_HI(net707));
 sg13g2_tiehi _8314__708 (.L_HI(net708));
 sg13g2_tiehi _8661__709 (.L_HI(net709));
 sg13g2_tiehi _8313__710 (.L_HI(net710));
 sg13g2_tiehi _8524__711 (.L_HI(net711));
 sg13g2_tiehi _8312__712 (.L_HI(net712));
 sg13g2_tiehi _8602__713 (.L_HI(net713));
 sg13g2_tiehi _8311__714 (.L_HI(net714));
 sg13g2_tiehi _8523__715 (.L_HI(net715));
 sg13g2_tiehi _8310__716 (.L_HI(net716));
 sg13g2_tiehi _8641__717 (.L_HI(net717));
 sg13g2_tiehi _8309__718 (.L_HI(net718));
 sg13g2_tiehi _8522__719 (.L_HI(net719));
 sg13g2_tiehi _8308__720 (.L_HI(net720));
 sg13g2_tiehi _8601__721 (.L_HI(net721));
 sg13g2_tiehi _8307__722 (.L_HI(net722));
 sg13g2_tiehi _8521__723 (.L_HI(net723));
 sg13g2_tiehi _8306__724 (.L_HI(net724));
 sg13g2_tiehi _8520__725 (.L_HI(net725));
 sg13g2_tiehi _8305__726 (.L_HI(net726));
 sg13g2_tiehi _8519__727 (.L_HI(net727));
 sg13g2_tiehi _8304__728 (.L_HI(net728));
 sg13g2_tiehi _8518__729 (.L_HI(net729));
 sg13g2_tiehi _8303__730 (.L_HI(net730));
 sg13g2_tiehi _8517__731 (.L_HI(net731));
 sg13g2_tiehi _8302__732 (.L_HI(net732));
 sg13g2_tiehi _8516__733 (.L_HI(net733));
 sg13g2_tiehi _8301__734 (.L_HI(net734));
 sg13g2_tiehi _8678__735 (.L_HI(net735));
 sg13g2_tiehi _8300__736 (.L_HI(net736));
 sg13g2_tiehi _8299__737 (.L_HI(net737));
 sg13g2_tiehi _8600__738 (.L_HI(net738));
 sg13g2_tiehi _8298__739 (.L_HI(net739));
 sg13g2_tiehi _8512__740 (.L_HI(net740));
 sg13g2_tiehi _8297__741 (.L_HI(net741));
 sg13g2_tiehi _8640__742 (.L_HI(net742));
 sg13g2_tiehi _8296__743 (.L_HI(net743));
 sg13g2_tiehi _8511__744 (.L_HI(net744));
 sg13g2_tiehi _8295__745 (.L_HI(net745));
 sg13g2_tiehi _8599__746 (.L_HI(net746));
 sg13g2_tiehi _8294__747 (.L_HI(net747));
 sg13g2_tiehi _8510__748 (.L_HI(net748));
 sg13g2_tiehi _8293__749 (.L_HI(net749));
 sg13g2_tiehi _8660__750 (.L_HI(net750));
 sg13g2_tiehi _8292__751 (.L_HI(net751));
 sg13g2_tiehi _8509__752 (.L_HI(net752));
 sg13g2_tiehi _8291__753 (.L_HI(net753));
 sg13g2_tiehi _8598__754 (.L_HI(net754));
 sg13g2_tiehi _8290__755 (.L_HI(net755));
 sg13g2_tiehi _8508__756 (.L_HI(net756));
 sg13g2_tiehi _8289__757 (.L_HI(net757));
 sg13g2_tiehi _8639__758 (.L_HI(net758));
 sg13g2_tiehi _7944__759 (.L_HI(net759));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_chrismoos_led_controller_7 (.L_LO(net7));
 sg13g2_tielo tt_um_chrismoos_led_controller_8 (.L_LO(net8));
 sg13g2_tielo tt_um_chrismoos_led_controller_9 (.L_LO(net9));
 sg13g2_tielo tt_um_chrismoos_led_controller_10 (.L_LO(net10));
 sg13g2_tielo tt_um_chrismoos_led_controller_11 (.L_LO(net11));
 sg13g2_tielo tt_um_chrismoos_led_controller_12 (.L_LO(net12));
 sg13g2_tielo tt_um_chrismoos_led_controller_13 (.L_LO(net13));
 sg13g2_tielo tt_um_chrismoos_led_controller_14 (.L_LO(net14));
 sg13g2_tielo tt_um_chrismoos_led_controller_15 (.L_LO(net15));
 sg13g2_tielo tt_um_chrismoos_led_controller_16 (.L_LO(net16));
 sg13g2_tielo tt_um_chrismoos_led_controller_17 (.L_LO(net17));
 sg13g2_tielo tt_um_chrismoos_led_controller_18 (.L_LO(net18));
 sg13g2_tielo tt_um_chrismoos_led_controller_19 (.L_LO(net19));
 sg13g2_tielo tt_um_chrismoos_led_controller_20 (.L_LO(net20));
 sg13g2_tielo tt_um_chrismoos_led_controller_21 (.L_LO(net21));
 sg13g2_tielo tt_um_chrismoos_led_controller_22 (.L_LO(net22));
 sg13g2_tielo tt_um_chrismoos_led_controller_23 (.L_LO(net23));
 sg13g2_tiehi _7942__24 (.L_HI(net24));
 sg13g2_buf_1 _9434_ (.A(\led_controller.o_spi_miso ),
    .X(uio_out[0]));
 sg13g2_buf_1 _9435_ (.A(\led_controller.flash.o_cs_n ),
    .X(uo_out[0]));
 sg13g2_buf_1 _9436_ (.A(\led_controller.flash.master.o_mosi ),
    .X(uo_out[1]));
 sg13g2_buf_1 _9437_ (.A(\led_controller.flash.master.o_sck ),
    .X(uo_out[2]));
 sg13g2_buf_1 _9438_ (.A(\led_controller.o_data ),
    .X(uo_out[3]));
 sg13g2_buf_8 fanout821 (.A(_2658_),
    .X(net821));
 sg13g2_buf_8 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_8 fanout823 (.A(_1689_),
    .X(net823));
 sg13g2_buf_8 fanout824 (.A(_1216_),
    .X(net824));
 sg13g2_buf_8 fanout825 (.A(_1206_),
    .X(net825));
 sg13g2_buf_8 fanout826 (.A(_2758_),
    .X(net826));
 sg13g2_buf_8 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_8 fanout828 (.A(_2452_),
    .X(net828));
 sg13g2_buf_8 fanout829 (.A(_1237_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_1237_),
    .X(net830));
 sg13g2_buf_8 fanout831 (.A(_1138_),
    .X(net831));
 sg13g2_buf_8 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_8 fanout833 (.A(_2595_),
    .X(net833));
 sg13g2_buf_8 fanout834 (.A(_1235_),
    .X(net834));
 sg13g2_buf_1 fanout835 (.A(_1235_),
    .X(net835));
 sg13g2_buf_8 fanout836 (.A(_2259_),
    .X(net836));
 sg13g2_buf_8 fanout837 (.A(_2186_),
    .X(net837));
 sg13g2_buf_8 fanout838 (.A(_2186_),
    .X(net838));
 sg13g2_buf_8 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_8 fanout840 (.A(net842),
    .X(net840));
 sg13g2_buf_8 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_8 fanout842 (.A(_2088_),
    .X(net842));
 sg13g2_buf_8 fanout843 (.A(_2054_),
    .X(net843));
 sg13g2_buf_8 fanout844 (.A(_2022_),
    .X(net844));
 sg13g2_buf_8 fanout845 (.A(_1989_),
    .X(net845));
 sg13g2_buf_8 fanout846 (.A(_1895_),
    .X(net846));
 sg13g2_buf_8 fanout847 (.A(net849),
    .X(net847));
 sg13g2_buf_8 fanout848 (.A(net849),
    .X(net848));
 sg13g2_buf_8 fanout849 (.A(_1227_),
    .X(net849));
 sg13g2_buf_8 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net855),
    .X(net851));
 sg13g2_buf_8 fanout852 (.A(net855),
    .X(net852));
 sg13g2_buf_8 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_8 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_8 fanout855 (.A(_1004_),
    .X(net855));
 sg13g2_buf_8 fanout856 (.A(net867),
    .X(net856));
 sg13g2_buf_1 fanout857 (.A(net867),
    .X(net857));
 sg13g2_buf_8 fanout858 (.A(net867),
    .X(net858));
 sg13g2_buf_1 fanout859 (.A(net867),
    .X(net859));
 sg13g2_buf_8 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_8 fanout861 (.A(net866),
    .X(net861));
 sg13g2_buf_8 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_8 fanout863 (.A(net866),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_1 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_8 fanout867 (.A(_0971_),
    .X(net867));
 sg13g2_buf_8 fanout868 (.A(_1953_),
    .X(net868));
 sg13g2_buf_1 fanout869 (.A(_1953_),
    .X(net869));
 sg13g2_buf_8 fanout870 (.A(_1918_),
    .X(net870));
 sg13g2_buf_8 fanout871 (.A(net873),
    .X(net871));
 sg13g2_buf_8 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_8 fanout873 (.A(_1419_),
    .X(net873));
 sg13g2_buf_8 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_8 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_8 fanout876 (.A(_1103_),
    .X(net876));
 sg13g2_buf_8 fanout877 (.A(_3532_),
    .X(net877));
 sg13g2_buf_8 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_8 fanout879 (.A(_3532_),
    .X(net879));
 sg13g2_buf_8 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_8 fanout881 (.A(net885),
    .X(net881));
 sg13g2_buf_8 fanout882 (.A(net884),
    .X(net882));
 sg13g2_buf_1 fanout883 (.A(net884),
    .X(net883));
 sg13g2_buf_8 fanout884 (.A(net885),
    .X(net884));
 sg13g2_buf_8 fanout885 (.A(_3493_),
    .X(net885));
 sg13g2_buf_8 fanout886 (.A(net889),
    .X(net886));
 sg13g2_buf_8 fanout887 (.A(net889),
    .X(net887));
 sg13g2_buf_8 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_8 fanout889 (.A(_3424_),
    .X(net889));
 sg13g2_buf_8 fanout890 (.A(net891),
    .X(net890));
 sg13g2_buf_8 fanout891 (.A(_3411_),
    .X(net891));
 sg13g2_buf_8 fanout892 (.A(net894),
    .X(net892));
 sg13g2_buf_8 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_8 fanout894 (.A(_1861_),
    .X(net894));
 sg13g2_buf_8 fanout895 (.A(_1785_),
    .X(net895));
 sg13g2_buf_8 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(net901),
    .X(net897));
 sg13g2_buf_8 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_8 fanout899 (.A(net901),
    .X(net899));
 sg13g2_buf_1 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_8 fanout901 (.A(_1529_),
    .X(net901));
 sg13g2_buf_8 fanout902 (.A(net903),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net907),
    .X(net903));
 sg13g2_buf_8 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_8 fanout905 (.A(net907),
    .X(net905));
 sg13g2_buf_1 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_8 fanout907 (.A(_1528_),
    .X(net907));
 sg13g2_buf_8 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_8 fanout909 (.A(_1526_),
    .X(net909));
 sg13g2_buf_8 fanout910 (.A(net912),
    .X(net910));
 sg13g2_buf_1 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_8 fanout912 (.A(_1526_),
    .X(net912));
 sg13g2_buf_8 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(_1418_),
    .X(net914));
 sg13g2_buf_8 fanout915 (.A(_1346_),
    .X(net915));
 sg13g2_buf_8 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_8 fanout917 (.A(_1123_),
    .X(net917));
 sg13g2_buf_8 fanout918 (.A(net920),
    .X(net918));
 sg13g2_buf_1 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_8 fanout920 (.A(_1121_),
    .X(net920));
 sg13g2_buf_8 fanout921 (.A(net923),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(net923),
    .X(net922));
 sg13g2_buf_8 fanout923 (.A(_1118_),
    .X(net923));
 sg13g2_buf_8 fanout924 (.A(_1117_),
    .X(net924));
 sg13g2_buf_8 fanout925 (.A(_1117_),
    .X(net925));
 sg13g2_buf_8 fanout926 (.A(net928),
    .X(net926));
 sg13g2_buf_1 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_8 fanout928 (.A(_1115_),
    .X(net928));
 sg13g2_buf_8 fanout929 (.A(net930),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(_1113_),
    .X(net930));
 sg13g2_buf_8 fanout931 (.A(net933),
    .X(net931));
 sg13g2_buf_1 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_8 fanout933 (.A(_1111_),
    .X(net933));
 sg13g2_buf_8 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_8 fanout935 (.A(net936),
    .X(net935));
 sg13g2_buf_8 fanout936 (.A(_1109_),
    .X(net936));
 sg13g2_buf_8 fanout937 (.A(net938),
    .X(net937));
 sg13g2_buf_1 fanout938 (.A(_1045_),
    .X(net938));
 sg13g2_buf_8 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_8 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_8 fanout941 (.A(net943),
    .X(net941));
 sg13g2_buf_8 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_1045_),
    .X(net943));
 sg13g2_buf_8 fanout944 (.A(net947),
    .X(net944));
 sg13g2_buf_8 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_8 fanout946 (.A(net947),
    .X(net946));
 sg13g2_buf_8 fanout947 (.A(_1045_),
    .X(net947));
 sg13g2_buf_8 fanout948 (.A(_1044_),
    .X(net948));
 sg13g2_buf_1 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_8 fanout950 (.A(_1044_),
    .X(net950));
 sg13g2_buf_8 fanout951 (.A(_1016_),
    .X(net951));
 sg13g2_buf_8 fanout952 (.A(_3574_),
    .X(net952));
 sg13g2_buf_1 fanout953 (.A(_3574_),
    .X(net953));
 sg13g2_buf_8 fanout954 (.A(_3264_),
    .X(net954));
 sg13g2_buf_8 fanout955 (.A(_3259_),
    .X(net955));
 sg13g2_buf_8 fanout956 (.A(_2769_),
    .X(net956));
 sg13g2_buf_8 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_8 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_8 fanout959 (.A(net965),
    .X(net959));
 sg13g2_buf_8 fanout960 (.A(net965),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net965),
    .X(net961));
 sg13g2_buf_8 fanout962 (.A(net964),
    .X(net962));
 sg13g2_buf_1 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_8 fanout964 (.A(net965),
    .X(net964));
 sg13g2_buf_8 fanout965 (.A(_2769_),
    .X(net965));
 sg13g2_buf_8 fanout966 (.A(_1774_),
    .X(net966));
 sg13g2_buf_8 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_8 fanout968 (.A(_1773_),
    .X(net968));
 sg13g2_buf_8 fanout969 (.A(_3236_),
    .X(net969));
 sg13g2_buf_8 fanout970 (.A(_2613_),
    .X(net970));
 sg13g2_buf_1 fanout971 (.A(_2613_),
    .X(net971));
 sg13g2_buf_8 fanout972 (.A(_2252_),
    .X(net972));
 sg13g2_buf_8 fanout973 (.A(net974),
    .X(net973));
 sg13g2_buf_8 fanout974 (.A(_2250_),
    .X(net974));
 sg13g2_buf_8 fanout975 (.A(net977),
    .X(net975));
 sg13g2_buf_1 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_8 fanout977 (.A(_2180_),
    .X(net977));
 sg13g2_buf_8 fanout978 (.A(net980),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(net980),
    .X(net979));
 sg13g2_buf_8 fanout980 (.A(_2179_),
    .X(net980));
 sg13g2_buf_8 fanout981 (.A(net982),
    .X(net981));
 sg13g2_buf_8 fanout982 (.A(_1822_),
    .X(net982));
 sg13g2_buf_8 fanout983 (.A(_0980_),
    .X(net983));
 sg13g2_buf_8 fanout984 (.A(_0980_),
    .X(net984));
 sg13g2_buf_8 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_8 fanout986 (.A(_0914_),
    .X(net986));
 sg13g2_buf_8 fanout987 (.A(net988),
    .X(net987));
 sg13g2_buf_8 fanout988 (.A(_0914_),
    .X(net988));
 sg13g2_buf_8 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_8 fanout990 (.A(_0914_),
    .X(net990));
 sg13g2_buf_8 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_8 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_8 fanout993 (.A(net1001),
    .X(net993));
 sg13g2_buf_8 fanout994 (.A(net995),
    .X(net994));
 sg13g2_buf_8 fanout995 (.A(net1001),
    .X(net995));
 sg13g2_buf_8 fanout996 (.A(net1000),
    .X(net996));
 sg13g2_buf_8 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_1 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_8 fanout999 (.A(net1000),
    .X(net999));
 sg13g2_buf_8 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_8 fanout1001 (.A(_0912_),
    .X(net1001));
 sg13g2_buf_8 fanout1002 (.A(_3475_),
    .X(net1002));
 sg13g2_buf_8 fanout1003 (.A(_3457_),
    .X(net1003));
 sg13g2_buf_8 fanout1004 (.A(_3255_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_3255_),
    .X(net1005));
 sg13g2_buf_8 fanout1006 (.A(net1009),
    .X(net1006));
 sg13g2_buf_8 fanout1007 (.A(net1008),
    .X(net1007));
 sg13g2_buf_8 fanout1008 (.A(net1009),
    .X(net1008));
 sg13g2_buf_8 fanout1009 (.A(_3241_),
    .X(net1009));
 sg13g2_buf_8 fanout1010 (.A(_3235_),
    .X(net1010));
 sg13g2_buf_8 fanout1011 (.A(_3191_),
    .X(net1011));
 sg13g2_buf_8 fanout1012 (.A(net1013),
    .X(net1012));
 sg13g2_buf_1 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_1 fanout1014 (.A(_2886_),
    .X(net1014));
 sg13g2_buf_8 fanout1015 (.A(_2873_),
    .X(net1015));
 sg13g2_buf_8 fanout1016 (.A(_2873_),
    .X(net1016));
 sg13g2_buf_8 fanout1017 (.A(net1019),
    .X(net1017));
 sg13g2_buf_8 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_8 fanout1019 (.A(_2450_),
    .X(net1019));
 sg13g2_buf_8 fanout1020 (.A(_1511_),
    .X(net1020));
 sg13g2_buf_8 fanout1021 (.A(net1784),
    .X(net1021));
 sg13g2_buf_1 fanout1022 (.A(net1784),
    .X(net1022));
 sg13g2_buf_8 fanout1023 (.A(net1025),
    .X(net1023));
 sg13g2_buf_1 fanout1024 (.A(net1025),
    .X(net1024));
 sg13g2_buf_8 fanout1025 (.A(net1030),
    .X(net1025));
 sg13g2_buf_8 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_8 fanout1027 (.A(net1030),
    .X(net1027));
 sg13g2_buf_8 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_8 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_8 fanout1030 (.A(net1042),
    .X(net1030));
 sg13g2_buf_8 fanout1031 (.A(net1033),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(net1036),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1036),
    .X(net1033));
 sg13g2_buf_8 fanout1034 (.A(net1036),
    .X(net1034));
 sg13g2_buf_1 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_8 fanout1036 (.A(net1042),
    .X(net1036));
 sg13g2_buf_8 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_8 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_8 fanout1039 (.A(net1042),
    .X(net1039));
 sg13g2_buf_8 fanout1040 (.A(net1041),
    .X(net1040));
 sg13g2_buf_8 fanout1041 (.A(net1042),
    .X(net1041));
 sg13g2_buf_8 fanout1042 (.A(_0905_),
    .X(net1042));
 sg13g2_buf_8 fanout1043 (.A(net1045),
    .X(net1043));
 sg13g2_buf_1 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_8 fanout1045 (.A(net1058),
    .X(net1045));
 sg13g2_buf_8 fanout1046 (.A(net1047),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1049),
    .X(net1047));
 sg13g2_buf_8 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_1 fanout1049 (.A(net1058),
    .X(net1049));
 sg13g2_buf_8 fanout1050 (.A(net1052),
    .X(net1050));
 sg13g2_buf_1 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_1 fanout1053 (.A(net1057),
    .X(net1053));
 sg13g2_buf_8 fanout1054 (.A(net1056),
    .X(net1054));
 sg13g2_buf_1 fanout1055 (.A(net1056),
    .X(net1055));
 sg13g2_buf_8 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_1 fanout1057 (.A(net1058),
    .X(net1057));
 sg13g2_buf_8 fanout1058 (.A(_0904_),
    .X(net1058));
 sg13g2_buf_8 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_8 fanout1060 (.A(_0904_),
    .X(net1060));
 sg13g2_buf_8 fanout1061 (.A(_3245_),
    .X(net1061));
 sg13g2_buf_8 fanout1062 (.A(_3242_),
    .X(net1062));
 sg13g2_buf_8 fanout1063 (.A(net1064),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_3239_),
    .X(net1064));
 sg13g2_buf_8 fanout1065 (.A(net1066),
    .X(net1065));
 sg13g2_buf_8 fanout1066 (.A(_3239_),
    .X(net1066));
 sg13g2_buf_8 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_8 fanout1068 (.A(_3223_),
    .X(net1068));
 sg13g2_buf_8 fanout1069 (.A(net1070),
    .X(net1069));
 sg13g2_buf_8 fanout1070 (.A(_3223_),
    .X(net1070));
 sg13g2_buf_8 fanout1071 (.A(net1075),
    .X(net1071));
 sg13g2_buf_8 fanout1072 (.A(net1075),
    .X(net1072));
 sg13g2_buf_8 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_8 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_8 fanout1075 (.A(_3220_),
    .X(net1075));
 sg13g2_buf_8 fanout1076 (.A(_2882_),
    .X(net1076));
 sg13g2_buf_8 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_8 fanout1078 (.A(_2876_),
    .X(net1078));
 sg13g2_buf_8 fanout1079 (.A(net1081),
    .X(net1079));
 sg13g2_buf_8 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_8 fanout1081 (.A(_2876_),
    .X(net1081));
 sg13g2_buf_8 fanout1082 (.A(_2872_),
    .X(net1082));
 sg13g2_buf_8 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_8 fanout1084 (.A(_2845_),
    .X(net1084));
 sg13g2_buf_8 fanout1085 (.A(net1087),
    .X(net1085));
 sg13g2_buf_8 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_8 fanout1087 (.A(_2845_),
    .X(net1087));
 sg13g2_buf_8 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_8 fanout1089 (.A(_2844_),
    .X(net1089));
 sg13g2_buf_8 fanout1090 (.A(net1092),
    .X(net1090));
 sg13g2_buf_8 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_8 fanout1092 (.A(_2844_),
    .X(net1092));
 sg13g2_buf_8 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_8 fanout1094 (.A(_2526_),
    .X(net1094));
 sg13g2_buf_8 fanout1095 (.A(_2451_),
    .X(net1095));
 sg13g2_buf_8 fanout1096 (.A(_1520_),
    .X(net1096));
 sg13g2_buf_8 fanout1097 (.A(_1506_),
    .X(net1097));
 sg13g2_buf_8 fanout1098 (.A(_0916_),
    .X(net1098));
 sg13g2_buf_8 fanout1099 (.A(net1102),
    .X(net1099));
 sg13g2_buf_8 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_8 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_8 fanout1102 (.A(_0894_),
    .X(net1102));
 sg13g2_buf_8 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_8 fanout1104 (.A(net1105),
    .X(net1104));
 sg13g2_buf_8 fanout1105 (.A(net1109),
    .X(net1105));
 sg13g2_buf_8 fanout1106 (.A(net1108),
    .X(net1106));
 sg13g2_buf_1 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_8 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(net1132),
    .X(net1109));
 sg13g2_buf_8 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_buf_8 fanout1111 (.A(net1117),
    .X(net1111));
 sg13g2_buf_8 fanout1112 (.A(net1116),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(net1116),
    .X(net1113));
 sg13g2_buf_8 fanout1114 (.A(net1116),
    .X(net1114));
 sg13g2_buf_1 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(net1132),
    .X(net1117));
 sg13g2_buf_8 fanout1118 (.A(net1120),
    .X(net1118));
 sg13g2_buf_8 fanout1119 (.A(net1120),
    .X(net1119));
 sg13g2_buf_8 fanout1120 (.A(net1122),
    .X(net1120));
 sg13g2_buf_8 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_8 fanout1122 (.A(net1132),
    .X(net1122));
 sg13g2_buf_8 fanout1123 (.A(net1127),
    .X(net1123));
 sg13g2_buf_8 fanout1124 (.A(net1127),
    .X(net1124));
 sg13g2_buf_8 fanout1125 (.A(net1126),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(net1127),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(net1132),
    .X(net1127));
 sg13g2_buf_8 fanout1128 (.A(net1131),
    .X(net1128));
 sg13g2_buf_8 fanout1129 (.A(net1131),
    .X(net1129));
 sg13g2_buf_1 fanout1130 (.A(net1131),
    .X(net1130));
 sg13g2_buf_8 fanout1131 (.A(net1132),
    .X(net1131));
 sg13g2_buf_8 fanout1132 (.A(_0884_),
    .X(net1132));
 sg13g2_buf_8 fanout1133 (.A(_0756_),
    .X(net1133));
 sg13g2_buf_8 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_8 fanout1135 (.A(_0755_),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_8 fanout1137 (.A(\led_controller.register_address[3] ),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_1 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(\led_controller.register_address[2] ),
    .X(net1141));
 sg13g2_buf_8 fanout1142 (.A(net1143),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(net1613),
    .X(net1143));
 sg13g2_buf_8 fanout1144 (.A(net1149),
    .X(net1144));
 sg13g2_buf_1 fanout1145 (.A(net1149),
    .X(net1145));
 sg13g2_buf_8 fanout1146 (.A(net1148),
    .X(net1146));
 sg13g2_buf_8 fanout1147 (.A(net1149),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_8 fanout1149 (.A(net1162),
    .X(net1149));
 sg13g2_buf_8 fanout1150 (.A(net1151),
    .X(net1150));
 sg13g2_buf_8 fanout1151 (.A(net1154),
    .X(net1151));
 sg13g2_buf_8 fanout1152 (.A(net1154),
    .X(net1152));
 sg13g2_buf_8 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_8 fanout1154 (.A(net1162),
    .X(net1154));
 sg13g2_buf_8 fanout1155 (.A(net1156),
    .X(net1155));
 sg13g2_buf_8 fanout1156 (.A(net1162),
    .X(net1156));
 sg13g2_buf_8 fanout1157 (.A(net1158),
    .X(net1157));
 sg13g2_buf_8 fanout1158 (.A(net1161),
    .X(net1158));
 sg13g2_buf_8 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_8 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_8 fanout1162 (.A(net2015),
    .X(net1162));
 sg13g2_buf_8 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_8 fanout1164 (.A(\led_controller.led_effect_pulse.color_1.counter[1] ),
    .X(net1164));
 sg13g2_buf_8 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_8 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_8 fanout1167 (.A(net2383),
    .X(net1167));
 sg13g2_buf_8 fanout1168 (.A(net2277),
    .X(net1168));
 sg13g2_buf_1 fanout1169 (.A(\led_controller.led_effect_pulse.brightness[4] ),
    .X(net1169));
 sg13g2_buf_8 fanout1170 (.A(net2336),
    .X(net1170));
 sg13g2_buf_1 fanout1171 (.A(\led_controller.led_effect_pulse.brightness[3] ),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(net2281),
    .X(net1172));
 sg13g2_buf_1 fanout1173 (.A(\led_controller.led_effect_pulse.brightness[2] ),
    .X(net1173));
 sg13g2_buf_8 fanout1174 (.A(net2372),
    .X(net1174));
 sg13g2_buf_8 fanout1175 (.A(net2365),
    .X(net1175));
 sg13g2_buf_8 fanout1176 (.A(net1608),
    .X(net1176));
 sg13g2_buf_8 fanout1177 (.A(net1178),
    .X(net1177));
 sg13g2_buf_8 fanout1178 (.A(net2382),
    .X(net1178));
 sg13g2_buf_8 fanout1179 (.A(net2371),
    .X(net1179));
 sg13g2_buf_8 fanout1180 (.A(net2356),
    .X(net1180));
 sg13g2_buf_8 fanout1181 (.A(net2378),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(net2368),
    .X(net1182));
 sg13g2_buf_8 fanout1183 (.A(net2377),
    .X(net1183));
 sg13g2_buf_8 fanout1184 (.A(net2362),
    .X(net1184));
 sg13g2_buf_8 fanout1185 (.A(\led_controller.cpu.register_x[0] ),
    .X(net1185));
 sg13g2_buf_8 fanout1186 (.A(net2381),
    .X(net1186));
 sg13g2_buf_8 fanout1187 (.A(net1188),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(\led_controller.led_effect_pulse.color_1.active ),
    .X(net1188));
 sg13g2_buf_8 fanout1189 (.A(net2376),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(net2333),
    .X(net1190));
 sg13g2_buf_8 fanout1191 (.A(net2353),
    .X(net1191));
 sg13g2_buf_8 fanout1192 (.A(net2087),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(net1936),
    .X(net1193));
 sg13g2_buf_8 fanout1194 (.A(net2374),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(_0003_),
    .X(net1195));
 sg13g2_buf_8 fanout1196 (.A(_0002_),
    .X(net1196));
 sg13g2_buf_8 fanout1197 (.A(net1199),
    .X(net1197));
 sg13g2_buf_1 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_8 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_8 fanout1200 (.A(_0001_),
    .X(net1200));
 sg13g2_buf_8 fanout1201 (.A(net1202),
    .X(net1201));
 sg13g2_buf_8 fanout1202 (.A(net1205),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(net1205),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(net1205),
    .X(net1204));
 sg13g2_buf_8 fanout1205 (.A(_0001_),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(net1223),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(net1223),
    .X(net1207));
 sg13g2_buf_8 fanout1208 (.A(net1210),
    .X(net1208));
 sg13g2_buf_1 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(net1223),
    .X(net1210));
 sg13g2_buf_8 fanout1211 (.A(net1214),
    .X(net1211));
 sg13g2_buf_1 fanout1212 (.A(net1214),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(net1214),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(net1222),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(net1222),
    .X(net1215));
 sg13g2_buf_1 fanout1216 (.A(net1222),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(net1221),
    .X(net1217));
 sg13g2_buf_1 fanout1218 (.A(net1221),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(net1221),
    .X(net1219));
 sg13g2_buf_1 fanout1220 (.A(net1221),
    .X(net1220));
 sg13g2_buf_1 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_8 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_8 fanout1223 (.A(_0000_),
    .X(net1223));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_tielo tt_um_chrismoos_led_controller_6 (.L_LO(net6));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_91_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_92_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\led_controller.reset.reset1 ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold2 (.A(\led_controller.spi_slave.sync_ss_n.data ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold3 (.A(\led_controller.spi_slave.sync_mosi.data ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold4 (.A(\led_controller.spi_slave.sync_sck.data ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold5 (.A(\led_controller.flash.cs_delay_counter[0] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0436_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold7 (.A(\led_controller.cpu.scratch_memory[6][4] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold8 (.A(\led_controller.cpu.scratch_memory[10][2] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0050_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold10 (.A(\led_controller.cpu.scratch_memory[6][5] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold11 (.A(\led_controller.cpu.scratch_memory[6][2] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold12 (.A(\led_controller.cpu.scratch_memory[6][7] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold13 (.A(\led_controller.cpu.scratch_memory[2][5] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold14 (.A(\led_controller.cpu.scratch_memory[10][7] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0055_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold16 (.A(\led_controller.cpu.scratch_memory[14][4] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold17 (.A(\led_controller.cpu.scratch_memory[6][3] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold18 (.A(\led_controller.cpu.scratch_memory[10][3] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0051_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold20 (.A(\led_controller.cpu.scratch_memory[6][0] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold21 (.A(\led_controller.cpu.scratch_memory[14][3] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold22 (.A(\led_controller.spi_slave.output_register[4] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0154_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold24 (.A(\led_controller.spi_slave.sck ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold25 (.A(\led_controller.cpu.scratch_memory[12][1] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold26 (.A(\led_controller.rgbw.counter[0] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0127_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold28 (.A(\led_controller.cpu.scratch_memory[14][7] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold29 (.A(\led_controller.cpu.scratch_memory[4][0] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold30 (.A(\led_controller.cpu.scratch_memory[7][2] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold31 (.A(\led_controller.cpu.scratch_memory[15][0] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold32 (.A(\led_controller.cpu.scratch_memory[6][6] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold33 (.A(\led_controller.cpu.scratch_memory[2][6] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold34 (.A(\led_controller.cpu.scratch_memory[9][7] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0039_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold36 (.A(\led_controller.cpu.scratch_memory[4][6] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold37 (.A(\led_controller.cpu.scratch_memory[10][6] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0054_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold39 (.A(\led_controller.cpu.scratch_memory[5][5] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold40 (.A(\led_controller.cpu.scratch_memory[0][2] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold41 (.A(\led_controller.cpu.scratch_memory[9][2] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0034_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold43 (.A(\led_controller.cpu.scratch_memory[14][1] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold44 (.A(\led_controller.cpu.scratch_memory[11][2] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0042_),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold46 (.A(\led_controller.cpu.scratch_memory[7][3] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold47 (.A(\led_controller.cpu.scratch_memory[10][0] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0048_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold49 (.A(\led_controller.cpu.scratch_memory[7][6] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0480_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold51 (.A(\led_controller.cpu.scratch_memory[1][4] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold52 (.A(\led_controller.cpu.scratch_memory[12][5] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold53 (.A(\led_controller.cpu.scratch_memory[11][4] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0044_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold55 (.A(\led_controller.cpu.scratch_memory[13][3] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold56 (.A(\led_controller.cpu.scratch_memory[6][1] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold57 (.A(\led_controller.cpu.scratch_memory[1][0] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold58 (.A(\led_controller.cpu.scratch_memory[0][7] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold59 (.A(\led_controller.cpu.scratch_memory[7][7] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold60 (.A(\led_controller.cpu.scratch_memory[4][3] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold61 (.A(\led_controller.cpu.scratch_memory[0][0] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold62 (.A(\led_controller.cpu.scratch_memory[15][7] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold63 (.A(\led_controller.cpu.scratch_memory[0][3] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold64 (.A(\led_controller.cpu.scratch_memory[11][1] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0041_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold66 (.A(\led_controller.cpu.scratch_memory[12][0] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold67 (.A(\led_controller.cpu.scratch_memory[0][6] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold68 (.A(\led_controller.cpu.scratch_memory[2][4] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold69 (.A(\led_controller.cpu.scratch_memory[8][7] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0739_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold71 (.A(\led_controller.spi_slave.output_register[1] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0151_),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold73 (.A(\led_controller.cpu.scratch_memory[1][6] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold74 (.A(\led_controller.led_effect_pulse.calc_color_out[8] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold75 (.A(\led_controller.cpu.scratch_memory[1][3] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold76 (.A(\led_controller.cpu.scratch_memory[5][6] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold77 (.A(\led_controller.cpu.scratch_memory[9][1] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0033_),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold79 (.A(\led_controller.cpu.scratch_memory[9][3] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0035_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold81 (.A(\led_controller.cpu.scratch_memory[8][1] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0733_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold83 (.A(\led_controller.cpu.scratch_memory[1][2] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold84 (.A(\led_controller.cpu.scratch_memory[13][4] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold85 (.A(\led_controller.cpu.scratch_memory[15][1] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold86 (.A(\led_controller.cpu.scratch_memory[2][3] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold87 (.A(\led_controller.cpu.scratch_memory[1][5] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold88 (.A(\led_controller.cpu.scratch_memory[9][5] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0037_),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold90 (.A(\led_controller.cpu.scratch_memory[7][1] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold91 (.A(\led_controller.cpu.scratch_memory[13][2] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold92 (.A(\led_controller.cpu.scratch_memory[5][1] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold93 (.A(\led_controller.cpu.scratch_memory[4][2] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold94 (.A(\led_controller.cpu.scratch_memory[8][5] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0737_),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold96 (.A(\led_controller.cpu.scratch_memory[8][4] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0736_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold98 (.A(\led_controller.cpu.scratch_memory[12][6] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold99 (.A(\led_controller.cpu.scratch_memory[0][5] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold100 (.A(\led_controller.cpu.scratch_memory[4][7] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold101 (.A(\led_controller.cpu.scratch_memory[11][3] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0043_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold103 (.A(\led_controller.flash.master.o_mosi ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0444_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold105 (.A(\led_controller.cpu.scratch_memory[12][3] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold106 (.A(\led_controller.cpu.scratch_memory[8][2] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0734_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold108 (.A(\led_controller.cpu.scratch_memory[3][4] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold109 (.A(\led_controller.cpu.scratch_memory[5][3] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold110 (.A(\led_controller.cpu.scratch_memory[13][5] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold111 (.A(\led_controller.cpu.scratch_memory[3][6] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold112 (.A(\led_controller.cpu.scratch_memory[14][0] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold113 (.A(\led_controller.cpu.scratch_memory[4][4] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold114 (.A(\led_controller.cpu.scratch_memory[2][1] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold115 (.A(\led_controller.cpu.scratch_memory[8][3] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0735_),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold117 (.A(\led_controller.cpu.scratch_memory[1][7] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold118 (.A(\led_controller.timer_100hz.div_counter[0] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold119 (.A(\led_controller.cpu.scratch_memory[1][1] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold120 (.A(\led_controller.cpu.scratch_memory[5][7] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold121 (.A(\led_controller.cpu.scratch_memory[13][7] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold122 (.A(\led_controller.cpu.scratch_memory[9][4] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0036_),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold124 (.A(\led_controller.cpu.scratch_memory[0][1] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold125 (.A(\led_controller.cpu.scratch_memory[12][7] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold126 (.A(\led_controller.cpu.scratch_memory[7][0] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold127 (.A(\led_controller.cpu.scratch_memory[7][5] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold128 (.A(\led_controller.cpu.scratch_memory[9][6] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0038_),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold130 (.A(\led_controller.cpu.scratch_memory[14][6] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold131 (.A(\led_controller.cpu.scratch_memory[15][5] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold132 (.A(\led_controller.led_effect_pulse.calc_color_out[12] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold133 (.A(\led_controller.cpu.scratch_memory[13][1] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0447_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold135 (.A(\led_controller.cpu.scratch_memory[11][0] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0040_),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold137 (.A(\led_controller.cpu.scratch_memory[3][3] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold138 (.A(\led_controller.cpu.scratch_memory[5][4] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold139 (.A(\led_controller.cpu.scratch_memory[11][7] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0047_),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold141 (.A(\led_controller.cpu.scratch_memory[8][0] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0732_),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold143 (.A(\led_controller.cpu.scratch_memory[15][6] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold144 (.A(\led_controller.timer_100hz.counter[30] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0205_),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold146 (.A(\led_controller.cpu.scratch_memory[4][5] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold147 (.A(\led_controller.cpu.scratch_memory[2][7] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold148 (.A(\led_controller.cpu.scratch_memory[9][0] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0032_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold150 (.A(\led_controller.spi_slave.output_register[3] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0153_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold152 (.A(\led_controller.cpu.scratch_memory[7][4] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold153 (.A(\led_controller.cpu.scratch_memory[8][6] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0738_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold155 (.A(\led_controller.cpu.scratch_memory[5][0] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold156 (.A(\led_controller.cpu.scratch_memory[13][6] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold157 (.A(\led_controller.cpu.scratch_memory[13][0] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold158 (.A(\led_controller.led_effect_pulse.calc_color_out[11] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold159 (.A(\led_controller.flash.addr[14] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0403_),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold161 (.A(\led_controller.cpu.scratch_memory[15][2] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold162 (.A(\led_controller.cpu.scratch_memory[3][5] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold163 (.A(\led_controller.flash.addr[11] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0400_),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold165 (.A(\led_controller.cpu.scratch_memory[10][1] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0049_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold167 (.A(\led_controller.flash.addr[12] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0401_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold169 (.A(\led_controller.cpu.scratch_memory[10][4] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0052_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold171 (.A(\led_controller.flash.master.sck ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0457_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold173 (.A(\led_controller.spi_slave.output_register[6] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0156_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold175 (.A(\led_controller.cpu.scratch_memory[5][2] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold176 (.A(\led_controller.cpu.scratch_memory[3][7] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold177 (.A(\led_controller.cpu.current_instruction[13] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0364_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold179 (.A(\led_controller.cpu.scratch_memory[4][1] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold180 (.A(\led_controller.cpu.scratch_memory[0][4] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold181 (.A(\led_controller.flash.addr[8] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0397_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold183 (.A(\led_controller.cpu.current_instruction[15] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0366_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold185 (.A(\led_controller.cpu.scratch_memory[3][0] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0080_),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold187 (.A(\led_controller.cpu.scratch_memory[12][2] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold188 (.A(\led_controller.cpu.scratch_memory[2][0] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold189 (.A(\led_controller.spi_slave.output_register[2] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0152_),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold191 (.A(\led_controller.flash.state[3] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0413_),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold193 (.A(\led_controller.led_effect_pulse.calc_color_out[14] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold194 (.A(\led_controller.flash.addr[13] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0402_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold196 (.A(\led_controller.led_effect_pulse.calc_color_out[15] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold197 (.A(\led_controller.cpu.current_instruction[14] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0365_),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold199 (.A(\led_controller.cpu.scratch_memory[11][5] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0045_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold201 (.A(\led_controller.cpu.scratch_memory[2][2] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold202 (.A(\led_controller.cpu.scratch_memory[11][6] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0046_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold204 (.A(\led_controller.effect_pulse_led_color[21] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0504_),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold206 (.A(\led_controller.effect_pulse_led_color[7] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0490_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold208 (.A(\led_controller.flash.addr[7] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0396_),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold210 (.A(\led_controller.cpu.scratch_memory[12][4] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold211 (.A(\led_controller.cpu.fetch_instruction[13] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0348_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold213 (.A(\led_controller.effect_pulse_led_color[20] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0503_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold215 (.A(\led_controller.cpu.scratch_memory[3][2] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold216 (.A(\led_controller.flash.addr[10] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0399_),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold218 (.A(\led_controller.led_effect_pulse.state[1] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0012_),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold220 (.A(\led_controller.flash.addr[5] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0394_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold222 (.A(\led_controller.flash.addr[9] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0398_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold224 (.A(\led_controller.cpu.scratch_memory[15][4] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold225 (.A(\led_controller.cpu.scratch_memory[10][5] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0053_),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold227 (.A(\led_controller.flash.addr[15] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0404_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold229 (.A(\led_controller.effect_pulse_led_color[22] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0505_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold231 (.A(\led_controller.spi_slave.output_register[5] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0155_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold233 (.A(\led_controller.cpu.scratch_memory[3][1] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold234 (.A(\led_controller.effect_pulse_led_color[2] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0485_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold236 (.A(\led_controller.flash.addr[6] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0395_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold238 (.A(\led_controller.flash.addr[1] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0390_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold240 (.A(\led_controller.effect_pulse_led_color[23] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0506_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold242 (.A(\led_controller.cpu.scratch_memory[14][2] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold243 (.A(\led_controller.timer_2hz.counter[1] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold244 (.A(_1386_),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0165_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold246 (.A(\led_controller.o_data ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold247 (.A(_1493_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0216_),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold249 (.A(\led_controller.led_effect_pulse.calc_color_out[13] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold250 (.A(\led_controller.effect_pulse_led_color[3] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0486_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold252 (.A(\led_controller.effect_pulse_led_color[30] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0513_),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold254 (.A(\led_controller.cpu.fetch_instruction[14] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0349_),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold256 (.A(\led_controller.cpu.fetch_instruction[15] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0350_),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold258 (.A(\led_controller.effect_pulse_led_color[9] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0492_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold260 (.A(\led_controller.effect_pulse_led_color[4] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0487_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold262 (.A(\led_controller.effect_pulse_led_color[5] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0488_),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold264 (.A(\led_controller.effect_pulse_led_color[0] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0483_),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold266 (.A(\led_controller.spi_slave.output_register[0] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0150_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold268 (.A(\led_controller.flash.addr[4] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0393_),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold270 (.A(\led_controller.effect_pulse_led_color[6] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0489_),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold272 (.A(\led_controller.cpu.current_instruction_valid ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold273 (.A(\led_controller.cpu.o_led_color[1] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0279_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold275 (.A(\led_controller.flash.addr[0] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0389_),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold277 (.A(\led_controller.led_effect_pulse.calc_color_out[5] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold278 (.A(\led_controller.cpu.fetch_instruction[11] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0346_),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold280 (.A(\led_controller.effect_pulse_led_color[11] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold281 (.A(\led_controller.cpu.current_instruction[6] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0357_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold283 (.A(\led_controller.cpu.current_instruction_pc[15] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0382_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold285 (.A(\led_controller.effect_pulse_led_color[10] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0493_),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold287 (.A(\led_controller.cpu.current_instruction_pc[13] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0380_),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold289 (.A(\led_controller.cpu.current_instruction_pc[3] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0370_),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold291 (.A(\led_controller.cpu.fetch_instruction[9] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0344_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold293 (.A(\led_controller.timer_100hz.counter[9] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0184_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold295 (.A(\led_controller.effect_pulse_led_color[26] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0509_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold297 (.A(\led_controller.cpu.fetch_instruction[10] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0345_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold299 (.A(\led_controller.cpu.current_instruction_pc[10] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0377_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold301 (.A(\led_controller.led_effect_pulse.calc_color_out[6] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold302 (.A(\led_controller.led_effect_pulse.calc_color_out[18] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0551_),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold304 (.A(\led_controller.effect_pulse_led_color[17] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0500_),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold306 (.A(\led_controller.effect_pulse_led_color[19] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0502_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold308 (.A(\led_controller.spi_slave.last_ss ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold309 (.A(_1329_),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold310 (.A(\led_controller.effect_pulse_led_color[29] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0512_),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold312 (.A(\led_controller.flash.addr[2] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0391_),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold314 (.A(\led_controller.cpu.current_instruction_pc[12] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0379_),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold316 (.A(\led_controller.cpu.o_led_color[0] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0278_),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold318 (.A(\led_controller.effect_pulse_led_color[13] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold319 (.A(\led_controller.effect_pulse_led_color[27] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0510_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold321 (.A(\led_controller.cpu.current_instruction_pc[2] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0369_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold323 (.A(\led_controller.cpu.current_instruction_pc[14] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0381_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold325 (.A(\led_controller.effect_pulse_led_color[16] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0499_),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold327 (.A(\led_controller.o_spi_miso ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0136_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold329 (.A(\led_controller.led_effect_pulse.calc_color_out[10] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold330 (.A(\led_controller.flash.addr[3] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0392_),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold332 (.A(\led_controller.spi_slave.data_bits[0] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0137_),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold334 (.A(\led_controller.cpu.current_instruction_pc[5] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0372_),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold336 (.A(\led_controller.spi_data_write[0] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0582_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold338 (.A(\led_controller.flash.state[2] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0998_),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0006_),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold341 (.A(\led_controller.cpu.current_instruction_pc[9] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0376_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold343 (.A(\led_controller.cpu.current_instruction_pc[8] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0375_),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold345 (.A(\led_controller.cpu.current_instruction[7] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0358_),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold347 (.A(\led_controller.effect_pulse_led_color[1] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0484_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold349 (.A(\led_controller.effect_pulse_led_color[8] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold350 (.A(\led_controller.effect_pulse_led_color[25] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0508_),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold352 (.A(\led_controller.timer_100hz.div_counter[2] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold353 (.A(_1185_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0066_),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold355 (.A(\led_controller.cpu.current_instruction_pc[11] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0378_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold357 (.A(\led_controller.flash.master.sck_counter[5] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold358 (.A(_2628_),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0422_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold360 (.A(\led_controller.flash.master.i_tx_data[0] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold361 (.A(_1779_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0270_),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold363 (.A(\led_controller.flash.master.sck_counter[2] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold364 (.A(_2622_),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0419_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold366 (.A(\led_controller.flash.state[5] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold367 (.A(_1005_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0007_),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold369 (.A(\led_controller.cpu.stall_counter[7] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0323_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold371 (.A(\led_controller.cpu.scratch_memory[14][5] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0029_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold373 (.A(\led_controller.effect_pulse_led_color[31] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0514_),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold375 (.A(\led_controller.cpu.o_bus_addr[13] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold376 (.A(_2514_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0339_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold378 (.A(\led_controller.led_effect_pulse.calc_color_out[4] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold379 (.A(\led_controller.cpu.fetch_instruction[12] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0347_),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold381 (.A(\led_controller.led_effect_chase.current_led[6] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold382 (.A(_2745_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0464_),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold384 (.A(\led_controller.timer_100hz.counter[31] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold385 (.A(_1480_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0206_),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold387 (.A(\led_controller.effect_pulse_led_color[24] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0507_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold389 (.A(\led_controller.cpu.current_instruction_pc[0] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0367_),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold391 (.A(\led_controller.cpu.current_instruction_pc[6] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0373_),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold393 (.A(\led_controller.flash.cs_delay_counter[2] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold394 (.A(_2648_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0438_),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold396 (.A(\led_controller.timer_10hz.counter[2] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold397 (.A(_1399_),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0172_),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold399 (.A(\led_controller.cpu.current_instruction_pc[4] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0371_),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold401 (.A(\led_controller.flash.master.sck_counter[0] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold402 (.A(_2620_),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0417_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold404 (.A(\led_controller.flash.cs_delay_counter[7] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0443_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold406 (.A(\led_controller.cpu_reset_counter[3] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold407 (.A(_3231_),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold408 (.A(\led_controller.effect_pulse_led_color[15] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold409 (.A(\led_controller.cpu.scratch_memory[15][3] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0469_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold411 (.A(\led_controller.cpu.fetch_instruction[8] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0343_),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold413 (.A(\led_controller.flash.state[0] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0996_),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0004_),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold416 (.A(\led_controller.led_effect_pulse.calc_color_out[26] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold417 (.A(_3196_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold418 (.A(\led_controller.led_effect_pulse.current_led[4] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold419 (.A(_2831_),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0520_),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold421 (.A(\led_controller.cpu_reset_counter[0] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold422 (.A(\led_controller.flash.master.i_tx_data[5] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold423 (.A(_1801_),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0275_),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold425 (.A(\led_controller.effect_pulse_led_color[18] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold426 (.A(\led_controller.rgbw.counter[2] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold427 (.A(_1319_),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0129_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold429 (.A(\led_controller.cpu.led_write_color[1] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold430 (.A(\led_controller.led_effect_pulse.current_led[3] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold431 (.A(_2829_),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0519_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold433 (.A(\led_controller.timer_100hz.counter[10] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold434 (.A(_1438_),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold435 (.A(\led_controller.cpu.current_instruction[5] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0356_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold437 (.A(\led_controller.effect_chase_led_strb ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold438 (.A(_2670_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0454_),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold440 (.A(\led_controller.cpu.o_bus_addr[10] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0336_),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold442 (.A(\led_controller.effect_pulse_led_color[12] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold443 (.A(\led_controller.flash.cs_delay_counter[6] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold444 (.A(_2652_),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0442_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold446 (.A(\led_controller.flash.master.o_busy ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0425_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold448 (.A(\led_controller.flash.master.i_tx_data[2] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0272_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold450 (.A(\led_controller.cpu.led_write_color[0] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold451 (.A(\led_controller.spi_data_write_strb ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold452 (.A(\led_controller.spi_data_write[7] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold453 (.A(_3369_),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold454 (.A(\led_controller.led_effect_pulse.calc_color_out[7] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold455 (.A(\led_controller.cpu.bus_hi_valid ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold456 (.A(_2571_),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold457 (.A(\led_controller.effect_pulse_led_color[28] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0511_),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold459 (.A(\led_controller.cpu.o_bus_addr[15] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold460 (.A(_2525_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0341_),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold462 (.A(\led_controller.cpu.current_instruction[4] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0355_),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold464 (.A(\led_controller.cpu.stall_counter[3] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0319_),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold466 (.A(\led_controller.cpu.i_bus_data[3] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0430_),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold468 (.A(\led_controller.timer_2hz.counter[2] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold469 (.A(_1388_),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0166_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold471 (.A(\led_controller.spi_data[6] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0604_),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold473 (.A(\led_controller.cpu.led_writing ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0280_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold475 (.A(\led_controller.rgbw.color[16] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold476 (.A(_1613_),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold477 (.A(\led_controller.rgbw.color[26] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold478 (.A(_1663_),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold479 (.A(\led_controller.rgbw.color[8] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold480 (.A(_1573_),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold481 (.A(\led_controller.effect_pulse_led_color[14] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold482 (.A(\led_controller.led_effect_pulse.calc_color_out[19] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold483 (.A(_3178_),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold484 (.A(\led_controller.rgbw.low_cycles[4] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold485 (.A(\led_controller.rgbw.color[17] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold486 (.A(_1618_),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold487 (.A(\led_controller.rgbw.color[1] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold488 (.A(_1538_),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold489 (.A(\led_controller.cpu.current_instruction_pc[1] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0368_),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold491 (.A(\led_controller.led_effect_chase.current_led[7] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0465_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold493 (.A(\led_controller.led_effect_pulse.calc_color_out[16] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold494 (.A(_3172_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold495 (.A(\led_controller.led_effect_pulse.calc_color_out[20] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold496 (.A(_3181_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold497 (.A(\led_controller.rgbw.color[7] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold498 (.A(_1568_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold499 (.A(\led_controller.rgbw.color[24] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold500 (.A(_1653_),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold501 (.A(\led_controller.rgbw.color[6] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold502 (.A(_1563_),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold503 (.A(\led_controller.spi_slave.data_bits[3] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0140_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold505 (.A(\led_controller.rgbw.color[18] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold506 (.A(_1623_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold507 (.A(\led_controller.rgbw.color[0] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold508 (.A(_1533_),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold509 (.A(\led_controller.rgbw.color[30] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold510 (.A(_1683_),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold511 (.A(\led_controller.rgbw.color[23] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold512 (.A(_1648_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold513 (.A(\led_controller.timer_2hz.counter[3] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold514 (.A(_1389_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold515 (.A(\led_controller.rgbw.color[20] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold516 (.A(_1633_),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold517 (.A(\led_controller.colors[46] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold518 (.A(_3501_),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold519 (.A(\led_controller.rgbw.color[21] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold520 (.A(_1638_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold521 (.A(\led_controller.flash.master.bit_counter[3] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold522 (.A(_2616_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0416_),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold524 (.A(\led_controller.rgbw.color[5] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold525 (.A(_1558_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold526 (.A(\led_controller.flash.master.tx_data[0] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold527 (.A(_2657_),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold528 (.A(\led_controller.led_effect_pulse.calc_color_out[23] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold529 (.A(_3190_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0556_),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold531 (.A(\led_controller.colors[66] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold532 (.A(_3524_),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold533 (.A(\led_controller.spi_data[5] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold534 (.A(_1354_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold535 (.A(\led_controller.timer_10hz.counter[0] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold536 (.A(_1396_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0170_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold538 (.A(\led_controller.rgbw.color[25] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold539 (.A(_1658_),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold540 (.A(\led_controller.rgbw.color[31] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold541 (.A(_1688_),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold542 (.A(\led_controller.rgbw.low_cycles[1] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold543 (.A(_1734_),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold544 (.A(\led_controller.cpu.i_bus_data[1] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold545 (.A(_0428_),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold546 (.A(\led_controller.led_effect_pulse.state[0] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0921_),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0011_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold549 (.A(\led_controller.rgbw.color[14] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold550 (.A(_1603_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold551 (.A(\led_controller.timer_2hz.counter[0] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold552 (.A(_1384_),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold553 (.A(_0164_),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold554 (.A(\led_controller.rgbw.color[10] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold555 (.A(_1583_),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold556 (.A(\led_controller.flash.cs_delay_counter[5] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold557 (.A(_2651_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0441_),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold559 (.A(\led_controller.rgbw.color[12] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold560 (.A(_1593_),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold561 (.A(\led_controller.rgbw.counter[3] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold562 (.A(_1321_),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold563 (.A(_0130_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold564 (.A(\led_controller.rgbw.color[29] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold565 (.A(_1678_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold566 (.A(\led_controller.cpu.o_bus_addr[2] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0328_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold568 (.A(\led_controller.rgbw.color[13] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold569 (.A(_1598_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold570 (.A(\led_controller.rgbw.pixel_counter[5] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0222_),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold572 (.A(\led_controller.cpu.i_bus_data[6] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0433_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold574 (.A(\led_controller.led_effect_pulse.color_index[0] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0524_),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold576 (.A(\led_controller.led_effect_pulse.current_led[7] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0523_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold578 (.A(\led_controller.rgbw.color[19] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold579 (.A(_1628_),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold580 (.A(\led_controller.cpu.fetch_instruction[7] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold581 (.A(_3212_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold582 (.A(\led_controller.spi_data_write[1] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold583 (.A(_3285_),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold584 (.A(\led_controller.colors[40] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold585 (.A(_3495_),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold586 (.A(\led_controller.spi_slave.mosi ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold587 (.A(_1349_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold588 (.A(\led_controller.colors[64] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold589 (.A(_3522_),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold590 (.A(\led_controller.colors[52] ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold591 (.A(_3508_),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold592 (.A(\led_controller.rgbw.color[28] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold593 (.A(_1673_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold594 (.A(\led_controller.cpu.fetch_instruction[1] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold595 (.A(_3206_),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold596 (.A(\led_controller.led_effect_pulse.calc_color_out[22] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold597 (.A(_3187_),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold598 (.A(\led_controller.rgbw.color[11] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold599 (.A(_1588_),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold600 (.A(\led_controller.colors[49] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold601 (.A(_3505_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold602 (.A(\led_controller.colors[44] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold603 (.A(_3499_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold604 (.A(\led_controller.cpu.i_bus_data[7] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold605 (.A(\led_controller.cpu.fetch_instruction[3] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold606 (.A(_3208_),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold607 (.A(\led_controller.cpu.i_bus_data[2] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold608 (.A(\led_controller.timer_100hz.counter[1] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold609 (.A(_1421_),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold610 (.A(_0176_),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold611 (.A(\led_controller.colors[70] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold612 (.A(_3528_),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold613 (.A(\led_controller.led_effect_pulse.current_led[1] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold614 (.A(_2825_),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold615 (.A(_0517_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold616 (.A(\led_controller.led_effect_pulse.calc_color_out[17] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold617 (.A(\led_controller.rgbw.color[15] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold618 (.A(_1608_),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold619 (.A(\led_controller.rgbw.color[22] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold620 (.A(_1643_),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold621 (.A(\led_controller.spi_slave.last_sck ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold622 (.A(_1334_),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold623 (.A(\led_controller.spi_data[2] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold624 (.A(_3384_),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold625 (.A(_0600_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold626 (.A(\led_controller.colors[92] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold627 (.A(_3555_),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold628 (.A(\led_controller.timer_2hz.counter[4] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold629 (.A(\led_controller.rgbw.color[4] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold630 (.A(_1553_),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold631 (.A(\led_controller.timer_100hz.div_counter[4] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold632 (.A(_1189_),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold633 (.A(_0068_),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold634 (.A(\led_controller.cpu.i_bus_data[4] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold635 (.A(\led_controller.spi_data[3] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold636 (.A(_3391_),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold637 (.A(_0601_),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold638 (.A(\led_controller.rgbw.counter[4] ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold639 (.A(_1323_),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold640 (.A(_0131_),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold641 (.A(\led_controller.flash.master.bit_counter[1] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold642 (.A(_2614_),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0414_),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold644 (.A(\led_controller.cpu.i_bus_data[5] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold645 (.A(\led_controller.cpu.current_instruction[12] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold646 (.A(\led_controller.led_effect_pulse.calc_color_out[9] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold647 (.A(_3160_),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold648 (.A(_0542_),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold649 (.A(\led_controller.timer_100hz.counter[28] ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold650 (.A(_1475_),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold651 (.A(_0203_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold652 (.A(\led_controller.colors[68] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold653 (.A(_3526_),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold654 (.A(\led_controller.cpu.o_bus_addr[5] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold655 (.A(_2475_),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0331_),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold657 (.A(\led_controller.colors[48] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold658 (.A(_3504_),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold659 (.A(\led_controller.spi_data_write[4] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold660 (.A(_3328_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold661 (.A(\led_controller.flash.master.sck_counter[3] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold662 (.A(_2624_),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold663 (.A(\led_controller.spi_slave.o_tx_start_strb ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold664 (.A(_0974_),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold665 (.A(_0016_),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold666 (.A(\led_controller.rgbw.counter[5] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0132_),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold668 (.A(\led_controller.colors[43] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold669 (.A(_3498_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold670 (.A(\led_controller.colors[65] ),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold671 (.A(_3523_),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold672 (.A(\led_controller.cpu.fetch_pc[7] ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold673 (.A(_0102_),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold674 (.A(\led_controller.cpu.fetch_pc_valid ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold675 (.A(_2572_),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold676 (.A(\led_controller.cpu.fetch_pc[11] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold677 (.A(_0106_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold678 (.A(\led_controller.cpu.current_instruction[10] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold679 (.A(\led_controller.colors[42] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold680 (.A(_3497_),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold681 (.A(\led_controller.timer_100hz.div_counter[3] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold682 (.A(_1187_),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold683 (.A(\led_controller.effect_pulse_led_strb ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0482_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold685 (.A(\led_controller.led_effect_pulse.calc_color_out[24] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold686 (.A(\led_controller.colors[95] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold687 (.A(_3558_),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold688 (.A(\led_controller.cpu.i_bus_data[0] ),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold689 (.A(\led_controller.cpu.fetch_instruction[4] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold690 (.A(_3209_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold691 (.A(\led_controller.led_effect_pulse.calc_color_out[31] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold692 (.A(\led_controller.colors[88] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold693 (.A(_3551_),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold694 (.A(\led_controller.cpu.o_bus_addr[4] ),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold695 (.A(_0330_),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold696 (.A(\led_controller.colors[41] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold697 (.A(_3496_),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold698 (.A(\led_controller.led_effect_pulse.current_led[2] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold699 (.A(_2828_),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold700 (.A(\led_controller.colors[47] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold701 (.A(_3502_),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold702 (.A(\led_controller.cpu.fetch_instruction[6] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold703 (.A(_3211_),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold704 (.A(\led_controller.colors[71] ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold705 (.A(_3529_),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold706 (.A(\led_controller.colors[94] ),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold707 (.A(_3557_),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold708 (.A(\led_controller.led_effect_pulse.calc_color_out[25] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold709 (.A(_0558_),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold710 (.A(\led_controller.rgbw.counter[1] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold711 (.A(_0128_),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold712 (.A(\led_controller.cpu.fetch_pc[9] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold713 (.A(_0104_),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold714 (.A(\led_controller.rgbw.state[0] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold715 (.A(_0013_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold716 (.A(\led_controller.timer_100hz.div_counter[5] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold717 (.A(\led_controller.led_effect_pulse.calc_color_out[2] ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold718 (.A(_3061_),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold719 (.A(_0535_),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold720 (.A(\led_controller.led_effect_pulse.current_led[6] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold721 (.A(_2835_),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold722 (.A(_0522_),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold723 (.A(\led_controller.colors[67] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold724 (.A(_3525_),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold725 (.A(\led_controller.spi_slave.data_bits[2] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold726 (.A(_1343_),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold727 (.A(_0139_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold728 (.A(\led_controller.rgbw.low_cycles[9] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold729 (.A(_0265_),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold730 (.A(\led_controller.flash.master.tx_data[4] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold731 (.A(_1797_),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold732 (.A(_0273_),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold733 (.A(\led_controller.timer_100hz.counter[13] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold734 (.A(_1444_),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold735 (.A(_0188_),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold736 (.A(\led_controller.led_effect_pulse.calc_color_out[0] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold737 (.A(\led_controller.flash.master.sck_counter[1] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold738 (.A(\led_controller.timer_100hz.counter[19] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold739 (.A(_1456_),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold740 (.A(_0194_),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold741 (.A(\led_controller.spi_slave.ss_n ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold742 (.A(\led_controller.cpu.fetch_pc[8] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold743 (.A(_0103_),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold744 (.A(\led_controller.spi_data[4] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold745 (.A(\led_controller.cpu.pc[8] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold746 (.A(\led_controller.cpu.fetch_instruction[5] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold747 (.A(_3210_),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold748 (.A(\led_controller.colors[24] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold749 (.A(_3460_),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold750 (.A(\led_controller.rgbw.color[2] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold751 (.A(_1543_),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold752 (.A(\led_controller.colors[69] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold753 (.A(_3527_),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold754 (.A(\led_controller.spi_data[7] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold755 (.A(\led_controller.cpu.fetch_pc[14] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold756 (.A(_0109_),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold757 (.A(\led_controller.colors[93] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold758 (.A(_3556_),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold759 (.A(\led_controller.led_effect_pulse.current_led[0] ),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold760 (.A(\led_controller.colors[76] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold761 (.A(_3537_),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold762 (.A(\led_controller.cpu.fetch_pc[6] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold763 (.A(_0101_),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold764 (.A(\led_controller.flash.master.sck_counter[6] ),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold765 (.A(_2630_),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold766 (.A(\led_controller.rgbw.counter[6] ),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold767 (.A(_0133_),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold768 (.A(\led_controller.timer_100hz.div_counter[1] ),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold769 (.A(\led_controller.led_effect_pulse.calc_color_out[28] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold770 (.A(_0561_),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold771 (.A(\led_controller.timer_100hz.counter[16] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold772 (.A(_1450_),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0191_),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold774 (.A(\led_controller.flash.state[1] ),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold775 (.A(_1002_),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold776 (.A(\led_controller.flash.master.tx_data[7] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold777 (.A(_1806_),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold778 (.A(_0276_),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold779 (.A(\led_controller.cpu.current_instruction[11] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold780 (.A(\led_controller.flash.o_cs_n ),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0388_),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold782 (.A(\led_controller.led_effect_pulse.calc_color_out[1] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold783 (.A(\led_controller.flash.master.tx_data[2] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold784 (.A(_1791_),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold785 (.A(_0271_),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold786 (.A(\led_controller.register_data[5] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold787 (.A(_0613_),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold788 (.A(\led_controller.led_effect_pulse.calc_color_out[21] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold789 (.A(_3184_),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold790 (.A(\led_controller.spi_data[1] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold791 (.A(_0599_),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold792 (.A(\led_controller.cpu.fetch_instruction[0] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold793 (.A(_3205_),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold794 (.A(\led_controller.flash.cs_delay_counter[4] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold795 (.A(_2650_),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold796 (.A(\led_controller.timer_100hz.counter[22] ),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold797 (.A(_1463_),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold798 (.A(_0197_),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold799 (.A(\led_controller.timer_10hz.counter[1] ),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold800 (.A(_1398_),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold801 (.A(_0171_),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold802 (.A(\led_controller.timer_100hz.counter[14] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold803 (.A(_1446_),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold804 (.A(\led_controller.spi_slave.data_bits[1] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold805 (.A(\led_controller.colors[16] ),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold806 (.A(_3442_),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold807 (.A(\led_controller.cpu.fetch_instruction[2] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold808 (.A(_3207_),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold809 (.A(\led_controller.cpu.fetch_pc[0] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold810 (.A(_2573_),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold811 (.A(_0386_),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold812 (.A(\led_controller.timer_100hz.div_counter[6] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold813 (.A(\led_controller.colors[89] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold814 (.A(_3552_),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold815 (.A(\led_controller.cpu.current_instruction_pc[7] ),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold816 (.A(\led_controller.rgbw.pixel_counter[3] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold817 (.A(_1513_),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold818 (.A(\led_controller.flash.master.tx_data[5] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold819 (.A(_1800_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold820 (.A(\led_controller.timer_10hz.counter[3] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold821 (.A(\led_controller.colors[54] ),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold822 (.A(_3510_),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold823 (.A(\led_controller.colors[34] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold824 (.A(_3482_),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold825 (.A(\led_controller.colors[72] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold826 (.A(_3533_),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold827 (.A(\led_controller.colors[36] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold828 (.A(_3486_),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold829 (.A(\led_controller.rgbw.color[3] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold830 (.A(_1548_),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold831 (.A(\led_controller.led_effect_pulse.calc_color_valid ),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold832 (.A(\led_controller.spi_data[0] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold833 (.A(\led_controller.clock_divider[5] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold834 (.A(\led_controller.colors[39] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold835 (.A(_3492_),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold836 (.A(\led_controller.colors[28] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold837 (.A(_3468_),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold838 (.A(\led_controller.register_data[3] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold839 (.A(_0611_),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold840 (.A(\led_controller.led_effect_pulse.color_index[1] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold841 (.A(_0525_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold842 (.A(\led_controller.rgbw.color[9] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold843 (.A(_1578_),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold844 (.A(\led_controller.colors[29] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold845 (.A(\led_controller.colors[78] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold846 (.A(_3539_),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold847 (.A(\led_controller.cpu.fetch_pc[3] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold848 (.A(_0098_),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold849 (.A(\led_controller.colors[91] ),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold850 (.A(\led_controller.spi_data_write[6] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold851 (.A(_3356_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold852 (.A(\led_controller.spi_state[1] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold853 (.A(\led_controller.led_effect_chase.i_reset_n ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold854 (.A(\led_controller.colors[17] ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold855 (.A(_3444_),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold856 (.A(\led_controller.colors[45] ),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold857 (.A(\led_controller.spi_data_write[2] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold858 (.A(_3300_),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold859 (.A(\led_controller.colors[20] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold860 (.A(_3450_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold861 (.A(\led_controller.timer_100hz.counter[8] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold862 (.A(_1436_),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold863 (.A(_0183_),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold864 (.A(\led_controller.rgbw.color[27] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold865 (.A(_1668_),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold866 (.A(\led_controller.rgbw.low_cycles[3] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold867 (.A(_0259_),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold868 (.A(\led_controller.colors[33] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold869 (.A(_3480_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold870 (.A(\led_controller.colors[80] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold871 (.A(_3542_),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold872 (.A(\led_controller.cpu.fetch_pc[15] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold873 (.A(_1295_),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold874 (.A(\led_controller.colors[38] ),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold875 (.A(_3490_),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold876 (.A(\led_controller.colors[90] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold877 (.A(_3553_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold878 (.A(\led_controller.spi_data_write[3] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold879 (.A(_3315_),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold880 (.A(\led_controller.register_data[7] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold881 (.A(_0711_),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold882 (.A(\led_controller.colors[74] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold883 (.A(_3535_),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold884 (.A(\led_controller.colors[53] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold885 (.A(\led_controller.register_data[4] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold886 (.A(\led_controller.colors[62] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold887 (.A(_3519_),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold888 (.A(\led_controller.led_effect_chase.current_led[3] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold889 (.A(_2735_),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold890 (.A(\led_controller.colors[55] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold891 (.A(\led_controller.colors[75] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold892 (.A(_3536_),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold893 (.A(\led_controller.cpu.current_instruction[9] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold894 (.A(\led_controller.cpu.pc[11] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold895 (.A(\led_controller.colors[26] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold896 (.A(_3464_),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold897 (.A(\led_controller.effect[3] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold898 (.A(\led_controller.cpu.pc[15] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold899 (.A(\led_controller.colors[35] ),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold900 (.A(\led_controller.colors[37] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold901 (.A(\led_controller.timer_100hz.counter[5] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold902 (.A(_1430_),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold903 (.A(_0180_),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold904 (.A(\led_controller.cpu.o_led_strb ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold905 (.A(_1807_),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold906 (.A(\led_controller.colors[32] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold907 (.A(_3478_),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold908 (.A(\led_controller.colors[56] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold909 (.A(_3513_),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold910 (.A(\led_controller.timer_100hz.counter[29] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold911 (.A(_1478_),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold912 (.A(_0204_),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold913 (.A(\led_controller.spi_data_write[5] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold914 (.A(_3342_),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold915 (.A(\led_controller.flash.state[4] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold916 (.A(_0010_),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold917 (.A(\led_controller.flash.master.bit_counter[2] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold918 (.A(_2615_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold919 (.A(\led_controller.rgbw.counter[7] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold920 (.A(\led_controller.register_address[5] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold921 (.A(_3399_),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold922 (.A(_3400_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold923 (.A(_3401_),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold924 (.A(\led_controller.cpu.i_num_leds[5] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold925 (.A(\led_controller.flash.state[6] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold926 (.A(\led_controller.colors[7] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold927 (.A(\led_controller.flash.master.i_tx_data[7] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold928 (.A(\led_controller.colors[4] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold929 (.A(\led_controller.register_data[2] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold930 (.A(\led_controller.rgbw.low_cycles[7] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold931 (.A(_1755_),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold932 (.A(\led_controller.timer_2hz.counter[5] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold933 (.A(\led_controller.timer_100hz.div_counter[7] ),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold934 (.A(\led_controller.rgbw.low_cycles[6] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold935 (.A(_1753_),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold936 (.A(\led_controller.colors[27] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold937 (.A(\led_controller.rgbw.low_cycles[8] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold938 (.A(\led_controller.flash.master.i_tx_data[3] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold939 (.A(\led_controller.cpu.o_bus_addr[3] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold940 (.A(_2466_),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold941 (.A(_0329_),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold942 (.A(\led_controller.timer_100hz.counter[6] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold943 (.A(_1432_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold944 (.A(_0181_),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold945 (.A(\led_controller.led_effect_chase.current_led[4] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold946 (.A(_2738_),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold947 (.A(\led_controller.rgbw.high_cycles[2] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold948 (.A(_0268_),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold949 (.A(\led_controller.clock_divider[7] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold950 (.A(\led_controller.rgbw.low_cycles[2] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold951 (.A(_0258_),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold952 (.A(\led_controller.led_effect_chase.current_led[5] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold953 (.A(_2741_),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold954 (.A(_0463_),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold955 (.A(\led_controller.flash.cs_delay_counter[3] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold956 (.A(\led_controller.effect[2] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold957 (.A(\led_controller.timer_100hz.counter[11] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold958 (.A(\led_controller.colors[22] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold959 (.A(_3454_),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold960 (.A(\led_controller.colors[2] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold961 (.A(_0610_),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold962 (.A(\led_controller.register_data[1] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold963 (.A(_0609_),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold964 (.A(\led_controller.colors[86] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold965 (.A(_3548_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold966 (.A(\led_controller.register_address[7] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold967 (.A(_0605_),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold968 (.A(\led_controller.led_effect_chase.current_led[2] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold969 (.A(_2731_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold970 (.A(\led_controller.clock_divider[4] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold971 (.A(\led_controller.colors[73] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold972 (.A(_3534_),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold973 (.A(\led_controller.colors[31] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold974 (.A(\led_controller.flash.master.i_tx_data[6] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold975 (.A(\led_controller.effect[1] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold976 (.A(\led_controller.cpu.led_write_pending ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold977 (.A(_1812_),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold978 (.A(\led_controller.register_data[6] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold979 (.A(_0614_),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold980 (.A(\led_controller.cpu.stall_counter[2] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold981 (.A(_0318_),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold982 (.A(\led_controller.clock_divider[3] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold983 (.A(\led_controller.colors[58] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold984 (.A(\led_controller.cpu.o_bus_addr[8] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold985 (.A(\led_controller.led_effect_pulse.current_led[5] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold986 (.A(_2833_),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold987 (.A(_0521_),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold988 (.A(\led_controller.colors[19] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold989 (.A(\led_controller.colors[87] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold990 (.A(\led_controller.cpu_reset_counter[2] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold991 (.A(_3230_),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold992 (.A(\led_controller.flash.master.i_tx_data[4] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold993 (.A(\led_controller.cpu.fetch_pc[4] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold994 (.A(_0099_),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold995 (.A(\led_controller.cpu.o_bus_addr[7] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold996 (.A(_2489_),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold997 (.A(\led_controller.timer_100hz.counter[0] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold998 (.A(_1420_),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold999 (.A(\led_controller.flash.master.sck_counter[7] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\led_controller.effect[0] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold1001 (.A(_0712_),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\led_controller.rgbw.low_cycles[5] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\led_controller.colors[84] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\led_controller.colors[85] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\led_controller.flash.master.sck_counter[4] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\led_controller.cpu.i_num_leds[6] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\led_controller.timer_100hz.counter[7] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold1008 (.A(_1434_),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_0182_),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\led_controller.rgbw.low_cycles[0] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\led_controller.colors[60] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\led_controller.timer_100hz.counter[26] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_1472_),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_0201_),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\led_controller.timer_100hz.counter[12] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\led_controller.colors[23] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\led_controller.colors[51] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\led_controller.colors[14] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold1019 (.A(_3437_),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\led_controller.timer_100hz.counter[18] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold1021 (.A(_1455_),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_0193_),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\led_controller.clock_divider[6] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\led_controller.cpu.status_zero ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\led_controller.clock_divider[2] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\led_controller.rgbw.high_cycles[1] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_0267_),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\led_controller.cpu.o_bus_addr[11] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_0337_),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\led_controller.cpu.current_instruction[8] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\led_controller.cpu.o_bus_addr[9] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_2499_),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\led_controller.clock_divider[1] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\led_controller.cpu.status_negative ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\led_controller.timer_100hz.counter[15] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold1036 (.A(_1449_),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\led_controller.colors[12] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\led_controller.timer_100hz.counter[2] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\led_controller.cpu.i_num_leds[4] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold1040 (.A(_0708_),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\led_controller.cpu.pc[10] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\led_controller.rgbw.pixel_counter[2] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold1043 (.A(_1510_),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\led_controller.colors[30] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\led_controller.colors[77] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\led_controller.cpu.i_num_leds[3] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold1047 (.A(_0707_),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\led_controller.cpu.register_y[2] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\led_controller.cpu.stall_counter[6] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold1050 (.A(_2439_),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\led_controller.rgbw.pixel_counter[4] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold1052 (.A(_1516_),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\led_controller.colors[83] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\led_controller.cpu.fetch_pc[2] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_0097_),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\led_controller.cpu.o_bus_addr[14] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_0340_),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\led_controller.cpu.o_bus_addr[6] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold1059 (.A(_2484_),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\led_controller.timer_100hz.counter[27] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold1061 (.A(_1474_),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\led_controller.cpu.fetch_pc[13] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_0108_),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\led_controller.cpu.fetch_pc[5] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold1065 (.A(_0100_),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\led_controller.led_effect_pulse.color_1.i_strb ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold1067 (.A(_2870_),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_0531_),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\led_controller.cpu.register_x[0] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\led_controller.cpu.stall_counter[0] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\led_controller.colors[50] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\led_controller.timer_100hz.counter[24] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold1073 (.A(_1468_),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\led_controller.cpu.o_bus_addr[12] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold1075 (.A(_2512_),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\led_controller.led_effect_pulse.finished ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold1077 (.A(_0515_),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\led_controller.led_effect_chase.current_led[0] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold1079 (.A(_2726_),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\led_controller.timer_100hz.counter[17] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\led_controller.flash.master.i_tx_data[1] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\led_controller.colors[63] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\led_controller.colors[59] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\led_controller.cpu.pc[13] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\led_controller.cpu.register_y[3] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\led_controller.cpu.pc[12] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\led_controller.colors[81] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\led_controller.colors[13] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\led_controller.colors[79] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\led_controller.cpu.i_num_leds[1] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_0705_),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\led_controller.colors[11] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold1093 (.A(_3431_),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\led_controller.cpu.register_x[6] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold1095 (.A(_0304_),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\led_controller.timer_100hz.counter[23] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_1466_),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold1098 (.A(_0198_),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\led_controller.colors[21] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\led_controller.colors[0] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_0608_),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\led_controller.cpu.i_num_colors[1] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\led_controller.colors[82] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\led_controller.cpu.current_instruction[1] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\led_controller.cpu.fetch_pc[10] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\led_controller.rgbw.high_cycles[0] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\led_controller.colors[18] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\led_controller.cpu.current_instruction[3] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\led_controller.colors[15] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\led_controller.cpu.fetch_pc[12] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold1111 (.A(_0107_),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\led_controller.colors[61] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\led_controller.timer_100hz.counter[21] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_1461_),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\led_controller.led_effect_pulse.brightness[4] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_0530_),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\led_controller.colors[10] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_3429_),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\led_controller.led_effect_pulse.brightness[2] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold1120 (.A(_0528_),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\led_controller.led_effect_pulse.fade_out ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\led_controller.led_effect_pulse.calc_color_out[29] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold1123 (.A(_3201_),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\led_controller.cpu.pc[9] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\led_controller.cpu.o_bus_addr[1] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\led_controller.cpu.stall_counter[1] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\led_controller.cpu.pc[14] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\led_controller.effect_chase_led_color[1] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_0456_),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\led_controller.cpu.current_instruction[2] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\led_controller.effect_chase_led_color[0] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold1132 (.A(_2685_),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\led_controller.cpu_reset_counter[0] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\led_controller.colors[57] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\led_controller.colors[9] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold1136 (.A(_3427_),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\led_controller.colors[25] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\led_controller.cpu.i_num_leds[2] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_0706_),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\led_controller.colors[8] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold1141 (.A(_3425_),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\led_controller.cpu.current_instruction[0] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\led_controller.register_address[4] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_3393_),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\led_controller.timer_100hz.counter[3] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\led_controller.flash.i_addr_width_24 ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_0581_),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\led_controller.flash.master.bit_counter[0] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\led_controller.led_effect_pulse.calc_color_out[30] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold1150 (.A(_3203_),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\led_controller.cpu.stall_counter[4] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\led_controller.register_data[0] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\led_controller.cpu.o_bus_addr_valid ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1154 (.A(_0342_),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\led_controller.spi_state[0] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\led_controller.cpu.register_y[7] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\led_controller.register_address[0] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_3381_),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\led_controller.cpu_reset_counter[1] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\led_controller.cpu.pc[4] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1161 (.A(_0286_),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\led_controller.timer_100hz.counter[25] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\led_controller.cpu.register_x[5] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\led_controller.cpu.i_num_leds[0] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\led_controller.led_effect_pulse.calc_color_out[27] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\led_controller.timer_100hz.counter[4] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1167 (.A(_1417_),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\led_controller.led_effect_chase.current_led[1] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_0459_),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\led_controller.cpu.register_x[3] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\led_controller.rgbw.pixel_counter[0] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_0217_),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\led_controller.cpu.register_y[6] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\led_controller.led_effect_pulse.brightness[3] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\led_controller.cpu.register_x[7] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_0305_),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\led_controller.cpu.fetch_pc[1] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1178 (.A(_0096_),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\led_controller.clock_divider[0] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\led_controller.cpu.stall_counter[5] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\led_controller.flash.cs_delay_counter[1] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1182 (.A(_0437_),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\led_controller.cpu.i_num_colors[0] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\led_controller.timer_100hz.counter[20] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\led_controller.timer_100hz.counter[20] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\led_controller.cpu.pc[6] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_2056_),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1188 (.A(_0288_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\led_controller.cpu.pc[2] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\led_controller.cpu.pc[3] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\led_controller.rgbw.state[2] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1192 (.A(_0015_),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\led_controller.flash.master.o_rx_data_valid ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\led_controller.cpu.register_y[1] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_2268_),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\led_controller.cpu.pc[5] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_2024_),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_0287_),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\led_controller.cpu.o_bus_addr_valid ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\led_controller.cpu.register_x[1] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\led_controller.cpu.pc[7] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\led_controller.cpu.led_write_strb ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\led_controller.led_effect_pulse.brightness[0] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\led_controller.led_effect_pulse.calc_color_out[3] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold1205 (.A(_3101_),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\led_controller.cpu.register_x[4] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\led_controller.cpu.pc[0] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\led_controller.flash.master.active ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\led_controller.cpu.register_y[4] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\led_controller.led_effect_pulse.brightness[1] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\led_controller.rgbw.state[1] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\led_controller.spi_state[2] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\led_controller.cpu.o_bus_addr[0] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\led_controller.rgbw.pixel_counter[1] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\led_controller.cpu.register_x[2] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\led_controller.cpu.register_y[0] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\led_controller.led_effect_chase.finished ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold1218 (.A(_2721_),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\led_controller.cpu.pc[1] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\led_controller.cpu.register_y[5] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\led_controller.led_effect_pulse.color_1.counter[0] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\led_controller.timer_100hz.counter[12] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_1445_),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\led_controller.timer_100hz.counter[7] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\led_controller.flash.master.sck_counter[4] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\led_controller.cpu.o_bus_addr[7] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\led_controller.cpu.current_instruction[2] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_1101_),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\led_controller.timer_100hz.div_counter[1] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\led_controller.cpu.register_x[6] ),
    .X(net2392));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_4 FILLER_0_77 ();
 sg13g2_fill_1 FILLER_0_81 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_4 FILLER_0_117 ();
 sg13g2_fill_2 FILLER_0_125 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_4 FILLER_0_175 ();
 sg13g2_fill_2 FILLER_0_179 ();
 sg13g2_fill_2 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_224 ();
 sg13g2_fill_1 FILLER_0_247 ();
 sg13g2_fill_2 FILLER_0_252 ();
 sg13g2_decap_4 FILLER_0_258 ();
 sg13g2_fill_1 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_267 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_fill_1 FILLER_0_288 ();
 sg13g2_fill_2 FILLER_0_293 ();
 sg13g2_decap_4 FILLER_0_317 ();
 sg13g2_fill_1 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_4 FILLER_0_333 ();
 sg13g2_fill_1 FILLER_0_337 ();
 sg13g2_fill_1 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_1 FILLER_0_407 ();
 sg13g2_decap_4 FILLER_0_412 ();
 sg13g2_fill_2 FILLER_0_416 ();
 sg13g2_fill_2 FILLER_0_445 ();
 sg13g2_decap_4 FILLER_0_452 ();
 sg13g2_fill_1 FILLER_0_456 ();
 sg13g2_decap_4 FILLER_0_465 ();
 sg13g2_fill_2 FILLER_0_469 ();
 sg13g2_fill_1 FILLER_0_480 ();
 sg13g2_decap_4 FILLER_0_485 ();
 sg13g2_fill_2 FILLER_0_489 ();
 sg13g2_fill_1 FILLER_0_535 ();
 sg13g2_decap_4 FILLER_0_544 ();
 sg13g2_fill_1 FILLER_0_548 ();
 sg13g2_decap_4 FILLER_0_558 ();
 sg13g2_decap_8 FILLER_0_571 ();
 sg13g2_decap_8 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_590 ();
 sg13g2_decap_4 FILLER_0_597 ();
 sg13g2_fill_1 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_646 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_754 ();
 sg13g2_fill_1 FILLER_0_795 ();
 sg13g2_fill_1 FILLER_0_810 ();
 sg13g2_fill_2 FILLER_0_826 ();
 sg13g2_fill_1 FILLER_0_828 ();
 sg13g2_fill_2 FILLER_0_860 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_51 ();
 sg13g2_fill_1 FILLER_1_68 ();
 sg13g2_fill_2 FILLER_1_85 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_fill_1 FILLER_1_115 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_228 ();
 sg13g2_fill_1 FILLER_1_238 ();
 sg13g2_fill_1 FILLER_1_254 ();
 sg13g2_decap_4 FILLER_1_311 ();
 sg13g2_fill_2 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_344 ();
 sg13g2_fill_2 FILLER_1_377 ();
 sg13g2_fill_1 FILLER_1_415 ();
 sg13g2_fill_2 FILLER_1_421 ();
 sg13g2_decap_4 FILLER_1_431 ();
 sg13g2_fill_1 FILLER_1_435 ();
 sg13g2_fill_2 FILLER_1_450 ();
 sg13g2_fill_2 FILLER_1_515 ();
 sg13g2_fill_2 FILLER_1_526 ();
 sg13g2_fill_1 FILLER_1_528 ();
 sg13g2_fill_2 FILLER_1_615 ();
 sg13g2_fill_1 FILLER_1_617 ();
 sg13g2_fill_2 FILLER_1_623 ();
 sg13g2_fill_1 FILLER_1_625 ();
 sg13g2_fill_2 FILLER_1_684 ();
 sg13g2_fill_1 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_696 ();
 sg13g2_decap_4 FILLER_1_703 ();
 sg13g2_fill_2 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_718 ();
 sg13g2_decap_8 FILLER_1_725 ();
 sg13g2_decap_8 FILLER_1_732 ();
 sg13g2_decap_8 FILLER_1_739 ();
 sg13g2_decap_8 FILLER_1_746 ();
 sg13g2_decap_8 FILLER_1_753 ();
 sg13g2_fill_2 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_25 ();
 sg13g2_decap_4 FILLER_2_92 ();
 sg13g2_fill_2 FILLER_2_96 ();
 sg13g2_fill_1 FILLER_2_119 ();
 sg13g2_decap_4 FILLER_2_138 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_fill_1 FILLER_2_147 ();
 sg13g2_decap_4 FILLER_2_169 ();
 sg13g2_fill_1 FILLER_2_173 ();
 sg13g2_fill_2 FILLER_2_183 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_fill_2 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_1 FILLER_2_242 ();
 sg13g2_fill_1 FILLER_2_249 ();
 sg13g2_fill_2 FILLER_2_258 ();
 sg13g2_fill_1 FILLER_2_260 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_fill_2 FILLER_2_305 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_fill_2 FILLER_2_340 ();
 sg13g2_fill_2 FILLER_2_364 ();
 sg13g2_fill_1 FILLER_2_366 ();
 sg13g2_fill_2 FILLER_2_394 ();
 sg13g2_fill_1 FILLER_2_406 ();
 sg13g2_fill_2 FILLER_2_437 ();
 sg13g2_decap_4 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_475 ();
 sg13g2_decap_8 FILLER_2_482 ();
 sg13g2_decap_4 FILLER_2_489 ();
 sg13g2_decap_4 FILLER_2_550 ();
 sg13g2_fill_1 FILLER_2_562 ();
 sg13g2_fill_2 FILLER_2_567 ();
 sg13g2_fill_1 FILLER_2_569 ();
 sg13g2_fill_2 FILLER_2_596 ();
 sg13g2_fill_1 FILLER_2_598 ();
 sg13g2_fill_1 FILLER_2_640 ();
 sg13g2_decap_4 FILLER_2_660 ();
 sg13g2_fill_2 FILLER_2_664 ();
 sg13g2_fill_1 FILLER_2_689 ();
 sg13g2_decap_8 FILLER_2_726 ();
 sg13g2_decap_8 FILLER_2_733 ();
 sg13g2_decap_8 FILLER_2_740 ();
 sg13g2_decap_4 FILLER_2_747 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_25 ();
 sg13g2_fill_2 FILLER_3_43 ();
 sg13g2_fill_1 FILLER_3_45 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_2 FILLER_3_73 ();
 sg13g2_fill_1 FILLER_3_75 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_decap_4 FILLER_3_87 ();
 sg13g2_decap_4 FILLER_3_99 ();
 sg13g2_fill_1 FILLER_3_103 ();
 sg13g2_decap_8 FILLER_3_124 ();
 sg13g2_decap_4 FILLER_3_131 ();
 sg13g2_fill_2 FILLER_3_135 ();
 sg13g2_fill_2 FILLER_3_142 ();
 sg13g2_decap_4 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_fill_2 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_fill_2 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_262 ();
 sg13g2_fill_2 FILLER_3_267 ();
 sg13g2_fill_1 FILLER_3_269 ();
 sg13g2_fill_1 FILLER_3_274 ();
 sg13g2_fill_2 FILLER_3_279 ();
 sg13g2_decap_4 FILLER_3_295 ();
 sg13g2_fill_2 FILLER_3_325 ();
 sg13g2_fill_2 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_418 ();
 sg13g2_decap_8 FILLER_3_425 ();
 sg13g2_decap_8 FILLER_3_432 ();
 sg13g2_fill_1 FILLER_3_439 ();
 sg13g2_fill_1 FILLER_3_452 ();
 sg13g2_fill_1 FILLER_3_475 ();
 sg13g2_decap_4 FILLER_3_489 ();
 sg13g2_fill_1 FILLER_3_503 ();
 sg13g2_fill_2 FILLER_3_509 ();
 sg13g2_fill_1 FILLER_3_511 ();
 sg13g2_fill_2 FILLER_3_581 ();
 sg13g2_decap_4 FILLER_3_596 ();
 sg13g2_fill_1 FILLER_3_630 ();
 sg13g2_fill_1 FILLER_3_635 ();
 sg13g2_fill_1 FILLER_3_650 ();
 sg13g2_fill_1 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_fill_1 FILLER_3_712 ();
 sg13g2_decap_8 FILLER_3_722 ();
 sg13g2_decap_8 FILLER_3_729 ();
 sg13g2_decap_4 FILLER_3_736 ();
 sg13g2_fill_2 FILLER_3_740 ();
 sg13g2_fill_2 FILLER_3_769 ();
 sg13g2_fill_2 FILLER_3_790 ();
 sg13g2_fill_1 FILLER_3_801 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_31 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_70 ();
 sg13g2_fill_2 FILLER_4_86 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_decap_8 FILLER_4_118 ();
 sg13g2_fill_1 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_166 ();
 sg13g2_decap_4 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_4 FILLER_4_189 ();
 sg13g2_fill_1 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_4 FILLER_4_205 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_2 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_decap_4 FILLER_4_243 ();
 sg13g2_fill_1 FILLER_4_247 ();
 sg13g2_decap_4 FILLER_4_265 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_fill_2 FILLER_4_326 ();
 sg13g2_fill_1 FILLER_4_328 ();
 sg13g2_decap_4 FILLER_4_337 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_decap_4 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_fill_2 FILLER_4_368 ();
 sg13g2_fill_1 FILLER_4_370 ();
 sg13g2_fill_1 FILLER_4_388 ();
 sg13g2_fill_1 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_4 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_481 ();
 sg13g2_fill_2 FILLER_4_540 ();
 sg13g2_fill_2 FILLER_4_564 ();
 sg13g2_decap_8 FILLER_4_570 ();
 sg13g2_decap_4 FILLER_4_577 ();
 sg13g2_fill_2 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_decap_8 FILLER_4_608 ();
 sg13g2_fill_2 FILLER_4_615 ();
 sg13g2_fill_1 FILLER_4_674 ();
 sg13g2_fill_2 FILLER_4_694 ();
 sg13g2_fill_1 FILLER_4_696 ();
 sg13g2_fill_1 FILLER_4_702 ();
 sg13g2_decap_8 FILLER_4_730 ();
 sg13g2_decap_8 FILLER_4_737 ();
 sg13g2_fill_2 FILLER_4_744 ();
 sg13g2_fill_1 FILLER_4_746 ();
 sg13g2_fill_2 FILLER_4_751 ();
 sg13g2_fill_1 FILLER_4_753 ();
 sg13g2_fill_2 FILLER_4_808 ();
 sg13g2_fill_1 FILLER_4_810 ();
 sg13g2_fill_2 FILLER_4_816 ();
 sg13g2_fill_2 FILLER_4_859 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_13 ();
 sg13g2_fill_2 FILLER_5_20 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_fill_2 FILLER_5_51 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_70 ();
 sg13g2_fill_2 FILLER_5_85 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_decap_8 FILLER_5_101 ();
 sg13g2_decap_4 FILLER_5_108 ();
 sg13g2_fill_1 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_fill_1 FILLER_5_161 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_fill_2 FILLER_5_307 ();
 sg13g2_decap_4 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_4 FILLER_5_365 ();
 sg13g2_fill_2 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_403 ();
 sg13g2_fill_1 FILLER_5_431 ();
 sg13g2_decap_4 FILLER_5_437 ();
 sg13g2_fill_1 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_446 ();
 sg13g2_decap_4 FILLER_5_453 ();
 sg13g2_fill_2 FILLER_5_457 ();
 sg13g2_decap_8 FILLER_5_463 ();
 sg13g2_decap_8 FILLER_5_484 ();
 sg13g2_decap_8 FILLER_5_491 ();
 sg13g2_decap_8 FILLER_5_498 ();
 sg13g2_decap_8 FILLER_5_505 ();
 sg13g2_decap_8 FILLER_5_534 ();
 sg13g2_fill_1 FILLER_5_541 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_fill_2 FILLER_5_584 ();
 sg13g2_fill_1 FILLER_5_586 ();
 sg13g2_decap_4 FILLER_5_623 ();
 sg13g2_fill_2 FILLER_5_627 ();
 sg13g2_fill_1 FILLER_5_639 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_4 FILLER_5_674 ();
 sg13g2_decap_4 FILLER_5_687 ();
 sg13g2_fill_2 FILLER_5_691 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_4 FILLER_5_704 ();
 sg13g2_fill_1 FILLER_5_712 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_fill_2 FILLER_5_729 ();
 sg13g2_decap_8 FILLER_5_748 ();
 sg13g2_fill_2 FILLER_5_755 ();
 sg13g2_fill_1 FILLER_5_757 ();
 sg13g2_fill_1 FILLER_5_804 ();
 sg13g2_fill_1 FILLER_5_818 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_9 ();
 sg13g2_fill_2 FILLER_6_38 ();
 sg13g2_fill_1 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_50 ();
 sg13g2_decap_8 FILLER_6_61 ();
 sg13g2_decap_8 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_75 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_162 ();
 sg13g2_decap_4 FILLER_6_169 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_179 ();
 sg13g2_decap_4 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_189 ();
 sg13g2_decap_4 FILLER_6_214 ();
 sg13g2_fill_1 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_decap_4 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_250 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_fill_1 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_4 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_4 FILLER_6_312 ();
 sg13g2_fill_1 FILLER_6_316 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_fill_1 FILLER_6_372 ();
 sg13g2_decap_4 FILLER_6_381 ();
 sg13g2_fill_2 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_fill_1 FILLER_6_416 ();
 sg13g2_decap_4 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_434 ();
 sg13g2_fill_1 FILLER_6_436 ();
 sg13g2_fill_1 FILLER_6_464 ();
 sg13g2_decap_8 FILLER_6_478 ();
 sg13g2_fill_2 FILLER_6_512 ();
 sg13g2_fill_1 FILLER_6_514 ();
 sg13g2_fill_1 FILLER_6_524 ();
 sg13g2_fill_2 FILLER_6_530 ();
 sg13g2_fill_1 FILLER_6_532 ();
 sg13g2_fill_2 FILLER_6_555 ();
 sg13g2_fill_2 FILLER_6_566 ();
 sg13g2_fill_1 FILLER_6_618 ();
 sg13g2_fill_2 FILLER_6_632 ();
 sg13g2_fill_1 FILLER_6_634 ();
 sg13g2_fill_2 FILLER_6_662 ();
 sg13g2_fill_2 FILLER_6_701 ();
 sg13g2_decap_4 FILLER_6_730 ();
 sg13g2_fill_2 FILLER_6_734 ();
 sg13g2_fill_1 FILLER_6_833 ();
 sg13g2_fill_1 FILLER_6_843 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_19 ();
 sg13g2_fill_2 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_28 ();
 sg13g2_fill_1 FILLER_7_33 ();
 sg13g2_decap_4 FILLER_7_38 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_48 ();
 sg13g2_fill_1 FILLER_7_65 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_fill_1 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_fill_2 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_decap_4 FILLER_7_160 ();
 sg13g2_fill_1 FILLER_7_164 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_1 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_258 ();
 sg13g2_decap_4 FILLER_7_333 ();
 sg13g2_fill_1 FILLER_7_337 ();
 sg13g2_fill_2 FILLER_7_360 ();
 sg13g2_fill_1 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_435 ();
 sg13g2_fill_1 FILLER_7_442 ();
 sg13g2_decap_4 FILLER_7_447 ();
 sg13g2_decap_4 FILLER_7_498 ();
 sg13g2_decap_4 FILLER_7_512 ();
 sg13g2_fill_2 FILLER_7_516 ();
 sg13g2_fill_1 FILLER_7_586 ();
 sg13g2_fill_1 FILLER_7_591 ();
 sg13g2_decap_8 FILLER_7_605 ();
 sg13g2_decap_8 FILLER_7_612 ();
 sg13g2_fill_2 FILLER_7_619 ();
 sg13g2_fill_1 FILLER_7_629 ();
 sg13g2_fill_1 FILLER_7_634 ();
 sg13g2_fill_2 FILLER_7_644 ();
 sg13g2_fill_1 FILLER_7_646 ();
 sg13g2_fill_2 FILLER_7_673 ();
 sg13g2_fill_2 FILLER_7_697 ();
 sg13g2_decap_8 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_737 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_751 ();
 sg13g2_fill_1 FILLER_7_787 ();
 sg13g2_fill_2 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_51 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_decap_4 FILLER_8_75 ();
 sg13g2_fill_1 FILLER_8_79 ();
 sg13g2_fill_2 FILLER_8_84 ();
 sg13g2_fill_1 FILLER_8_86 ();
 sg13g2_fill_2 FILLER_8_100 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_107 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_decap_8 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_143 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_fill_2 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_242 ();
 sg13g2_fill_2 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_276 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_decap_4 FILLER_8_302 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_311 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_fill_1 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_408 ();
 sg13g2_decap_4 FILLER_8_415 ();
 sg13g2_fill_1 FILLER_8_419 ();
 sg13g2_fill_1 FILLER_8_441 ();
 sg13g2_fill_1 FILLER_8_488 ();
 sg13g2_decap_8 FILLER_8_516 ();
 sg13g2_fill_1 FILLER_8_523 ();
 sg13g2_fill_2 FILLER_8_537 ();
 sg13g2_fill_1 FILLER_8_539 ();
 sg13g2_decap_4 FILLER_8_545 ();
 sg13g2_fill_1 FILLER_8_549 ();
 sg13g2_fill_2 FILLER_8_555 ();
 sg13g2_decap_4 FILLER_8_584 ();
 sg13g2_fill_2 FILLER_8_588 ();
 sg13g2_fill_2 FILLER_8_608 ();
 sg13g2_fill_1 FILLER_8_610 ();
 sg13g2_fill_2 FILLER_8_643 ();
 sg13g2_fill_1 FILLER_8_645 ();
 sg13g2_fill_2 FILLER_8_711 ();
 sg13g2_fill_1 FILLER_8_713 ();
 sg13g2_fill_1 FILLER_8_727 ();
 sg13g2_fill_2 FILLER_8_859 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_15 ();
 sg13g2_decap_4 FILLER_9_22 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_2 FILLER_9_45 ();
 sg13g2_fill_1 FILLER_9_47 ();
 sg13g2_fill_1 FILLER_9_76 ();
 sg13g2_decap_4 FILLER_9_96 ();
 sg13g2_fill_1 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_121 ();
 sg13g2_fill_2 FILLER_9_128 ();
 sg13g2_decap_4 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_decap_4 FILLER_9_215 ();
 sg13g2_fill_2 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_decap_4 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_4 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_1 FILLER_9_299 ();
 sg13g2_decap_4 FILLER_9_313 ();
 sg13g2_decap_4 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_decap_4 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_335 ();
 sg13g2_fill_2 FILLER_9_354 ();
 sg13g2_decap_4 FILLER_9_396 ();
 sg13g2_fill_1 FILLER_9_400 ();
 sg13g2_fill_1 FILLER_9_432 ();
 sg13g2_decap_4 FILLER_9_438 ();
 sg13g2_fill_1 FILLER_9_442 ();
 sg13g2_decap_8 FILLER_9_447 ();
 sg13g2_decap_8 FILLER_9_454 ();
 sg13g2_fill_1 FILLER_9_461 ();
 sg13g2_fill_2 FILLER_9_480 ();
 sg13g2_fill_2 FILLER_9_491 ();
 sg13g2_fill_1 FILLER_9_493 ();
 sg13g2_fill_2 FILLER_9_498 ();
 sg13g2_fill_2 FILLER_9_507 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_fill_1 FILLER_9_529 ();
 sg13g2_fill_1 FILLER_9_543 ();
 sg13g2_fill_1 FILLER_9_574 ();
 sg13g2_decap_4 FILLER_9_632 ();
 sg13g2_decap_4 FILLER_9_649 ();
 sg13g2_fill_1 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_663 ();
 sg13g2_fill_1 FILLER_9_670 ();
 sg13g2_fill_2 FILLER_9_675 ();
 sg13g2_fill_1 FILLER_9_690 ();
 sg13g2_fill_2 FILLER_9_718 ();
 sg13g2_fill_1 FILLER_9_720 ();
 sg13g2_fill_1 FILLER_9_734 ();
 sg13g2_decap_4 FILLER_9_757 ();
 sg13g2_fill_2 FILLER_9_761 ();
 sg13g2_fill_1 FILLER_9_785 ();
 sg13g2_fill_1 FILLER_9_810 ();
 sg13g2_fill_1 FILLER_9_825 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_34 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_4 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_decap_4 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_decap_4 FILLER_10_246 ();
 sg13g2_fill_2 FILLER_10_292 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_355 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_decap_4 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_409 ();
 sg13g2_fill_1 FILLER_10_411 ();
 sg13g2_fill_1 FILLER_10_465 ();
 sg13g2_fill_2 FILLER_10_479 ();
 sg13g2_fill_2 FILLER_10_486 ();
 sg13g2_fill_1 FILLER_10_493 ();
 sg13g2_fill_2 FILLER_10_500 ();
 sg13g2_fill_2 FILLER_10_521 ();
 sg13g2_fill_2 FILLER_10_559 ();
 sg13g2_fill_1 FILLER_10_561 ();
 sg13g2_fill_2 FILLER_10_619 ();
 sg13g2_fill_1 FILLER_10_621 ();
 sg13g2_fill_2 FILLER_10_676 ();
 sg13g2_fill_1 FILLER_10_678 ();
 sg13g2_fill_2 FILLER_10_701 ();
 sg13g2_fill_2 FILLER_10_716 ();
 sg13g2_fill_1 FILLER_10_718 ();
 sg13g2_fill_2 FILLER_10_761 ();
 sg13g2_fill_2 FILLER_10_815 ();
 sg13g2_fill_1 FILLER_10_817 ();
 sg13g2_fill_1 FILLER_10_836 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_2 FILLER_11_31 ();
 sg13g2_fill_1 FILLER_11_33 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_87 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_decap_4 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_fill_2 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_fill_2 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_263 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_decap_4 FILLER_11_367 ();
 sg13g2_fill_2 FILLER_11_450 ();
 sg13g2_fill_2 FILLER_11_474 ();
 sg13g2_fill_1 FILLER_11_485 ();
 sg13g2_decap_4 FILLER_11_493 ();
 sg13g2_decap_4 FILLER_11_505 ();
 sg13g2_fill_1 FILLER_11_509 ();
 sg13g2_decap_8 FILLER_11_545 ();
 sg13g2_decap_4 FILLER_11_584 ();
 sg13g2_fill_1 FILLER_11_588 ();
 sg13g2_fill_1 FILLER_11_625 ();
 sg13g2_fill_1 FILLER_11_630 ();
 sg13g2_decap_4 FILLER_11_636 ();
 sg13g2_fill_1 FILLER_11_640 ();
 sg13g2_fill_2 FILLER_11_645 ();
 sg13g2_fill_1 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_656 ();
 sg13g2_fill_1 FILLER_11_663 ();
 sg13g2_fill_2 FILLER_11_762 ();
 sg13g2_fill_2 FILLER_11_772 ();
 sg13g2_fill_2 FILLER_11_823 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_12 ();
 sg13g2_fill_1 FILLER_12_43 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_decap_8 FILLER_12_66 ();
 sg13g2_decap_4 FILLER_12_73 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_decap_4 FILLER_12_186 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_fill_2 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_287 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_339 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_fill_2 FILLER_12_356 ();
 sg13g2_fill_1 FILLER_12_358 ();
 sg13g2_fill_2 FILLER_12_380 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_fill_2 FILLER_12_392 ();
 sg13g2_fill_1 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_4 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_428 ();
 sg13g2_fill_2 FILLER_12_435 ();
 sg13g2_fill_1 FILLER_12_437 ();
 sg13g2_fill_2 FILLER_12_455 ();
 sg13g2_fill_1 FILLER_12_484 ();
 sg13g2_decap_8 FILLER_12_489 ();
 sg13g2_decap_8 FILLER_12_496 ();
 sg13g2_decap_4 FILLER_12_503 ();
 sg13g2_fill_1 FILLER_12_507 ();
 sg13g2_decap_4 FILLER_12_521 ();
 sg13g2_fill_1 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_4 FILLER_12_550 ();
 sg13g2_fill_1 FILLER_12_554 ();
 sg13g2_decap_8 FILLER_12_559 ();
 sg13g2_fill_1 FILLER_12_566 ();
 sg13g2_fill_2 FILLER_12_580 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_fill_2 FILLER_12_597 ();
 sg13g2_fill_1 FILLER_12_635 ();
 sg13g2_fill_2 FILLER_12_676 ();
 sg13g2_fill_1 FILLER_12_697 ();
 sg13g2_fill_2 FILLER_12_734 ();
 sg13g2_fill_1 FILLER_12_736 ();
 sg13g2_fill_2 FILLER_12_804 ();
 sg13g2_fill_1 FILLER_12_806 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_23 ();
 sg13g2_fill_2 FILLER_13_32 ();
 sg13g2_decap_4 FILLER_13_46 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_4 FILLER_13_172 ();
 sg13g2_fill_2 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_fill_2 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_228 ();
 sg13g2_fill_2 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_decap_4 FILLER_13_279 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_365 ();
 sg13g2_fill_2 FILLER_13_415 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_decap_4 FILLER_13_472 ();
 sg13g2_fill_1 FILLER_13_476 ();
 sg13g2_fill_2 FILLER_13_481 ();
 sg13g2_fill_1 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_516 ();
 sg13g2_decap_4 FILLER_13_523 ();
 sg13g2_fill_2 FILLER_13_570 ();
 sg13g2_fill_1 FILLER_13_572 ();
 sg13g2_fill_2 FILLER_13_595 ();
 sg13g2_fill_1 FILLER_13_597 ();
 sg13g2_fill_2 FILLER_13_615 ();
 sg13g2_decap_4 FILLER_13_632 ();
 sg13g2_fill_2 FILLER_13_645 ();
 sg13g2_decap_8 FILLER_13_709 ();
 sg13g2_fill_2 FILLER_13_716 ();
 sg13g2_fill_1 FILLER_13_726 ();
 sg13g2_fill_1 FILLER_13_772 ();
 sg13g2_fill_2 FILLER_13_812 ();
 sg13g2_fill_1 FILLER_13_814 ();
 sg13g2_fill_2 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_29 ();
 sg13g2_decap_8 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_54 ();
 sg13g2_decap_8 FILLER_14_65 ();
 sg13g2_decap_8 FILLER_14_72 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_fill_1 FILLER_14_94 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_4 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_2 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_327 ();
 sg13g2_fill_2 FILLER_14_337 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_4 FILLER_14_419 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_fill_2 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_454 ();
 sg13g2_fill_2 FILLER_14_461 ();
 sg13g2_fill_2 FILLER_14_472 ();
 sg13g2_fill_1 FILLER_14_474 ();
 sg13g2_fill_2 FILLER_14_489 ();
 sg13g2_fill_1 FILLER_14_491 ();
 sg13g2_fill_1 FILLER_14_505 ();
 sg13g2_fill_2 FILLER_14_535 ();
 sg13g2_fill_1 FILLER_14_537 ();
 sg13g2_fill_2 FILLER_14_556 ();
 sg13g2_decap_4 FILLER_14_607 ();
 sg13g2_fill_2 FILLER_14_611 ();
 sg13g2_fill_2 FILLER_14_640 ();
 sg13g2_fill_2 FILLER_14_647 ();
 sg13g2_fill_1 FILLER_14_649 ();
 sg13g2_decap_8 FILLER_14_667 ();
 sg13g2_decap_4 FILLER_14_678 ();
 sg13g2_fill_2 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_4 FILLER_14_705 ();
 sg13g2_fill_1 FILLER_14_709 ();
 sg13g2_fill_1 FILLER_14_715 ();
 sg13g2_fill_2 FILLER_14_726 ();
 sg13g2_fill_1 FILLER_14_737 ();
 sg13g2_fill_1 FILLER_14_777 ();
 sg13g2_fill_2 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_59 ();
 sg13g2_fill_2 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_75 ();
 sg13g2_fill_2 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_122 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_decap_4 FILLER_15_214 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_234 ();
 sg13g2_decap_4 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_253 ();
 sg13g2_fill_2 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_fill_1 FILLER_15_283 ();
 sg13g2_decap_4 FILLER_15_302 ();
 sg13g2_decap_4 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_437 ();
 sg13g2_decap_4 FILLER_15_444 ();
 sg13g2_fill_1 FILLER_15_475 ();
 sg13g2_fill_2 FILLER_15_507 ();
 sg13g2_fill_1 FILLER_15_545 ();
 sg13g2_fill_2 FILLER_15_555 ();
 sg13g2_fill_1 FILLER_15_557 ();
 sg13g2_fill_1 FILLER_15_566 ();
 sg13g2_fill_2 FILLER_15_576 ();
 sg13g2_fill_2 FILLER_15_615 ();
 sg13g2_fill_1 FILLER_15_617 ();
 sg13g2_fill_2 FILLER_15_622 ();
 sg13g2_fill_1 FILLER_15_624 ();
 sg13g2_fill_1 FILLER_15_684 ();
 sg13g2_fill_2 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_4 FILLER_15_707 ();
 sg13g2_fill_1 FILLER_15_721 ();
 sg13g2_fill_1 FILLER_15_730 ();
 sg13g2_fill_2 FILLER_15_749 ();
 sg13g2_fill_1 FILLER_15_751 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_fill_1 FILLER_16_18 ();
 sg13g2_decap_4 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_61 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_decap_4 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_decap_4 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_159 ();
 sg13g2_decap_4 FILLER_16_166 ();
 sg13g2_decap_4 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_fill_1 FILLER_16_313 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_fill_1 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_394 ();
 sg13g2_fill_1 FILLER_16_402 ();
 sg13g2_fill_1 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_fill_1 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_434 ();
 sg13g2_fill_2 FILLER_16_447 ();
 sg13g2_fill_1 FILLER_16_449 ();
 sg13g2_fill_1 FILLER_16_471 ();
 sg13g2_fill_2 FILLER_16_488 ();
 sg13g2_fill_1 FILLER_16_512 ();
 sg13g2_fill_1 FILLER_16_607 ();
 sg13g2_decap_8 FILLER_16_621 ();
 sg13g2_fill_2 FILLER_16_628 ();
 sg13g2_decap_8 FILLER_16_643 ();
 sg13g2_fill_2 FILLER_16_650 ();
 sg13g2_decap_4 FILLER_16_656 ();
 sg13g2_fill_2 FILLER_16_660 ();
 sg13g2_fill_2 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_768 ();
 sg13g2_decap_4 FILLER_16_775 ();
 sg13g2_fill_2 FILLER_16_832 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_44 ();
 sg13g2_decap_4 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_58 ();
 sg13g2_decap_4 FILLER_17_65 ();
 sg13g2_decap_4 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_94 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_135 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_decap_4 FILLER_17_232 ();
 sg13g2_decap_4 FILLER_17_241 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_decap_4 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_4 FILLER_17_296 ();
 sg13g2_decap_4 FILLER_17_314 ();
 sg13g2_fill_2 FILLER_17_318 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_4 FILLER_17_414 ();
 sg13g2_fill_1 FILLER_17_418 ();
 sg13g2_fill_2 FILLER_17_429 ();
 sg13g2_decap_4 FILLER_17_436 ();
 sg13g2_fill_2 FILLER_17_440 ();
 sg13g2_fill_1 FILLER_17_448 ();
 sg13g2_fill_2 FILLER_17_475 ();
 sg13g2_fill_1 FILLER_17_477 ();
 sg13g2_fill_2 FILLER_17_495 ();
 sg13g2_decap_4 FILLER_17_505 ();
 sg13g2_fill_1 FILLER_17_557 ();
 sg13g2_fill_1 FILLER_17_572 ();
 sg13g2_fill_2 FILLER_17_587 ();
 sg13g2_fill_2 FILLER_17_602 ();
 sg13g2_fill_1 FILLER_17_604 ();
 sg13g2_decap_8 FILLER_17_660 ();
 sg13g2_fill_2 FILLER_17_685 ();
 sg13g2_decap_8 FILLER_17_692 ();
 sg13g2_decap_4 FILLER_17_699 ();
 sg13g2_fill_1 FILLER_17_703 ();
 sg13g2_decap_8 FILLER_17_717 ();
 sg13g2_decap_4 FILLER_17_724 ();
 sg13g2_fill_2 FILLER_17_741 ();
 sg13g2_fill_1 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_fill_1 FILLER_17_777 ();
 sg13g2_fill_2 FILLER_17_806 ();
 sg13g2_fill_2 FILLER_17_821 ();
 sg13g2_fill_1 FILLER_17_843 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_17 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_51 ();
 sg13g2_decap_4 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_decap_4 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_278 ();
 sg13g2_fill_2 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_fill_2 FILLER_18_416 ();
 sg13g2_fill_2 FILLER_18_431 ();
 sg13g2_fill_1 FILLER_18_433 ();
 sg13g2_decap_8 FILLER_18_443 ();
 sg13g2_fill_1 FILLER_18_450 ();
 sg13g2_fill_1 FILLER_18_466 ();
 sg13g2_decap_4 FILLER_18_472 ();
 sg13g2_fill_1 FILLER_18_476 ();
 sg13g2_fill_2 FILLER_18_498 ();
 sg13g2_fill_2 FILLER_18_531 ();
 sg13g2_fill_2 FILLER_18_552 ();
 sg13g2_fill_2 FILLER_18_558 ();
 sg13g2_fill_2 FILLER_18_570 ();
 sg13g2_fill_1 FILLER_18_572 ();
 sg13g2_fill_1 FILLER_18_619 ();
 sg13g2_decap_4 FILLER_18_628 ();
 sg13g2_fill_1 FILLER_18_632 ();
 sg13g2_fill_1 FILLER_18_647 ();
 sg13g2_fill_2 FILLER_18_661 ();
 sg13g2_fill_1 FILLER_18_663 ();
 sg13g2_decap_4 FILLER_18_672 ();
 sg13g2_fill_2 FILLER_18_676 ();
 sg13g2_fill_2 FILLER_18_688 ();
 sg13g2_fill_1 FILLER_18_690 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_fill_1 FILLER_18_730 ();
 sg13g2_fill_2 FILLER_18_736 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_4 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_fill_2 FILLER_18_823 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_decap_8 FILLER_19_40 ();
 sg13g2_decap_8 FILLER_19_47 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_decap_8 FILLER_19_83 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_fill_2 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_176 ();
 sg13g2_decap_4 FILLER_19_183 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_309 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_decap_4 FILLER_19_385 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_fill_2 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_442 ();
 sg13g2_decap_4 FILLER_19_449 ();
 sg13g2_fill_1 FILLER_19_453 ();
 sg13g2_fill_2 FILLER_19_460 ();
 sg13g2_fill_1 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_fill_1 FILLER_19_492 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_fill_1 FILLER_19_522 ();
 sg13g2_fill_1 FILLER_19_574 ();
 sg13g2_fill_1 FILLER_19_593 ();
 sg13g2_fill_2 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_615 ();
 sg13g2_fill_1 FILLER_19_622 ();
 sg13g2_fill_1 FILLER_19_639 ();
 sg13g2_fill_2 FILLER_19_684 ();
 sg13g2_fill_2 FILLER_19_702 ();
 sg13g2_decap_8 FILLER_19_717 ();
 sg13g2_decap_8 FILLER_19_724 ();
 sg13g2_fill_2 FILLER_19_740 ();
 sg13g2_fill_1 FILLER_19_742 ();
 sg13g2_fill_1 FILLER_19_747 ();
 sg13g2_fill_2 FILLER_19_788 ();
 sg13g2_fill_2 FILLER_19_832 ();
 sg13g2_fill_1 FILLER_19_834 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_10 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_319 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_453 ();
 sg13g2_decap_4 FILLER_20_460 ();
 sg13g2_fill_1 FILLER_20_495 ();
 sg13g2_fill_1 FILLER_20_532 ();
 sg13g2_fill_2 FILLER_20_537 ();
 sg13g2_fill_2 FILLER_20_580 ();
 sg13g2_fill_2 FILLER_20_645 ();
 sg13g2_fill_2 FILLER_20_656 ();
 sg13g2_fill_1 FILLER_20_671 ();
 sg13g2_fill_2 FILLER_20_686 ();
 sg13g2_fill_2 FILLER_20_697 ();
 sg13g2_decap_4 FILLER_20_704 ();
 sg13g2_fill_2 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_fill_2 FILLER_20_745 ();
 sg13g2_fill_1 FILLER_20_778 ();
 sg13g2_fill_2 FILLER_20_815 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_65 ();
 sg13g2_fill_2 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_decap_4 FILLER_21_333 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_fill_1 FILLER_21_384 ();
 sg13g2_fill_1 FILLER_21_394 ();
 sg13g2_fill_1 FILLER_21_470 ();
 sg13g2_decap_4 FILLER_21_498 ();
 sg13g2_fill_1 FILLER_21_502 ();
 sg13g2_fill_2 FILLER_21_508 ();
 sg13g2_fill_1 FILLER_21_510 ();
 sg13g2_fill_2 FILLER_21_546 ();
 sg13g2_fill_2 FILLER_21_561 ();
 sg13g2_fill_1 FILLER_21_563 ();
 sg13g2_fill_2 FILLER_21_581 ();
 sg13g2_fill_2 FILLER_21_596 ();
 sg13g2_fill_2 FILLER_21_611 ();
 sg13g2_decap_8 FILLER_21_617 ();
 sg13g2_decap_4 FILLER_21_624 ();
 sg13g2_fill_1 FILLER_21_669 ();
 sg13g2_decap_8 FILLER_21_774 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_decap_4 FILLER_22_94 ();
 sg13g2_decap_4 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_decap_4 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_425 ();
 sg13g2_decap_8 FILLER_22_432 ();
 sg13g2_fill_2 FILLER_22_439 ();
 sg13g2_fill_1 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_446 ();
 sg13g2_decap_4 FILLER_22_453 ();
 sg13g2_fill_1 FILLER_22_457 ();
 sg13g2_fill_1 FILLER_22_494 ();
 sg13g2_fill_1 FILLER_22_535 ();
 sg13g2_fill_2 FILLER_22_563 ();
 sg13g2_fill_2 FILLER_22_597 ();
 sg13g2_fill_2 FILLER_22_639 ();
 sg13g2_fill_2 FILLER_22_646 ();
 sg13g2_fill_1 FILLER_22_648 ();
 sg13g2_fill_2 FILLER_22_653 ();
 sg13g2_fill_1 FILLER_22_655 ();
 sg13g2_fill_2 FILLER_22_673 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_fill_1 FILLER_22_700 ();
 sg13g2_fill_2 FILLER_22_732 ();
 sg13g2_fill_1 FILLER_22_734 ();
 sg13g2_fill_1 FILLER_22_748 ();
 sg13g2_decap_8 FILLER_22_762 ();
 sg13g2_decap_8 FILLER_22_769 ();
 sg13g2_decap_4 FILLER_22_776 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_1 FILLER_23_31 ();
 sg13g2_fill_1 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_64 ();
 sg13g2_decap_4 FILLER_23_87 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_106 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_4 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_decap_4 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_318 ();
 sg13g2_fill_2 FILLER_23_351 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_fill_2 FILLER_23_464 ();
 sg13g2_fill_1 FILLER_23_466 ();
 sg13g2_fill_2 FILLER_23_476 ();
 sg13g2_fill_1 FILLER_23_478 ();
 sg13g2_fill_1 FILLER_23_493 ();
 sg13g2_fill_2 FILLER_23_522 ();
 sg13g2_fill_1 FILLER_23_524 ();
 sg13g2_fill_1 FILLER_23_543 ();
 sg13g2_fill_2 FILLER_23_610 ();
 sg13g2_fill_1 FILLER_23_612 ();
 sg13g2_fill_1 FILLER_23_639 ();
 sg13g2_decap_4 FILLER_23_689 ();
 sg13g2_fill_1 FILLER_23_693 ();
 sg13g2_fill_1 FILLER_23_753 ();
 sg13g2_fill_1 FILLER_23_785 ();
 sg13g2_fill_2 FILLER_23_808 ();
 sg13g2_fill_1 FILLER_23_810 ();
 sg13g2_fill_1 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_10 ();
 sg13g2_fill_1 FILLER_24_12 ();
 sg13g2_decap_8 FILLER_24_17 ();
 sg13g2_fill_2 FILLER_24_24 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_decap_4 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_fill_2 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_4 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_24_421 ();
 sg13g2_decap_8 FILLER_24_436 ();
 sg13g2_fill_2 FILLER_24_443 ();
 sg13g2_fill_1 FILLER_24_445 ();
 sg13g2_decap_4 FILLER_24_450 ();
 sg13g2_fill_2 FILLER_24_454 ();
 sg13g2_fill_2 FILLER_24_474 ();
 sg13g2_fill_1 FILLER_24_476 ();
 sg13g2_decap_4 FILLER_24_517 ();
 sg13g2_fill_1 FILLER_24_521 ();
 sg13g2_fill_2 FILLER_24_562 ();
 sg13g2_fill_1 FILLER_24_564 ();
 sg13g2_fill_1 FILLER_24_578 ();
 sg13g2_fill_2 FILLER_24_588 ();
 sg13g2_fill_2 FILLER_24_629 ();
 sg13g2_fill_1 FILLER_24_631 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_4 FILLER_24_665 ();
 sg13g2_fill_1 FILLER_24_669 ();
 sg13g2_fill_2 FILLER_24_714 ();
 sg13g2_fill_1 FILLER_24_716 ();
 sg13g2_fill_1 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_855 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_decap_4 FILLER_25_103 ();
 sg13g2_fill_2 FILLER_25_111 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_fill_2 FILLER_25_490 ();
 sg13g2_fill_1 FILLER_25_492 ();
 sg13g2_fill_2 FILLER_25_549 ();
 sg13g2_fill_1 FILLER_25_551 ();
 sg13g2_fill_2 FILLER_25_592 ();
 sg13g2_fill_1 FILLER_25_594 ();
 sg13g2_fill_2 FILLER_25_631 ();
 sg13g2_decap_4 FILLER_25_674 ();
 sg13g2_fill_1 FILLER_25_678 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_4 FILLER_25_690 ();
 sg13g2_fill_1 FILLER_25_694 ();
 sg13g2_fill_2 FILLER_25_722 ();
 sg13g2_fill_2 FILLER_25_733 ();
 sg13g2_fill_1 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_767 ();
 sg13g2_fill_2 FILLER_25_778 ();
 sg13g2_fill_1 FILLER_25_780 ();
 sg13g2_decap_8 FILLER_25_836 ();
 sg13g2_decap_8 FILLER_25_843 ();
 sg13g2_decap_8 FILLER_25_850 ();
 sg13g2_decap_4 FILLER_25_857 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_11 ();
 sg13g2_fill_1 FILLER_26_24 ();
 sg13g2_fill_2 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_decap_4 FILLER_26_145 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_404 ();
 sg13g2_decap_4 FILLER_26_414 ();
 sg13g2_fill_1 FILLER_26_440 ();
 sg13g2_decap_4 FILLER_26_446 ();
 sg13g2_fill_2 FILLER_26_450 ();
 sg13g2_fill_2 FILLER_26_465 ();
 sg13g2_fill_1 FILLER_26_467 ();
 sg13g2_decap_4 FILLER_26_473 ();
 sg13g2_fill_2 FILLER_26_504 ();
 sg13g2_fill_1 FILLER_26_551 ();
 sg13g2_fill_1 FILLER_26_598 ();
 sg13g2_fill_1 FILLER_26_621 ();
 sg13g2_fill_1 FILLER_26_673 ();
 sg13g2_fill_2 FILLER_26_777 ();
 sg13g2_fill_2 FILLER_26_787 ();
 sg13g2_decap_8 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_855 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_59 ();
 sg13g2_decap_4 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_decap_4 FILLER_27_349 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_432 ();
 sg13g2_fill_1 FILLER_27_434 ();
 sg13g2_fill_2 FILLER_27_467 ();
 sg13g2_fill_1 FILLER_27_469 ();
 sg13g2_fill_2 FILLER_27_500 ();
 sg13g2_fill_1 FILLER_27_502 ();
 sg13g2_fill_2 FILLER_27_556 ();
 sg13g2_fill_1 FILLER_27_558 ();
 sg13g2_fill_2 FILLER_27_604 ();
 sg13g2_fill_1 FILLER_27_606 ();
 sg13g2_fill_2 FILLER_27_634 ();
 sg13g2_fill_1 FILLER_27_636 ();
 sg13g2_decap_8 FILLER_27_668 ();
 sg13g2_fill_2 FILLER_27_675 ();
 sg13g2_fill_1 FILLER_27_677 ();
 sg13g2_decap_8 FILLER_27_682 ();
 sg13g2_decap_8 FILLER_27_689 ();
 sg13g2_fill_1 FILLER_27_700 ();
 sg13g2_fill_2 FILLER_27_709 ();
 sg13g2_fill_1 FILLER_27_729 ();
 sg13g2_fill_2 FILLER_27_753 ();
 sg13g2_fill_2 FILLER_27_763 ();
 sg13g2_fill_1 FILLER_27_793 ();
 sg13g2_fill_2 FILLER_27_798 ();
 sg13g2_fill_1 FILLER_27_800 ();
 sg13g2_fill_2 FILLER_27_808 ();
 sg13g2_fill_1 FILLER_27_827 ();
 sg13g2_decap_8 FILLER_27_841 ();
 sg13g2_decap_8 FILLER_27_848 ();
 sg13g2_decap_8 FILLER_27_855 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_411 ();
 sg13g2_fill_1 FILLER_28_413 ();
 sg13g2_fill_1 FILLER_28_417 ();
 sg13g2_fill_2 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_435 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_fill_2 FILLER_28_519 ();
 sg13g2_fill_1 FILLER_28_521 ();
 sg13g2_decap_4 FILLER_28_531 ();
 sg13g2_fill_2 FILLER_28_567 ();
 sg13g2_fill_2 FILLER_28_577 ();
 sg13g2_fill_1 FILLER_28_632 ();
 sg13g2_decap_4 FILLER_28_668 ();
 sg13g2_fill_1 FILLER_28_672 ();
 sg13g2_fill_1 FILLER_28_701 ();
 sg13g2_fill_1 FILLER_28_751 ();
 sg13g2_fill_2 FILLER_28_803 ();
 sg13g2_fill_2 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_decap_4 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_424 ();
 sg13g2_decap_8 FILLER_29_461 ();
 sg13g2_fill_2 FILLER_29_468 ();
 sg13g2_decap_4 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_550 ();
 sg13g2_fill_2 FILLER_29_557 ();
 sg13g2_fill_1 FILLER_29_559 ();
 sg13g2_fill_2 FILLER_29_564 ();
 sg13g2_fill_1 FILLER_29_566 ();
 sg13g2_decap_4 FILLER_29_572 ();
 sg13g2_fill_2 FILLER_29_576 ();
 sg13g2_fill_2 FILLER_29_602 ();
 sg13g2_fill_1 FILLER_29_604 ();
 sg13g2_decap_4 FILLER_29_673 ();
 sg13g2_fill_2 FILLER_29_677 ();
 sg13g2_fill_2 FILLER_29_702 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_decap_4 FILLER_29_740 ();
 sg13g2_fill_1 FILLER_29_764 ();
 sg13g2_fill_2 FILLER_29_787 ();
 sg13g2_fill_1 FILLER_29_789 ();
 sg13g2_fill_2 FILLER_29_799 ();
 sg13g2_fill_1 FILLER_29_801 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_decap_8 FILLER_30_407 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_4 FILLER_30_434 ();
 sg13g2_fill_1 FILLER_30_438 ();
 sg13g2_decap_8 FILLER_30_443 ();
 sg13g2_decap_8 FILLER_30_450 ();
 sg13g2_fill_1 FILLER_30_485 ();
 sg13g2_decap_4 FILLER_30_503 ();
 sg13g2_fill_1 FILLER_30_507 ();
 sg13g2_decap_8 FILLER_30_536 ();
 sg13g2_decap_4 FILLER_30_543 ();
 sg13g2_fill_2 FILLER_30_630 ();
 sg13g2_fill_2 FILLER_30_643 ();
 sg13g2_fill_2 FILLER_30_744 ();
 sg13g2_fill_2 FILLER_30_758 ();
 sg13g2_fill_1 FILLER_30_760 ();
 sg13g2_fill_2 FILLER_30_833 ();
 sg13g2_fill_1 FILLER_30_835 ();
 sg13g2_fill_2 FILLER_30_845 ();
 sg13g2_fill_1 FILLER_30_847 ();
 sg13g2_decap_4 FILLER_31_116 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_4 FILLER_31_371 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_decap_8 FILLER_31_438 ();
 sg13g2_fill_2 FILLER_31_445 ();
 sg13g2_decap_8 FILLER_31_451 ();
 sg13g2_decap_4 FILLER_31_458 ();
 sg13g2_fill_1 FILLER_31_466 ();
 sg13g2_decap_4 FILLER_31_485 ();
 sg13g2_fill_2 FILLER_31_522 ();
 sg13g2_fill_1 FILLER_31_524 ();
 sg13g2_fill_2 FILLER_31_585 ();
 sg13g2_fill_1 FILLER_31_587 ();
 sg13g2_fill_2 FILLER_31_647 ();
 sg13g2_fill_1 FILLER_31_658 ();
 sg13g2_fill_1 FILLER_31_668 ();
 sg13g2_fill_2 FILLER_31_678 ();
 sg13g2_fill_1 FILLER_31_680 ();
 sg13g2_decap_4 FILLER_31_694 ();
 sg13g2_fill_1 FILLER_31_698 ();
 sg13g2_fill_2 FILLER_31_708 ();
 sg13g2_fill_1 FILLER_31_710 ();
 sg13g2_fill_1 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_734 ();
 sg13g2_fill_1 FILLER_31_741 ();
 sg13g2_fill_1 FILLER_31_784 ();
 sg13g2_decap_4 FILLER_31_794 ();
 sg13g2_fill_2 FILLER_31_798 ();
 sg13g2_fill_2 FILLER_31_826 ();
 sg13g2_fill_1 FILLER_31_828 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_9 ();
 sg13g2_fill_2 FILLER_32_16 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_45 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_decap_4 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_decap_4 FILLER_32_400 ();
 sg13g2_fill_1 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_499 ();
 sg13g2_decap_4 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_513 ();
 sg13g2_fill_2 FILLER_32_519 ();
 sg13g2_fill_1 FILLER_32_521 ();
 sg13g2_fill_1 FILLER_32_531 ();
 sg13g2_decap_4 FILLER_32_545 ();
 sg13g2_fill_2 FILLER_32_549 ();
 sg13g2_fill_1 FILLER_32_556 ();
 sg13g2_fill_1 FILLER_32_576 ();
 sg13g2_fill_2 FILLER_32_628 ();
 sg13g2_fill_2 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_717 ();
 sg13g2_fill_1 FILLER_32_724 ();
 sg13g2_fill_1 FILLER_32_741 ();
 sg13g2_fill_2 FILLER_32_755 ();
 sg13g2_fill_1 FILLER_32_757 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_10 ();
 sg13g2_decap_8 FILLER_33_17 ();
 sg13g2_decap_8 FILLER_33_44 ();
 sg13g2_decap_4 FILLER_33_51 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_83 ();
 sg13g2_decap_8 FILLER_33_90 ();
 sg13g2_decap_4 FILLER_33_97 ();
 sg13g2_decap_8 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_113 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_4 FILLER_33_142 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_245 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_271 ();
 sg13g2_decap_8 FILLER_33_278 ();
 sg13g2_decap_4 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_324 ();
 sg13g2_decap_4 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_450 ();
 sg13g2_fill_2 FILLER_33_454 ();
 sg13g2_fill_2 FILLER_33_475 ();
 sg13g2_fill_1 FILLER_33_477 ();
 sg13g2_fill_1 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_538 ();
 sg13g2_decap_4 FILLER_33_545 ();
 sg13g2_fill_1 FILLER_33_566 ();
 sg13g2_fill_1 FILLER_33_579 ();
 sg13g2_fill_2 FILLER_33_584 ();
 sg13g2_fill_1 FILLER_33_586 ();
 sg13g2_decap_4 FILLER_33_614 ();
 sg13g2_fill_2 FILLER_33_629 ();
 sg13g2_fill_1 FILLER_33_640 ();
 sg13g2_fill_2 FILLER_33_687 ();
 sg13g2_fill_1 FILLER_33_689 ();
 sg13g2_fill_1 FILLER_33_708 ();
 sg13g2_fill_2 FILLER_33_722 ();
 sg13g2_fill_1 FILLER_33_724 ();
 sg13g2_decap_8 FILLER_33_739 ();
 sg13g2_decap_4 FILLER_33_746 ();
 sg13g2_fill_1 FILLER_33_750 ();
 sg13g2_fill_1 FILLER_33_756 ();
 sg13g2_fill_2 FILLER_33_794 ();
 sg13g2_fill_1 FILLER_33_796 ();
 sg13g2_fill_2 FILLER_33_849 ();
 sg13g2_fill_1 FILLER_33_851 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_43 ();
 sg13g2_fill_1 FILLER_34_47 ();
 sg13g2_fill_2 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_116 ();
 sg13g2_decap_4 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_139 ();
 sg13g2_decap_4 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_decap_4 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_446 ();
 sg13g2_decap_8 FILLER_34_451 ();
 sg13g2_fill_2 FILLER_34_458 ();
 sg13g2_fill_2 FILLER_34_466 ();
 sg13g2_fill_2 FILLER_34_474 ();
 sg13g2_fill_1 FILLER_34_495 ();
 sg13g2_fill_1 FILLER_34_510 ();
 sg13g2_fill_1 FILLER_34_548 ();
 sg13g2_fill_2 FILLER_34_563 ();
 sg13g2_fill_1 FILLER_34_565 ();
 sg13g2_fill_2 FILLER_34_632 ();
 sg13g2_fill_1 FILLER_34_644 ();
 sg13g2_decap_4 FILLER_34_697 ();
 sg13g2_fill_2 FILLER_34_708 ();
 sg13g2_fill_2 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_725 ();
 sg13g2_fill_1 FILLER_34_732 ();
 sg13g2_decap_4 FILLER_34_741 ();
 sg13g2_fill_1 FILLER_34_745 ();
 sg13g2_fill_1 FILLER_34_762 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_decap_4 FILLER_35_90 ();
 sg13g2_decap_4 FILLER_35_106 ();
 sg13g2_decap_8 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_125 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_1 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_decap_8 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_decap_4 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_398 ();
 sg13g2_fill_1 FILLER_35_400 ();
 sg13g2_fill_1 FILLER_35_412 ();
 sg13g2_fill_2 FILLER_35_423 ();
 sg13g2_fill_1 FILLER_35_425 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_fill_2 FILLER_35_476 ();
 sg13g2_fill_2 FILLER_35_497 ();
 sg13g2_fill_1 FILLER_35_499 ();
 sg13g2_fill_2 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_fill_2 FILLER_35_546 ();
 sg13g2_fill_2 FILLER_35_572 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_fill_2 FILLER_35_595 ();
 sg13g2_decap_4 FILLER_35_612 ();
 sg13g2_fill_1 FILLER_35_616 ();
 sg13g2_fill_2 FILLER_35_622 ();
 sg13g2_fill_1 FILLER_35_624 ();
 sg13g2_fill_2 FILLER_35_636 ();
 sg13g2_fill_1 FILLER_35_638 ();
 sg13g2_fill_1 FILLER_35_655 ();
 sg13g2_decap_8 FILLER_35_701 ();
 sg13g2_fill_2 FILLER_35_708 ();
 sg13g2_fill_1 FILLER_35_710 ();
 sg13g2_fill_2 FILLER_35_732 ();
 sg13g2_fill_2 FILLER_35_762 ();
 sg13g2_fill_2 FILLER_35_777 ();
 sg13g2_fill_1 FILLER_35_779 ();
 sg13g2_fill_1 FILLER_35_793 ();
 sg13g2_fill_1 FILLER_35_831 ();
 sg13g2_fill_2 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_decap_4 FILLER_36_23 ();
 sg13g2_decap_4 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_decap_8 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_fill_2 FILLER_36_430 ();
 sg13g2_fill_1 FILLER_36_432 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_fill_1 FILLER_36_462 ();
 sg13g2_fill_1 FILLER_36_475 ();
 sg13g2_fill_1 FILLER_36_481 ();
 sg13g2_fill_1 FILLER_36_505 ();
 sg13g2_fill_1 FILLER_36_510 ();
 sg13g2_fill_1 FILLER_36_553 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_fill_1 FILLER_36_614 ();
 sg13g2_fill_2 FILLER_36_623 ();
 sg13g2_fill_1 FILLER_36_625 ();
 sg13g2_decap_4 FILLER_36_658 ();
 sg13g2_fill_2 FILLER_36_674 ();
 sg13g2_fill_1 FILLER_36_695 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_fill_2 FILLER_36_707 ();
 sg13g2_fill_1 FILLER_36_709 ();
 sg13g2_fill_2 FILLER_36_737 ();
 sg13g2_fill_1 FILLER_36_739 ();
 sg13g2_decap_4 FILLER_36_748 ();
 sg13g2_fill_1 FILLER_36_768 ();
 sg13g2_fill_1 FILLER_36_815 ();
 sg13g2_fill_2 FILLER_36_820 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_146 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_4 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_decap_4 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_394 ();
 sg13g2_fill_2 FILLER_37_399 ();
 sg13g2_fill_1 FILLER_37_401 ();
 sg13g2_fill_2 FILLER_37_411 ();
 sg13g2_fill_1 FILLER_37_413 ();
 sg13g2_fill_1 FILLER_37_455 ();
 sg13g2_fill_1 FILLER_37_482 ();
 sg13g2_fill_2 FILLER_37_487 ();
 sg13g2_fill_1 FILLER_37_489 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_fill_1 FILLER_37_539 ();
 sg13g2_fill_1 FILLER_37_558 ();
 sg13g2_decap_8 FILLER_37_572 ();
 sg13g2_decap_8 FILLER_37_579 ();
 sg13g2_decap_8 FILLER_37_586 ();
 sg13g2_fill_1 FILLER_37_593 ();
 sg13g2_fill_2 FILLER_37_606 ();
 sg13g2_fill_1 FILLER_37_608 ();
 sg13g2_decap_8 FILLER_37_620 ();
 sg13g2_decap_8 FILLER_37_627 ();
 sg13g2_decap_8 FILLER_37_634 ();
 sg13g2_fill_1 FILLER_37_641 ();
 sg13g2_fill_2 FILLER_37_647 ();
 sg13g2_fill_1 FILLER_37_654 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_fill_1 FILLER_37_772 ();
 sg13g2_fill_2 FILLER_37_785 ();
 sg13g2_decap_4 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_decap_4 FILLER_38_53 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_171 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_4 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_decap_8 FILLER_38_443 ();
 sg13g2_decap_8 FILLER_38_450 ();
 sg13g2_fill_2 FILLER_38_463 ();
 sg13g2_fill_1 FILLER_38_465 ();
 sg13g2_decap_4 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_484 ();
 sg13g2_fill_1 FILLER_38_491 ();
 sg13g2_decap_4 FILLER_38_497 ();
 sg13g2_fill_1 FILLER_38_538 ();
 sg13g2_decap_4 FILLER_38_586 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_fill_2 FILLER_38_617 ();
 sg13g2_fill_1 FILLER_38_619 ();
 sg13g2_fill_2 FILLER_38_629 ();
 sg13g2_fill_1 FILLER_38_631 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_fill_2 FILLER_38_658 ();
 sg13g2_fill_1 FILLER_38_664 ();
 sg13g2_fill_1 FILLER_38_675 ();
 sg13g2_fill_2 FILLER_38_681 ();
 sg13g2_fill_1 FILLER_38_683 ();
 sg13g2_fill_1 FILLER_38_709 ();
 sg13g2_fill_2 FILLER_38_734 ();
 sg13g2_fill_2 FILLER_38_764 ();
 sg13g2_fill_1 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_45 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_56 ();
 sg13g2_fill_2 FILLER_39_129 ();
 sg13g2_decap_4 FILLER_39_207 ();
 sg13g2_fill_2 FILLER_39_248 ();
 sg13g2_decap_4 FILLER_39_260 ();
 sg13g2_fill_2 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_283 ();
 sg13g2_fill_2 FILLER_39_314 ();
 sg13g2_fill_1 FILLER_39_316 ();
 sg13g2_decap_4 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_326 ();
 sg13g2_decap_4 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_decap_4 FILLER_39_402 ();
 sg13g2_fill_1 FILLER_39_411 ();
 sg13g2_decap_8 FILLER_39_418 ();
 sg13g2_decap_8 FILLER_39_425 ();
 sg13g2_decap_4 FILLER_39_445 ();
 sg13g2_fill_1 FILLER_39_457 ();
 sg13g2_fill_2 FILLER_39_477 ();
 sg13g2_fill_1 FILLER_39_479 ();
 sg13g2_decap_4 FILLER_39_512 ();
 sg13g2_fill_1 FILLER_39_544 ();
 sg13g2_decap_8 FILLER_39_573 ();
 sg13g2_decap_8 FILLER_39_580 ();
 sg13g2_fill_1 FILLER_39_587 ();
 sg13g2_decap_8 FILLER_39_592 ();
 sg13g2_decap_8 FILLER_39_599 ();
 sg13g2_decap_4 FILLER_39_606 ();
 sg13g2_fill_2 FILLER_39_610 ();
 sg13g2_decap_4 FILLER_39_640 ();
 sg13g2_fill_1 FILLER_39_676 ();
 sg13g2_fill_2 FILLER_39_691 ();
 sg13g2_fill_1 FILLER_39_693 ();
 sg13g2_fill_2 FILLER_39_708 ();
 sg13g2_fill_1 FILLER_39_817 ();
 sg13g2_fill_2 FILLER_39_827 ();
 sg13g2_fill_1 FILLER_39_838 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_13 ();
 sg13g2_fill_2 FILLER_40_20 ();
 sg13g2_fill_1 FILLER_40_22 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_49 ();
 sg13g2_fill_1 FILLER_40_111 ();
 sg13g2_decap_4 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_194 ();
 sg13g2_fill_2 FILLER_40_235 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_249 ();
 sg13g2_decap_4 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_259 ();
 sg13g2_fill_1 FILLER_40_288 ();
 sg13g2_fill_1 FILLER_40_327 ();
 sg13g2_decap_4 FILLER_40_334 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_fill_1 FILLER_40_379 ();
 sg13g2_fill_2 FILLER_40_390 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_decap_4 FILLER_40_426 ();
 sg13g2_fill_1 FILLER_40_430 ();
 sg13g2_fill_1 FILLER_40_444 ();
 sg13g2_decap_8 FILLER_40_450 ();
 sg13g2_fill_2 FILLER_40_461 ();
 sg13g2_fill_1 FILLER_40_479 ();
 sg13g2_fill_1 FILLER_40_520 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_decap_8 FILLER_40_571 ();
 sg13g2_fill_1 FILLER_40_578 ();
 sg13g2_decap_4 FILLER_40_611 ();
 sg13g2_fill_2 FILLER_40_615 ();
 sg13g2_decap_8 FILLER_40_621 ();
 sg13g2_fill_2 FILLER_40_628 ();
 sg13g2_fill_1 FILLER_40_630 ();
 sg13g2_decap_4 FILLER_40_671 ();
 sg13g2_fill_2 FILLER_40_703 ();
 sg13g2_fill_1 FILLER_40_705 ();
 sg13g2_fill_2 FILLER_40_710 ();
 sg13g2_fill_2 FILLER_40_767 ();
 sg13g2_fill_1 FILLER_40_769 ();
 sg13g2_decap_8 FILLER_40_778 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_fill_2 FILLER_40_792 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_fill_1 FILLER_40_846 ();
 sg13g2_decap_4 FILLER_40_856 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_43 ();
 sg13g2_fill_2 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_73 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_fill_2 FILLER_41_114 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_decap_4 FILLER_41_199 ();
 sg13g2_fill_1 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_263 ();
 sg13g2_decap_4 FILLER_41_270 ();
 sg13g2_fill_2 FILLER_41_291 ();
 sg13g2_fill_2 FILLER_41_322 ();
 sg13g2_decap_4 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_354 ();
 sg13g2_decap_4 FILLER_41_377 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_decap_4 FILLER_41_407 ();
 sg13g2_decap_4 FILLER_41_417 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_fill_1 FILLER_41_452 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_494 ();
 sg13g2_fill_2 FILLER_41_501 ();
 sg13g2_fill_1 FILLER_41_503 ();
 sg13g2_decap_4 FILLER_41_530 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_fill_1 FILLER_41_592 ();
 sg13g2_decap_4 FILLER_41_621 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_decap_4 FILLER_41_640 ();
 sg13g2_fill_2 FILLER_41_644 ();
 sg13g2_fill_1 FILLER_41_681 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_fill_2 FILLER_41_742 ();
 sg13g2_fill_2 FILLER_41_757 ();
 sg13g2_fill_1 FILLER_41_759 ();
 sg13g2_fill_1 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_fill_1 FILLER_41_810 ();
 sg13g2_fill_2 FILLER_41_823 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_4 ();
 sg13g2_decap_4 FILLER_42_10 ();
 sg13g2_fill_2 FILLER_42_118 ();
 sg13g2_fill_1 FILLER_42_120 ();
 sg13g2_decap_8 FILLER_42_125 ();
 sg13g2_decap_8 FILLER_42_132 ();
 sg13g2_decap_8 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_213 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_fill_1 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_fill_1 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_433 ();
 sg13g2_fill_1 FILLER_42_440 ();
 sg13g2_decap_8 FILLER_42_446 ();
 sg13g2_fill_1 FILLER_42_453 ();
 sg13g2_fill_1 FILLER_42_472 ();
 sg13g2_decap_8 FILLER_42_499 ();
 sg13g2_fill_2 FILLER_42_506 ();
 sg13g2_fill_1 FILLER_42_508 ();
 sg13g2_decap_8 FILLER_42_522 ();
 sg13g2_fill_1 FILLER_42_529 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_4 FILLER_42_560 ();
 sg13g2_fill_1 FILLER_42_568 ();
 sg13g2_fill_2 FILLER_42_590 ();
 sg13g2_fill_1 FILLER_42_592 ();
 sg13g2_fill_2 FILLER_42_610 ();
 sg13g2_fill_1 FILLER_42_612 ();
 sg13g2_fill_2 FILLER_42_617 ();
 sg13g2_fill_1 FILLER_42_619 ();
 sg13g2_fill_1 FILLER_42_648 ();
 sg13g2_fill_1 FILLER_42_677 ();
 sg13g2_fill_2 FILLER_42_703 ();
 sg13g2_fill_2 FILLER_42_708 ();
 sg13g2_fill_2 FILLER_42_734 ();
 sg13g2_fill_2 FILLER_42_763 ();
 sg13g2_fill_2 FILLER_42_774 ();
 sg13g2_fill_1 FILLER_42_776 ();
 sg13g2_fill_2 FILLER_42_782 ();
 sg13g2_fill_1 FILLER_42_784 ();
 sg13g2_fill_1 FILLER_42_821 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_4 ();
 sg13g2_fill_2 FILLER_43_10 ();
 sg13g2_fill_1 FILLER_43_12 ();
 sg13g2_decap_8 FILLER_43_80 ();
 sg13g2_fill_1 FILLER_43_87 ();
 sg13g2_decap_4 FILLER_43_96 ();
 sg13g2_decap_8 FILLER_43_109 ();
 sg13g2_decap_4 FILLER_43_116 ();
 sg13g2_fill_1 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_188 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_decap_4 FILLER_43_195 ();
 sg13g2_decap_4 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_decap_8 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_240 ();
 sg13g2_decap_8 FILLER_43_260 ();
 sg13g2_fill_2 FILLER_43_313 ();
 sg13g2_fill_2 FILLER_43_381 ();
 sg13g2_fill_1 FILLER_43_383 ();
 sg13g2_fill_1 FILLER_43_412 ();
 sg13g2_fill_2 FILLER_43_441 ();
 sg13g2_fill_1 FILLER_43_443 ();
 sg13g2_fill_1 FILLER_43_453 ();
 sg13g2_decap_4 FILLER_43_458 ();
 sg13g2_fill_2 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_471 ();
 sg13g2_fill_1 FILLER_43_478 ();
 sg13g2_fill_1 FILLER_43_485 ();
 sg13g2_decap_8 FILLER_43_519 ();
 sg13g2_fill_2 FILLER_43_554 ();
 sg13g2_fill_1 FILLER_43_556 ();
 sg13g2_fill_1 FILLER_43_561 ();
 sg13g2_fill_1 FILLER_43_583 ();
 sg13g2_fill_2 FILLER_43_629 ();
 sg13g2_fill_1 FILLER_43_631 ();
 sg13g2_decap_8 FILLER_43_645 ();
 sg13g2_decap_8 FILLER_43_652 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_fill_1 FILLER_43_666 ();
 sg13g2_fill_2 FILLER_43_675 ();
 sg13g2_fill_1 FILLER_43_705 ();
 sg13g2_fill_2 FILLER_43_776 ();
 sg13g2_decap_8 FILLER_43_797 ();
 sg13g2_decap_8 FILLER_43_804 ();
 sg13g2_fill_2 FILLER_43_811 ();
 sg13g2_fill_1 FILLER_43_813 ();
 sg13g2_decap_8 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_841 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_48 ();
 sg13g2_decap_4 FILLER_44_138 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_149 ();
 sg13g2_fill_2 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_156 ();
 sg13g2_decap_4 FILLER_44_213 ();
 sg13g2_fill_1 FILLER_44_217 ();
 sg13g2_decap_4 FILLER_44_278 ();
 sg13g2_fill_2 FILLER_44_282 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_fill_1 FILLER_44_331 ();
 sg13g2_fill_2 FILLER_44_361 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_fill_2 FILLER_44_415 ();
 sg13g2_fill_1 FILLER_44_417 ();
 sg13g2_decap_4 FILLER_44_422 ();
 sg13g2_fill_2 FILLER_44_477 ();
 sg13g2_fill_2 FILLER_44_488 ();
 sg13g2_fill_1 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_509 ();
 sg13g2_fill_2 FILLER_44_570 ();
 sg13g2_fill_2 FILLER_44_590 ();
 sg13g2_fill_1 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_653 ();
 sg13g2_fill_2 FILLER_44_660 ();
 sg13g2_decap_4 FILLER_44_675 ();
 sg13g2_fill_1 FILLER_44_715 ();
 sg13g2_fill_2 FILLER_44_726 ();
 sg13g2_decap_4 FILLER_44_758 ();
 sg13g2_fill_2 FILLER_44_779 ();
 sg13g2_fill_1 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_787 ();
 sg13g2_decap_4 FILLER_44_794 ();
 sg13g2_fill_2 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_827 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_855 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_20 ();
 sg13g2_fill_1 FILLER_45_22 ();
 sg13g2_fill_1 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_55 ();
 sg13g2_fill_2 FILLER_45_90 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_decap_4 FILLER_45_121 ();
 sg13g2_fill_2 FILLER_45_125 ();
 sg13g2_fill_2 FILLER_45_132 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_fill_2 FILLER_45_158 ();
 sg13g2_fill_1 FILLER_45_173 ();
 sg13g2_decap_8 FILLER_45_187 ();
 sg13g2_decap_4 FILLER_45_194 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_45_216 ();
 sg13g2_fill_2 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_decap_4 FILLER_45_398 ();
 sg13g2_fill_1 FILLER_45_415 ();
 sg13g2_decap_4 FILLER_45_421 ();
 sg13g2_decap_4 FILLER_45_430 ();
 sg13g2_fill_1 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_440 ();
 sg13g2_fill_1 FILLER_45_447 ();
 sg13g2_fill_2 FILLER_45_490 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_fill_2 FILLER_45_552 ();
 sg13g2_fill_2 FILLER_45_563 ();
 sg13g2_fill_1 FILLER_45_565 ();
 sg13g2_fill_2 FILLER_45_584 ();
 sg13g2_fill_1 FILLER_45_643 ();
 sg13g2_fill_1 FILLER_45_685 ();
 sg13g2_fill_1 FILLER_45_709 ();
 sg13g2_fill_1 FILLER_45_727 ();
 sg13g2_fill_2 FILLER_45_765 ();
 sg13g2_fill_1 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_4 FILLER_45_857 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_fill_2 FILLER_46_40 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_fill_2 FILLER_46_50 ();
 sg13g2_fill_1 FILLER_46_52 ();
 sg13g2_fill_1 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_117 ();
 sg13g2_fill_1 FILLER_46_144 ();
 sg13g2_decap_4 FILLER_46_176 ();
 sg13g2_fill_1 FILLER_46_212 ();
 sg13g2_decap_4 FILLER_46_223 ();
 sg13g2_fill_2 FILLER_46_227 ();
 sg13g2_decap_4 FILLER_46_232 ();
 sg13g2_fill_1 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_260 ();
 sg13g2_fill_2 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_300 ();
 sg13g2_fill_2 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_fill_2 FILLER_46_356 ();
 sg13g2_fill_2 FILLER_46_379 ();
 sg13g2_fill_1 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_fill_2 FILLER_46_395 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_411 ();
 sg13g2_fill_2 FILLER_46_425 ();
 sg13g2_fill_1 FILLER_46_466 ();
 sg13g2_fill_2 FILLER_46_494 ();
 sg13g2_fill_1 FILLER_46_496 ();
 sg13g2_decap_4 FILLER_46_510 ();
 sg13g2_fill_2 FILLER_46_514 ();
 sg13g2_fill_2 FILLER_46_575 ();
 sg13g2_fill_2 FILLER_46_592 ();
 sg13g2_fill_1 FILLER_46_603 ();
 sg13g2_fill_1 FILLER_46_613 ();
 sg13g2_decap_4 FILLER_46_654 ();
 sg13g2_fill_2 FILLER_46_662 ();
 sg13g2_fill_1 FILLER_46_677 ();
 sg13g2_fill_2 FILLER_46_711 ();
 sg13g2_fill_1 FILLER_46_713 ();
 sg13g2_fill_2 FILLER_46_760 ();
 sg13g2_fill_2 FILLER_46_767 ();
 sg13g2_fill_2 FILLER_46_774 ();
 sg13g2_fill_1 FILLER_46_776 ();
 sg13g2_fill_1 FILLER_46_804 ();
 sg13g2_fill_2 FILLER_46_816 ();
 sg13g2_fill_2 FILLER_46_827 ();
 sg13g2_fill_1 FILLER_46_829 ();
 sg13g2_decap_4 FILLER_46_858 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_4 ();
 sg13g2_fill_2 FILLER_47_9 ();
 sg13g2_fill_1 FILLER_47_11 ();
 sg13g2_decap_4 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_fill_1 FILLER_47_71 ();
 sg13g2_fill_1 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_110 ();
 sg13g2_fill_1 FILLER_47_112 ();
 sg13g2_fill_2 FILLER_47_122 ();
 sg13g2_fill_1 FILLER_47_124 ();
 sg13g2_fill_2 FILLER_47_141 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_decap_8 FILLER_47_174 ();
 sg13g2_fill_2 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_201 ();
 sg13g2_fill_2 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_301 ();
 sg13g2_decap_4 FILLER_47_316 ();
 sg13g2_decap_8 FILLER_47_325 ();
 sg13g2_fill_2 FILLER_47_332 ();
 sg13g2_fill_1 FILLER_47_334 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_decap_4 FILLER_47_360 ();
 sg13g2_fill_2 FILLER_47_379 ();
 sg13g2_fill_1 FILLER_47_381 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_decap_8 FILLER_47_410 ();
 sg13g2_decap_4 FILLER_47_417 ();
 sg13g2_fill_2 FILLER_47_421 ();
 sg13g2_decap_4 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_47_436 ();
 sg13g2_decap_4 FILLER_47_443 ();
 sg13g2_fill_1 FILLER_47_447 ();
 sg13g2_fill_1 FILLER_47_479 ();
 sg13g2_decap_4 FILLER_47_490 ();
 sg13g2_decap_4 FILLER_47_520 ();
 sg13g2_fill_2 FILLER_47_539 ();
 sg13g2_fill_2 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_566 ();
 sg13g2_fill_2 FILLER_47_573 ();
 sg13g2_fill_1 FILLER_47_581 ();
 sg13g2_fill_1 FILLER_47_634 ();
 sg13g2_fill_2 FILLER_47_691 ();
 sg13g2_fill_1 FILLER_47_693 ();
 sg13g2_fill_2 FILLER_47_700 ();
 sg13g2_fill_1 FILLER_47_702 ();
 sg13g2_decap_8 FILLER_47_712 ();
 sg13g2_fill_1 FILLER_47_732 ();
 sg13g2_fill_1 FILLER_47_773 ();
 sg13g2_fill_2 FILLER_47_789 ();
 sg13g2_fill_2 FILLER_47_810 ();
 sg13g2_fill_1 FILLER_47_812 ();
 sg13g2_fill_2 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_32 ();
 sg13g2_decap_4 FILLER_48_47 ();
 sg13g2_decap_4 FILLER_48_106 ();
 sg13g2_fill_2 FILLER_48_114 ();
 sg13g2_fill_1 FILLER_48_120 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_169 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_231 ();
 sg13g2_decap_4 FILLER_48_277 ();
 sg13g2_fill_1 FILLER_48_359 ();
 sg13g2_decap_8 FILLER_48_466 ();
 sg13g2_decap_4 FILLER_48_473 ();
 sg13g2_fill_2 FILLER_48_477 ();
 sg13g2_fill_2 FILLER_48_507 ();
 sg13g2_fill_2 FILLER_48_537 ();
 sg13g2_decap_4 FILLER_48_544 ();
 sg13g2_fill_1 FILLER_48_548 ();
 sg13g2_fill_1 FILLER_48_554 ();
 sg13g2_fill_2 FILLER_48_561 ();
 sg13g2_fill_1 FILLER_48_579 ();
 sg13g2_fill_2 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_597 ();
 sg13g2_fill_1 FILLER_48_618 ();
 sg13g2_decap_8 FILLER_48_648 ();
 sg13g2_decap_4 FILLER_48_655 ();
 sg13g2_fill_2 FILLER_48_659 ();
 sg13g2_decap_8 FILLER_48_675 ();
 sg13g2_fill_1 FILLER_48_682 ();
 sg13g2_fill_2 FILLER_48_692 ();
 sg13g2_decap_4 FILLER_48_703 ();
 sg13g2_fill_2 FILLER_48_716 ();
 sg13g2_fill_1 FILLER_48_752 ();
 sg13g2_fill_2 FILLER_48_793 ();
 sg13g2_fill_2 FILLER_48_832 ();
 sg13g2_fill_1 FILLER_49_27 ();
 sg13g2_fill_2 FILLER_49_33 ();
 sg13g2_fill_2 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_110 ();
 sg13g2_decap_4 FILLER_49_143 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_197 ();
 sg13g2_fill_1 FILLER_49_203 ();
 sg13g2_fill_1 FILLER_49_235 ();
 sg13g2_decap_4 FILLER_49_254 ();
 sg13g2_fill_2 FILLER_49_258 ();
 sg13g2_fill_2 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_4 FILLER_49_329 ();
 sg13g2_fill_2 FILLER_49_333 ();
 sg13g2_fill_2 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_8 FILLER_49_411 ();
 sg13g2_fill_1 FILLER_49_418 ();
 sg13g2_fill_2 FILLER_49_437 ();
 sg13g2_fill_1 FILLER_49_474 ();
 sg13g2_fill_2 FILLER_49_508 ();
 sg13g2_fill_1 FILLER_49_525 ();
 sg13g2_decap_4 FILLER_49_550 ();
 sg13g2_fill_2 FILLER_49_564 ();
 sg13g2_fill_1 FILLER_49_566 ();
 sg13g2_fill_1 FILLER_49_603 ();
 sg13g2_fill_2 FILLER_49_625 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_decap_4 FILLER_49_649 ();
 sg13g2_fill_1 FILLER_49_666 ();
 sg13g2_decap_8 FILLER_49_680 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_793 ();
 sg13g2_fill_1 FILLER_49_811 ();
 sg13g2_fill_2 FILLER_49_816 ();
 sg13g2_fill_1 FILLER_49_818 ();
 sg13g2_fill_2 FILLER_49_832 ();
 sg13g2_fill_1 FILLER_49_834 ();
 sg13g2_decap_4 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_11 ();
 sg13g2_fill_1 FILLER_50_15 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_100 ();
 sg13g2_fill_1 FILLER_50_102 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_fill_2 FILLER_50_119 ();
 sg13g2_fill_1 FILLER_50_121 ();
 sg13g2_decap_4 FILLER_50_139 ();
 sg13g2_decap_8 FILLER_50_156 ();
 sg13g2_decap_4 FILLER_50_163 ();
 sg13g2_decap_4 FILLER_50_220 ();
 sg13g2_fill_2 FILLER_50_224 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_fill_1 FILLER_50_261 ();
 sg13g2_decap_4 FILLER_50_283 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_fill_1 FILLER_50_320 ();
 sg13g2_fill_1 FILLER_50_331 ();
 sg13g2_decap_4 FILLER_50_349 ();
 sg13g2_fill_2 FILLER_50_353 ();
 sg13g2_fill_2 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_395 ();
 sg13g2_fill_1 FILLER_50_397 ();
 sg13g2_fill_1 FILLER_50_438 ();
 sg13g2_fill_2 FILLER_50_471 ();
 sg13g2_fill_1 FILLER_50_473 ();
 sg13g2_fill_2 FILLER_50_502 ();
 sg13g2_fill_1 FILLER_50_504 ();
 sg13g2_fill_2 FILLER_50_539 ();
 sg13g2_fill_1 FILLER_50_541 ();
 sg13g2_fill_2 FILLER_50_548 ();
 sg13g2_fill_1 FILLER_50_550 ();
 sg13g2_fill_1 FILLER_50_556 ();
 sg13g2_fill_1 FILLER_50_574 ();
 sg13g2_decap_4 FILLER_50_581 ();
 sg13g2_fill_2 FILLER_50_585 ();
 sg13g2_fill_1 FILLER_50_591 ();
 sg13g2_decap_4 FILLER_50_596 ();
 sg13g2_fill_1 FILLER_50_616 ();
 sg13g2_fill_1 FILLER_50_621 ();
 sg13g2_fill_2 FILLER_50_640 ();
 sg13g2_decap_8 FILLER_50_656 ();
 sg13g2_fill_2 FILLER_50_695 ();
 sg13g2_decap_4 FILLER_50_701 ();
 sg13g2_fill_1 FILLER_50_705 ();
 sg13g2_decap_4 FILLER_50_711 ();
 sg13g2_fill_2 FILLER_50_715 ();
 sg13g2_fill_2 FILLER_50_736 ();
 sg13g2_fill_1 FILLER_50_738 ();
 sg13g2_decap_4 FILLER_50_755 ();
 sg13g2_fill_2 FILLER_50_759 ();
 sg13g2_fill_2 FILLER_50_778 ();
 sg13g2_decap_8 FILLER_50_787 ();
 sg13g2_fill_2 FILLER_50_794 ();
 sg13g2_fill_1 FILLER_50_796 ();
 sg13g2_fill_2 FILLER_50_802 ();
 sg13g2_fill_2 FILLER_50_809 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_fill_2 FILLER_50_826 ();
 sg13g2_fill_1 FILLER_50_828 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_30 ();
 sg13g2_decap_8 FILLER_51_45 ();
 sg13g2_decap_4 FILLER_51_52 ();
 sg13g2_fill_2 FILLER_51_69 ();
 sg13g2_fill_1 FILLER_51_71 ();
 sg13g2_decap_4 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_121 ();
 sg13g2_decap_8 FILLER_51_153 ();
 sg13g2_fill_2 FILLER_51_160 ();
 sg13g2_decap_4 FILLER_51_166 ();
 sg13g2_fill_1 FILLER_51_170 ();
 sg13g2_fill_1 FILLER_51_202 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_255 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_decap_8 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_51_354 ();
 sg13g2_decap_4 FILLER_51_397 ();
 sg13g2_fill_1 FILLER_51_401 ();
 sg13g2_fill_2 FILLER_51_460 ();
 sg13g2_fill_1 FILLER_51_462 ();
 sg13g2_fill_1 FILLER_51_468 ();
 sg13g2_fill_1 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_493 ();
 sg13g2_fill_1 FILLER_51_495 ();
 sg13g2_fill_2 FILLER_51_505 ();
 sg13g2_decap_8 FILLER_51_599 ();
 sg13g2_decap_4 FILLER_51_649 ();
 sg13g2_decap_8 FILLER_51_659 ();
 sg13g2_fill_2 FILLER_51_706 ();
 sg13g2_fill_1 FILLER_51_708 ();
 sg13g2_fill_2 FILLER_51_759 ();
 sg13g2_fill_2 FILLER_51_779 ();
 sg13g2_fill_2 FILLER_51_793 ();
 sg13g2_decap_4 FILLER_51_820 ();
 sg13g2_fill_1 FILLER_51_824 ();
 sg13g2_decap_4 FILLER_51_830 ();
 sg13g2_fill_2 FILLER_51_834 ();
 sg13g2_fill_1 FILLER_51_852 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_34 ();
 sg13g2_fill_2 FILLER_52_66 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_fill_2 FILLER_52_93 ();
 sg13g2_fill_2 FILLER_52_102 ();
 sg13g2_fill_1 FILLER_52_117 ();
 sg13g2_decap_4 FILLER_52_151 ();
 sg13g2_fill_2 FILLER_52_155 ();
 sg13g2_decap_4 FILLER_52_226 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_fill_2 FILLER_52_271 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_315 ();
 sg13g2_fill_1 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_327 ();
 sg13g2_fill_1 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_410 ();
 sg13g2_decap_4 FILLER_52_417 ();
 sg13g2_decap_4 FILLER_52_434 ();
 sg13g2_fill_2 FILLER_52_438 ();
 sg13g2_fill_1 FILLER_52_453 ();
 sg13g2_fill_2 FILLER_52_510 ();
 sg13g2_fill_2 FILLER_52_566 ();
 sg13g2_fill_1 FILLER_52_587 ();
 sg13g2_fill_1 FILLER_52_631 ();
 sg13g2_decap_8 FILLER_52_658 ();
 sg13g2_fill_2 FILLER_52_665 ();
 sg13g2_fill_1 FILLER_52_667 ();
 sg13g2_decap_8 FILLER_52_681 ();
 sg13g2_fill_2 FILLER_52_688 ();
 sg13g2_fill_1 FILLER_52_744 ();
 sg13g2_fill_2 FILLER_52_770 ();
 sg13g2_fill_1 FILLER_52_781 ();
 sg13g2_fill_2 FILLER_52_787 ();
 sg13g2_fill_1 FILLER_52_789 ();
 sg13g2_decap_8 FILLER_52_794 ();
 sg13g2_fill_2 FILLER_52_824 ();
 sg13g2_fill_1 FILLER_52_834 ();
 sg13g2_fill_2 FILLER_52_844 ();
 sg13g2_decap_8 FILLER_52_851 ();
 sg13g2_decap_4 FILLER_52_858 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_42 ();
 sg13g2_fill_1 FILLER_53_80 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_decap_4 FILLER_53_162 ();
 sg13g2_fill_1 FILLER_53_194 ();
 sg13g2_decap_4 FILLER_53_248 ();
 sg13g2_fill_1 FILLER_53_303 ();
 sg13g2_fill_2 FILLER_53_323 ();
 sg13g2_fill_2 FILLER_53_331 ();
 sg13g2_fill_2 FILLER_53_356 ();
 sg13g2_fill_1 FILLER_53_358 ();
 sg13g2_fill_2 FILLER_53_373 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_fill_1 FILLER_53_387 ();
 sg13g2_decap_4 FILLER_53_407 ();
 sg13g2_fill_1 FILLER_53_411 ();
 sg13g2_decap_4 FILLER_53_440 ();
 sg13g2_fill_2 FILLER_53_480 ();
 sg13g2_fill_1 FILLER_53_488 ();
 sg13g2_fill_2 FILLER_53_539 ();
 sg13g2_fill_2 FILLER_53_550 ();
 sg13g2_fill_1 FILLER_53_565 ();
 sg13g2_fill_2 FILLER_53_594 ();
 sg13g2_decap_4 FILLER_53_605 ();
 sg13g2_fill_1 FILLER_53_609 ();
 sg13g2_fill_2 FILLER_53_636 ();
 sg13g2_fill_1 FILLER_53_638 ();
 sg13g2_fill_2 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_720 ();
 sg13g2_fill_2 FILLER_53_769 ();
 sg13g2_fill_1 FILLER_53_799 ();
 sg13g2_decap_4 FILLER_53_813 ();
 sg13g2_fill_2 FILLER_53_817 ();
 sg13g2_fill_2 FILLER_53_823 ();
 sg13g2_fill_1 FILLER_53_825 ();
 sg13g2_decap_4 FILLER_53_829 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_fill_2 FILLER_54_59 ();
 sg13g2_fill_1 FILLER_54_61 ();
 sg13g2_fill_1 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_163 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_fill_2 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_fill_2 FILLER_54_227 ();
 sg13g2_decap_8 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_251 ();
 sg13g2_fill_2 FILLER_54_265 ();
 sg13g2_fill_2 FILLER_54_275 ();
 sg13g2_fill_2 FILLER_54_296 ();
 sg13g2_fill_1 FILLER_54_298 ();
 sg13g2_decap_4 FILLER_54_303 ();
 sg13g2_fill_1 FILLER_54_356 ();
 sg13g2_decap_4 FILLER_54_390 ();
 sg13g2_fill_1 FILLER_54_394 ();
 sg13g2_decap_8 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_54_424 ();
 sg13g2_decap_8 FILLER_54_468 ();
 sg13g2_fill_2 FILLER_54_518 ();
 sg13g2_fill_2 FILLER_54_562 ();
 sg13g2_fill_1 FILLER_54_564 ();
 sg13g2_decap_4 FILLER_54_587 ();
 sg13g2_fill_1 FILLER_54_591 ();
 sg13g2_fill_2 FILLER_54_607 ();
 sg13g2_fill_1 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_653 ();
 sg13g2_fill_2 FILLER_54_660 ();
 sg13g2_decap_4 FILLER_54_679 ();
 sg13g2_fill_2 FILLER_54_735 ();
 sg13g2_fill_2 FILLER_54_750 ();
 sg13g2_fill_1 FILLER_54_752 ();
 sg13g2_fill_1 FILLER_54_769 ();
 sg13g2_decap_8 FILLER_54_773 ();
 sg13g2_fill_1 FILLER_54_784 ();
 sg13g2_decap_4 FILLER_54_798 ();
 sg13g2_fill_2 FILLER_54_807 ();
 sg13g2_fill_1 FILLER_54_809 ();
 sg13g2_decap_8 FILLER_54_823 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_fill_1 FILLER_55_27 ();
 sg13g2_fill_1 FILLER_55_37 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_fill_2 FILLER_55_127 ();
 sg13g2_fill_2 FILLER_55_147 ();
 sg13g2_decap_4 FILLER_55_172 ();
 sg13g2_fill_2 FILLER_55_176 ();
 sg13g2_decap_4 FILLER_55_210 ();
 sg13g2_decap_4 FILLER_55_250 ();
 sg13g2_fill_2 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_fill_2 FILLER_55_360 ();
 sg13g2_decap_8 FILLER_55_375 ();
 sg13g2_decap_8 FILLER_55_382 ();
 sg13g2_fill_1 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_426 ();
 sg13g2_decap_8 FILLER_55_433 ();
 sg13g2_fill_2 FILLER_55_440 ();
 sg13g2_fill_1 FILLER_55_442 ();
 sg13g2_decap_8 FILLER_55_452 ();
 sg13g2_decap_4 FILLER_55_468 ();
 sg13g2_fill_1 FILLER_55_472 ();
 sg13g2_fill_2 FILLER_55_550 ();
 sg13g2_fill_1 FILLER_55_552 ();
 sg13g2_fill_2 FILLER_55_570 ();
 sg13g2_fill_1 FILLER_55_572 ();
 sg13g2_fill_2 FILLER_55_583 ();
 sg13g2_decap_8 FILLER_55_596 ();
 sg13g2_fill_2 FILLER_55_603 ();
 sg13g2_fill_1 FILLER_55_605 ();
 sg13g2_decap_4 FILLER_55_633 ();
 sg13g2_fill_1 FILLER_55_687 ();
 sg13g2_fill_2 FILLER_55_701 ();
 sg13g2_decap_8 FILLER_55_707 ();
 sg13g2_fill_2 FILLER_55_755 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_4 FILLER_55_784 ();
 sg13g2_fill_2 FILLER_55_788 ();
 sg13g2_decap_4 FILLER_55_794 ();
 sg13g2_fill_2 FILLER_55_803 ();
 sg13g2_fill_1 FILLER_55_805 ();
 sg13g2_fill_2 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_fill_2 FILLER_55_835 ();
 sg13g2_fill_1 FILLER_55_837 ();
 sg13g2_decap_8 FILLER_55_848 ();
 sg13g2_decap_8 FILLER_55_855 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_4 ();
 sg13g2_fill_2 FILLER_56_9 ();
 sg13g2_fill_1 FILLER_56_11 ();
 sg13g2_fill_1 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_187 ();
 sg13g2_fill_1 FILLER_56_189 ();
 sg13g2_decap_4 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_199 ();
 sg13g2_decap_4 FILLER_56_203 ();
 sg13g2_fill_1 FILLER_56_207 ();
 sg13g2_fill_1 FILLER_56_229 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_decap_8 FILLER_56_267 ();
 sg13g2_fill_2 FILLER_56_274 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_fill_2 FILLER_56_301 ();
 sg13g2_fill_1 FILLER_56_303 ();
 sg13g2_fill_1 FILLER_56_313 ();
 sg13g2_fill_2 FILLER_56_348 ();
 sg13g2_fill_1 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_362 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_378 ();
 sg13g2_fill_2 FILLER_56_421 ();
 sg13g2_fill_1 FILLER_56_423 ();
 sg13g2_fill_2 FILLER_56_443 ();
 sg13g2_fill_1 FILLER_56_445 ();
 sg13g2_decap_8 FILLER_56_454 ();
 sg13g2_fill_2 FILLER_56_515 ();
 sg13g2_fill_1 FILLER_56_517 ();
 sg13g2_fill_2 FILLER_56_524 ();
 sg13g2_fill_1 FILLER_56_526 ();
 sg13g2_fill_2 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_573 ();
 sg13g2_fill_1 FILLER_56_606 ();
 sg13g2_fill_2 FILLER_56_613 ();
 sg13g2_fill_1 FILLER_56_615 ();
 sg13g2_fill_2 FILLER_56_644 ();
 sg13g2_fill_1 FILLER_56_646 ();
 sg13g2_fill_2 FILLER_56_664 ();
 sg13g2_fill_1 FILLER_56_666 ();
 sg13g2_fill_2 FILLER_56_700 ();
 sg13g2_fill_1 FILLER_56_702 ();
 sg13g2_decap_8 FILLER_56_708 ();
 sg13g2_fill_2 FILLER_56_715 ();
 sg13g2_fill_1 FILLER_56_721 ();
 sg13g2_decap_8 FILLER_56_730 ();
 sg13g2_decap_4 FILLER_56_737 ();
 sg13g2_fill_2 FILLER_56_741 ();
 sg13g2_fill_2 FILLER_56_750 ();
 sg13g2_fill_1 FILLER_56_752 ();
 sg13g2_decap_4 FILLER_56_757 ();
 sg13g2_fill_1 FILLER_56_761 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_decap_4 FILLER_56_774 ();
 sg13g2_fill_2 FILLER_56_787 ();
 sg13g2_fill_2 FILLER_56_793 ();
 sg13g2_fill_1 FILLER_56_811 ();
 sg13g2_fill_2 FILLER_56_833 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_43 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_1 FILLER_57_99 ();
 sg13g2_fill_1 FILLER_57_116 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_decap_8 FILLER_57_246 ();
 sg13g2_decap_4 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_257 ();
 sg13g2_fill_2 FILLER_57_287 ();
 sg13g2_fill_1 FILLER_57_289 ();
 sg13g2_decap_4 FILLER_57_345 ();
 sg13g2_fill_2 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_386 ();
 sg13g2_fill_2 FILLER_57_409 ();
 sg13g2_fill_1 FILLER_57_411 ();
 sg13g2_decap_4 FILLER_57_429 ();
 sg13g2_fill_1 FILLER_57_469 ();
 sg13g2_fill_1 FILLER_57_504 ();
 sg13g2_decap_4 FILLER_57_510 ();
 sg13g2_fill_2 FILLER_57_514 ();
 sg13g2_decap_8 FILLER_57_571 ();
 sg13g2_decap_8 FILLER_57_578 ();
 sg13g2_fill_2 FILLER_57_585 ();
 sg13g2_fill_1 FILLER_57_587 ();
 sg13g2_decap_8 FILLER_57_598 ();
 sg13g2_fill_1 FILLER_57_605 ();
 sg13g2_decap_8 FILLER_57_632 ();
 sg13g2_decap_8 FILLER_57_657 ();
 sg13g2_fill_2 FILLER_57_664 ();
 sg13g2_fill_1 FILLER_57_666 ();
 sg13g2_fill_1 FILLER_57_680 ();
 sg13g2_fill_1 FILLER_57_698 ();
 sg13g2_decap_8 FILLER_57_719 ();
 sg13g2_decap_4 FILLER_57_726 ();
 sg13g2_fill_2 FILLER_57_730 ();
 sg13g2_decap_8 FILLER_57_752 ();
 sg13g2_decap_4 FILLER_57_759 ();
 sg13g2_fill_1 FILLER_57_771 ();
 sg13g2_fill_2 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_804 ();
 sg13g2_decap_8 FILLER_57_820 ();
 sg13g2_decap_8 FILLER_57_827 ();
 sg13g2_decap_4 FILLER_57_834 ();
 sg13g2_fill_1 FILLER_57_838 ();
 sg13g2_fill_1 FILLER_57_843 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_4 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_decap_8 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_192 ();
 sg13g2_decap_4 FILLER_58_198 ();
 sg13g2_fill_1 FILLER_58_202 ();
 sg13g2_fill_2 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_218 ();
 sg13g2_decap_4 FILLER_58_223 ();
 sg13g2_decap_8 FILLER_58_230 ();
 sg13g2_decap_4 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_250 ();
 sg13g2_fill_2 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_303 ();
 sg13g2_decap_4 FILLER_58_328 ();
 sg13g2_decap_4 FILLER_58_348 ();
 sg13g2_fill_2 FILLER_58_352 ();
 sg13g2_fill_2 FILLER_58_373 ();
 sg13g2_fill_1 FILLER_58_375 ();
 sg13g2_decap_4 FILLER_58_382 ();
 sg13g2_fill_2 FILLER_58_392 ();
 sg13g2_fill_2 FILLER_58_412 ();
 sg13g2_decap_4 FILLER_58_423 ();
 sg13g2_fill_1 FILLER_58_427 ();
 sg13g2_decap_8 FILLER_58_433 ();
 sg13g2_decap_4 FILLER_58_440 ();
 sg13g2_fill_1 FILLER_58_448 ();
 sg13g2_fill_2 FILLER_58_455 ();
 sg13g2_fill_1 FILLER_58_457 ();
 sg13g2_fill_1 FILLER_58_473 ();
 sg13g2_decap_4 FILLER_58_483 ();
 sg13g2_decap_8 FILLER_58_518 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_fill_2 FILLER_58_532 ();
 sg13g2_decap_4 FILLER_58_538 ();
 sg13g2_fill_2 FILLER_58_542 ();
 sg13g2_fill_2 FILLER_58_550 ();
 sg13g2_fill_1 FILLER_58_552 ();
 sg13g2_fill_2 FILLER_58_564 ();
 sg13g2_fill_2 FILLER_58_572 ();
 sg13g2_decap_4 FILLER_58_591 ();
 sg13g2_fill_1 FILLER_58_599 ();
 sg13g2_fill_2 FILLER_58_616 ();
 sg13g2_fill_1 FILLER_58_624 ();
 sg13g2_decap_8 FILLER_58_638 ();
 sg13g2_decap_8 FILLER_58_645 ();
 sg13g2_decap_4 FILLER_58_652 ();
 sg13g2_fill_2 FILLER_58_656 ();
 sg13g2_decap_8 FILLER_58_662 ();
 sg13g2_decap_8 FILLER_58_669 ();
 sg13g2_fill_2 FILLER_58_676 ();
 sg13g2_fill_1 FILLER_58_678 ();
 sg13g2_fill_1 FILLER_58_700 ();
 sg13g2_fill_2 FILLER_58_741 ();
 sg13g2_fill_1 FILLER_58_743 ();
 sg13g2_fill_2 FILLER_58_754 ();
 sg13g2_fill_1 FILLER_58_756 ();
 sg13g2_decap_4 FILLER_58_775 ();
 sg13g2_fill_2 FILLER_58_779 ();
 sg13g2_fill_2 FILLER_58_785 ();
 sg13g2_fill_1 FILLER_58_787 ();
 sg13g2_fill_2 FILLER_58_793 ();
 sg13g2_fill_1 FILLER_58_800 ();
 sg13g2_fill_1 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_823 ();
 sg13g2_fill_1 FILLER_58_830 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_33 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_decap_4 FILLER_59_93 ();
 sg13g2_fill_2 FILLER_59_97 ();
 sg13g2_fill_2 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_173 ();
 sg13g2_fill_1 FILLER_59_175 ();
 sg13g2_fill_1 FILLER_59_204 ();
 sg13g2_fill_2 FILLER_59_269 ();
 sg13g2_fill_2 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_301 ();
 sg13g2_decap_4 FILLER_59_323 ();
 sg13g2_decap_8 FILLER_59_347 ();
 sg13g2_fill_1 FILLER_59_354 ();
 sg13g2_decap_4 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_412 ();
 sg13g2_fill_1 FILLER_59_414 ();
 sg13g2_fill_1 FILLER_59_482 ();
 sg13g2_fill_1 FILLER_59_505 ();
 sg13g2_fill_2 FILLER_59_523 ();
 sg13g2_fill_1 FILLER_59_562 ();
 sg13g2_fill_1 FILLER_59_574 ();
 sg13g2_decap_4 FILLER_59_590 ();
 sg13g2_fill_1 FILLER_59_600 ();
 sg13g2_fill_2 FILLER_59_615 ();
 sg13g2_fill_2 FILLER_59_686 ();
 sg13g2_fill_1 FILLER_59_698 ();
 sg13g2_fill_2 FILLER_59_709 ();
 sg13g2_fill_1 FILLER_59_711 ();
 sg13g2_decap_8 FILLER_59_733 ();
 sg13g2_decap_4 FILLER_59_740 ();
 sg13g2_fill_1 FILLER_59_762 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_decap_4 FILLER_59_773 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_fill_2 FILLER_59_812 ();
 sg13g2_fill_2 FILLER_59_818 ();
 sg13g2_decap_4 FILLER_59_840 ();
 sg13g2_fill_1 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_853 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_fill_1 FILLER_60_47 ();
 sg13g2_fill_2 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_178 ();
 sg13g2_decap_4 FILLER_60_185 ();
 sg13g2_fill_2 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_195 ();
 sg13g2_decap_8 FILLER_60_202 ();
 sg13g2_decap_8 FILLER_60_209 ();
 sg13g2_fill_1 FILLER_60_216 ();
 sg13g2_decap_8 FILLER_60_225 ();
 sg13g2_decap_8 FILLER_60_232 ();
 sg13g2_decap_8 FILLER_60_243 ();
 sg13g2_fill_2 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_284 ();
 sg13g2_fill_2 FILLER_60_326 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_fill_1 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_430 ();
 sg13g2_decap_4 FILLER_60_437 ();
 sg13g2_fill_1 FILLER_60_441 ();
 sg13g2_fill_1 FILLER_60_479 ();
 sg13g2_fill_2 FILLER_60_514 ();
 sg13g2_fill_1 FILLER_60_516 ();
 sg13g2_fill_2 FILLER_60_534 ();
 sg13g2_fill_2 FILLER_60_550 ();
 sg13g2_fill_1 FILLER_60_552 ();
 sg13g2_fill_2 FILLER_60_586 ();
 sg13g2_fill_1 FILLER_60_588 ();
 sg13g2_decap_4 FILLER_60_614 ();
 sg13g2_fill_2 FILLER_60_618 ();
 sg13g2_fill_2 FILLER_60_629 ();
 sg13g2_decap_8 FILLER_60_644 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_fill_2 FILLER_60_665 ();
 sg13g2_decap_8 FILLER_60_675 ();
 sg13g2_fill_2 FILLER_60_682 ();
 sg13g2_fill_2 FILLER_60_705 ();
 sg13g2_fill_1 FILLER_60_707 ();
 sg13g2_decap_4 FILLER_60_741 ();
 sg13g2_fill_2 FILLER_60_745 ();
 sg13g2_fill_1 FILLER_60_767 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_4 FILLER_60_787 ();
 sg13g2_fill_1 FILLER_60_791 ();
 sg13g2_decap_8 FILLER_60_797 ();
 sg13g2_fill_2 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_fill_1 FILLER_60_835 ();
 sg13g2_fill_1 FILLER_60_844 ();
 sg13g2_decap_4 FILLER_60_858 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_decap_8 FILLER_61_9 ();
 sg13g2_fill_1 FILLER_61_16 ();
 sg13g2_decap_4 FILLER_61_49 ();
 sg13g2_fill_2 FILLER_61_57 ();
 sg13g2_fill_1 FILLER_61_59 ();
 sg13g2_decap_4 FILLER_61_97 ();
 sg13g2_fill_2 FILLER_61_171 ();
 sg13g2_fill_2 FILLER_61_213 ();
 sg13g2_decap_4 FILLER_61_256 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_decap_4 FILLER_61_265 ();
 sg13g2_fill_2 FILLER_61_269 ();
 sg13g2_fill_2 FILLER_61_280 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_decap_4 FILLER_61_345 ();
 sg13g2_fill_1 FILLER_61_349 ();
 sg13g2_decap_4 FILLER_61_372 ();
 sg13g2_fill_2 FILLER_61_389 ();
 sg13g2_fill_1 FILLER_61_391 ();
 sg13g2_fill_2 FILLER_61_412 ();
 sg13g2_fill_1 FILLER_61_414 ();
 sg13g2_decap_4 FILLER_61_428 ();
 sg13g2_fill_2 FILLER_61_432 ();
 sg13g2_fill_2 FILLER_61_439 ();
 sg13g2_fill_1 FILLER_61_441 ();
 sg13g2_fill_2 FILLER_61_463 ();
 sg13g2_fill_1 FILLER_61_465 ();
 sg13g2_decap_4 FILLER_61_494 ();
 sg13g2_fill_2 FILLER_61_498 ();
 sg13g2_fill_2 FILLER_61_518 ();
 sg13g2_decap_4 FILLER_61_557 ();
 sg13g2_fill_1 FILLER_61_573 ();
 sg13g2_fill_1 FILLER_61_602 ();
 sg13g2_fill_1 FILLER_61_609 ();
 sg13g2_fill_1 FILLER_61_637 ();
 sg13g2_fill_2 FILLER_61_718 ();
 sg13g2_fill_1 FILLER_61_720 ();
 sg13g2_decap_8 FILLER_61_748 ();
 sg13g2_fill_2 FILLER_61_755 ();
 sg13g2_fill_1 FILLER_61_757 ();
 sg13g2_decap_8 FILLER_61_773 ();
 sg13g2_fill_2 FILLER_61_780 ();
 sg13g2_decap_4 FILLER_61_795 ();
 sg13g2_decap_8 FILLER_61_804 ();
 sg13g2_decap_4 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_836 ();
 sg13g2_fill_2 FILLER_61_843 ();
 sg13g2_fill_1 FILLER_61_845 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_9 ();
 sg13g2_fill_2 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_16 ();
 sg13g2_fill_2 FILLER_62_36 ();
 sg13g2_fill_2 FILLER_62_43 ();
 sg13g2_fill_1 FILLER_62_45 ();
 sg13g2_decap_4 FILLER_62_59 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_decap_4 FILLER_62_82 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_decap_8 FILLER_62_193 ();
 sg13g2_decap_8 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_207 ();
 sg13g2_fill_2 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_344 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_fill_2 FILLER_62_373 ();
 sg13g2_fill_1 FILLER_62_375 ();
 sg13g2_fill_2 FILLER_62_394 ();
 sg13g2_fill_2 FILLER_62_402 ();
 sg13g2_fill_1 FILLER_62_438 ();
 sg13g2_fill_2 FILLER_62_445 ();
 sg13g2_fill_1 FILLER_62_447 ();
 sg13g2_decap_4 FILLER_62_489 ();
 sg13g2_fill_1 FILLER_62_516 ();
 sg13g2_fill_1 FILLER_62_534 ();
 sg13g2_decap_8 FILLER_62_548 ();
 sg13g2_fill_2 FILLER_62_555 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_fill_2 FILLER_62_650 ();
 sg13g2_fill_1 FILLER_62_652 ();
 sg13g2_fill_2 FILLER_62_666 ();
 sg13g2_fill_1 FILLER_62_668 ();
 sg13g2_fill_2 FILLER_62_682 ();
 sg13g2_fill_1 FILLER_62_684 ();
 sg13g2_fill_1 FILLER_62_707 ();
 sg13g2_fill_2 FILLER_62_717 ();
 sg13g2_fill_1 FILLER_62_719 ();
 sg13g2_fill_2 FILLER_62_756 ();
 sg13g2_fill_1 FILLER_62_758 ();
 sg13g2_fill_2 FILLER_62_767 ();
 sg13g2_decap_8 FILLER_62_786 ();
 sg13g2_decap_4 FILLER_62_793 ();
 sg13g2_fill_1 FILLER_62_797 ();
 sg13g2_decap_8 FILLER_62_814 ();
 sg13g2_fill_2 FILLER_62_821 ();
 sg13g2_decap_4 FILLER_62_834 ();
 sg13g2_fill_2 FILLER_62_838 ();
 sg13g2_fill_1 FILLER_62_844 ();
 sg13g2_decap_4 FILLER_62_858 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_4 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_fill_1 FILLER_63_34 ();
 sg13g2_decap_4 FILLER_63_98 ();
 sg13g2_fill_1 FILLER_63_102 ();
 sg13g2_decap_8 FILLER_63_186 ();
 sg13g2_decap_4 FILLER_63_193 ();
 sg13g2_fill_1 FILLER_63_197 ();
 sg13g2_fill_2 FILLER_63_251 ();
 sg13g2_fill_1 FILLER_63_253 ();
 sg13g2_fill_1 FILLER_63_295 ();
 sg13g2_decap_4 FILLER_63_336 ();
 sg13g2_fill_2 FILLER_63_340 ();
 sg13g2_fill_1 FILLER_63_359 ();
 sg13g2_fill_2 FILLER_63_375 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_fill_2 FILLER_63_391 ();
 sg13g2_fill_2 FILLER_63_424 ();
 sg13g2_fill_1 FILLER_63_432 ();
 sg13g2_fill_2 FILLER_63_438 ();
 sg13g2_fill_1 FILLER_63_440 ();
 sg13g2_fill_2 FILLER_63_445 ();
 sg13g2_fill_1 FILLER_63_447 ();
 sg13g2_fill_2 FILLER_63_471 ();
 sg13g2_fill_2 FILLER_63_478 ();
 sg13g2_fill_1 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_506 ();
 sg13g2_fill_2 FILLER_63_576 ();
 sg13g2_fill_2 FILLER_63_634 ();
 sg13g2_fill_1 FILLER_63_636 ();
 sg13g2_fill_2 FILLER_63_642 ();
 sg13g2_fill_1 FILLER_63_644 ();
 sg13g2_fill_1 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_4 FILLER_63_693 ();
 sg13g2_fill_1 FILLER_63_724 ();
 sg13g2_fill_2 FILLER_63_738 ();
 sg13g2_fill_2 FILLER_63_746 ();
 sg13g2_fill_1 FILLER_63_757 ();
 sg13g2_decap_4 FILLER_63_787 ();
 sg13g2_decap_4 FILLER_63_814 ();
 sg13g2_fill_2 FILLER_63_818 ();
 sg13g2_fill_2 FILLER_63_833 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_4 ();
 sg13g2_fill_1 FILLER_64_42 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_80 ();
 sg13g2_fill_2 FILLER_64_127 ();
 sg13g2_fill_2 FILLER_64_221 ();
 sg13g2_fill_2 FILLER_64_264 ();
 sg13g2_fill_2 FILLER_64_279 ();
 sg13g2_fill_2 FILLER_64_287 ();
 sg13g2_fill_1 FILLER_64_289 ();
 sg13g2_fill_2 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_376 ();
 sg13g2_fill_2 FILLER_64_443 ();
 sg13g2_fill_1 FILLER_64_504 ();
 sg13g2_decap_8 FILLER_64_529 ();
 sg13g2_fill_2 FILLER_64_536 ();
 sg13g2_fill_1 FILLER_64_538 ();
 sg13g2_fill_1 FILLER_64_562 ();
 sg13g2_fill_2 FILLER_64_584 ();
 sg13g2_fill_2 FILLER_64_605 ();
 sg13g2_fill_1 FILLER_64_607 ();
 sg13g2_fill_2 FILLER_64_612 ();
 sg13g2_fill_2 FILLER_64_659 ();
 sg13g2_fill_1 FILLER_64_661 ();
 sg13g2_fill_1 FILLER_64_684 ();
 sg13g2_fill_2 FILLER_64_754 ();
 sg13g2_fill_1 FILLER_64_774 ();
 sg13g2_fill_2 FILLER_64_851 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_fill_2 FILLER_65_63 ();
 sg13g2_fill_2 FILLER_65_79 ();
 sg13g2_fill_1 FILLER_65_107 ();
 sg13g2_fill_2 FILLER_65_170 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_fill_1 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_200 ();
 sg13g2_decap_4 FILLER_65_207 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_2 FILLER_65_252 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_1 FILLER_65_311 ();
 sg13g2_fill_2 FILLER_65_331 ();
 sg13g2_fill_2 FILLER_65_350 ();
 sg13g2_fill_1 FILLER_65_352 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_438 ();
 sg13g2_fill_2 FILLER_65_445 ();
 sg13g2_fill_1 FILLER_65_447 ();
 sg13g2_fill_1 FILLER_65_490 ();
 sg13g2_fill_1 FILLER_65_504 ();
 sg13g2_fill_2 FILLER_65_539 ();
 sg13g2_fill_1 FILLER_65_557 ();
 sg13g2_decap_4 FILLER_65_609 ();
 sg13g2_fill_2 FILLER_65_621 ();
 sg13g2_fill_1 FILLER_65_623 ();
 sg13g2_fill_2 FILLER_65_646 ();
 sg13g2_fill_1 FILLER_65_648 ();
 sg13g2_fill_2 FILLER_65_662 ();
 sg13g2_decap_4 FILLER_65_678 ();
 sg13g2_fill_1 FILLER_65_682 ();
 sg13g2_fill_1 FILLER_65_745 ();
 sg13g2_fill_1 FILLER_65_760 ();
 sg13g2_fill_2 FILLER_65_779 ();
 sg13g2_fill_2 FILLER_65_807 ();
 sg13g2_decap_4 FILLER_65_813 ();
 sg13g2_decap_4 FILLER_65_825 ();
 sg13g2_fill_1 FILLER_65_829 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_90 ();
 sg13g2_fill_2 FILLER_66_119 ();
 sg13g2_fill_2 FILLER_66_146 ();
 sg13g2_fill_1 FILLER_66_148 ();
 sg13g2_fill_2 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_194 ();
 sg13g2_decap_4 FILLER_66_199 ();
 sg13g2_fill_1 FILLER_66_203 ();
 sg13g2_decap_4 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_212 ();
 sg13g2_decap_8 FILLER_66_227 ();
 sg13g2_decap_8 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_269 ();
 sg13g2_fill_2 FILLER_66_292 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_decap_4 FILLER_66_351 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_391 ();
 sg13g2_fill_1 FILLER_66_402 ();
 sg13g2_fill_1 FILLER_66_416 ();
 sg13g2_fill_1 FILLER_66_480 ();
 sg13g2_fill_2 FILLER_66_518 ();
 sg13g2_fill_1 FILLER_66_520 ();
 sg13g2_fill_1 FILLER_66_634 ();
 sg13g2_fill_1 FILLER_66_656 ();
 sg13g2_fill_1 FILLER_66_692 ();
 sg13g2_fill_2 FILLER_66_727 ();
 sg13g2_fill_1 FILLER_66_729 ();
 sg13g2_fill_1 FILLER_66_804 ();
 sg13g2_fill_2 FILLER_66_819 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_113 ();
 sg13g2_fill_2 FILLER_67_126 ();
 sg13g2_fill_1 FILLER_67_128 ();
 sg13g2_fill_2 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_fill_1 FILLER_67_173 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_fill_2 FILLER_67_195 ();
 sg13g2_fill_2 FILLER_67_291 ();
 sg13g2_fill_2 FILLER_67_327 ();
 sg13g2_fill_2 FILLER_67_424 ();
 sg13g2_fill_1 FILLER_67_426 ();
 sg13g2_decap_8 FILLER_67_440 ();
 sg13g2_fill_1 FILLER_67_447 ();
 sg13g2_fill_1 FILLER_67_452 ();
 sg13g2_fill_2 FILLER_67_518 ();
 sg13g2_fill_1 FILLER_67_520 ();
 sg13g2_fill_1 FILLER_67_543 ();
 sg13g2_fill_2 FILLER_67_557 ();
 sg13g2_fill_1 FILLER_67_559 ();
 sg13g2_fill_2 FILLER_67_610 ();
 sg13g2_decap_4 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_620 ();
 sg13g2_fill_2 FILLER_67_640 ();
 sg13g2_fill_2 FILLER_67_681 ();
 sg13g2_fill_1 FILLER_67_683 ();
 sg13g2_fill_2 FILLER_67_693 ();
 sg13g2_fill_1 FILLER_67_695 ();
 sg13g2_fill_1 FILLER_67_706 ();
 sg13g2_fill_1 FILLER_67_728 ();
 sg13g2_fill_2 FILLER_67_778 ();
 sg13g2_fill_1 FILLER_67_780 ();
 sg13g2_decap_4 FILLER_67_845 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_1 FILLER_68_56 ();
 sg13g2_decap_4 FILLER_68_201 ();
 sg13g2_decap_8 FILLER_68_209 ();
 sg13g2_decap_4 FILLER_68_216 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_2 FILLER_68_266 ();
 sg13g2_fill_1 FILLER_68_268 ();
 sg13g2_fill_1 FILLER_68_345 ();
 sg13g2_fill_2 FILLER_68_355 ();
 sg13g2_decap_4 FILLER_68_421 ();
 sg13g2_fill_2 FILLER_68_425 ();
 sg13g2_fill_1 FILLER_68_432 ();
 sg13g2_fill_2 FILLER_68_511 ();
 sg13g2_fill_1 FILLER_68_513 ();
 sg13g2_fill_2 FILLER_68_583 ();
 sg13g2_fill_1 FILLER_68_585 ();
 sg13g2_fill_2 FILLER_68_610 ();
 sg13g2_fill_1 FILLER_68_612 ();
 sg13g2_fill_2 FILLER_68_623 ();
 sg13g2_fill_2 FILLER_68_630 ();
 sg13g2_fill_2 FILLER_68_702 ();
 sg13g2_fill_1 FILLER_68_704 ();
 sg13g2_fill_1 FILLER_68_723 ();
 sg13g2_fill_2 FILLER_68_790 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_fill_1 FILLER_68_803 ();
 sg13g2_decap_4 FILLER_68_808 ();
 sg13g2_decap_4 FILLER_68_817 ();
 sg13g2_fill_2 FILLER_68_825 ();
 sg13g2_fill_2 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_41 ();
 sg13g2_fill_1 FILLER_69_43 ();
 sg13g2_fill_2 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_55 ();
 sg13g2_decap_4 FILLER_69_101 ();
 sg13g2_decap_4 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_136 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_181 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_227 ();
 sg13g2_fill_1 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_250 ();
 sg13g2_fill_1 FILLER_69_270 ();
 sg13g2_fill_1 FILLER_69_280 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_fill_2 FILLER_69_295 ();
 sg13g2_fill_1 FILLER_69_297 ();
 sg13g2_fill_1 FILLER_69_324 ();
 sg13g2_fill_2 FILLER_69_329 ();
 sg13g2_fill_1 FILLER_69_331 ();
 sg13g2_decap_8 FILLER_69_349 ();
 sg13g2_fill_1 FILLER_69_356 ();
 sg13g2_decap_8 FILLER_69_365 ();
 sg13g2_fill_1 FILLER_69_372 ();
 sg13g2_decap_8 FILLER_69_433 ();
 sg13g2_fill_2 FILLER_69_440 ();
 sg13g2_decap_8 FILLER_69_446 ();
 sg13g2_decap_8 FILLER_69_457 ();
 sg13g2_decap_4 FILLER_69_464 ();
 sg13g2_fill_2 FILLER_69_472 ();
 sg13g2_fill_1 FILLER_69_474 ();
 sg13g2_fill_2 FILLER_69_506 ();
 sg13g2_fill_1 FILLER_69_508 ();
 sg13g2_decap_8 FILLER_69_518 ();
 sg13g2_fill_2 FILLER_69_525 ();
 sg13g2_fill_2 FILLER_69_531 ();
 sg13g2_fill_2 FILLER_69_541 ();
 sg13g2_fill_1 FILLER_69_552 ();
 sg13g2_fill_2 FILLER_69_575 ();
 sg13g2_fill_2 FILLER_69_617 ();
 sg13g2_fill_1 FILLER_69_649 ();
 sg13g2_fill_2 FILLER_69_676 ();
 sg13g2_fill_1 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_683 ();
 sg13g2_fill_1 FILLER_69_711 ();
 sg13g2_fill_1 FILLER_69_726 ();
 sg13g2_fill_2 FILLER_69_732 ();
 sg13g2_fill_1 FILLER_69_752 ();
 sg13g2_decap_4 FILLER_69_779 ();
 sg13g2_fill_1 FILLER_69_783 ();
 sg13g2_fill_2 FILLER_69_801 ();
 sg13g2_fill_2 FILLER_69_820 ();
 sg13g2_fill_1 FILLER_69_822 ();
 sg13g2_fill_2 FILLER_69_832 ();
 sg13g2_fill_1 FILLER_69_834 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_4 ();
 sg13g2_fill_1 FILLER_70_48 ();
 sg13g2_fill_1 FILLER_70_67 ();
 sg13g2_decap_8 FILLER_70_85 ();
 sg13g2_fill_1 FILLER_70_92 ();
 sg13g2_fill_2 FILLER_70_98 ();
 sg13g2_fill_2 FILLER_70_117 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_fill_2 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_211 ();
 sg13g2_decap_4 FILLER_70_221 ();
 sg13g2_fill_2 FILLER_70_225 ();
 sg13g2_fill_2 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_266 ();
 sg13g2_fill_2 FILLER_70_359 ();
 sg13g2_fill_1 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_70_366 ();
 sg13g2_fill_1 FILLER_70_368 ();
 sg13g2_fill_2 FILLER_70_374 ();
 sg13g2_decap_4 FILLER_70_397 ();
 sg13g2_decap_4 FILLER_70_414 ();
 sg13g2_decap_8 FILLER_70_422 ();
 sg13g2_decap_8 FILLER_70_429 ();
 sg13g2_fill_1 FILLER_70_436 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_fill_1 FILLER_70_475 ();
 sg13g2_fill_2 FILLER_70_508 ();
 sg13g2_decap_4 FILLER_70_523 ();
 sg13g2_fill_2 FILLER_70_540 ();
 sg13g2_fill_2 FILLER_70_575 ();
 sg13g2_fill_1 FILLER_70_577 ();
 sg13g2_fill_1 FILLER_70_608 ();
 sg13g2_fill_2 FILLER_70_615 ();
 sg13g2_fill_1 FILLER_70_617 ();
 sg13g2_fill_1 FILLER_70_649 ();
 sg13g2_fill_2 FILLER_70_659 ();
 sg13g2_fill_1 FILLER_70_741 ();
 sg13g2_decap_8 FILLER_70_761 ();
 sg13g2_decap_8 FILLER_70_768 ();
 sg13g2_decap_4 FILLER_70_775 ();
 sg13g2_fill_2 FILLER_70_779 ();
 sg13g2_fill_2 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_31 ();
 sg13g2_fill_1 FILLER_71_33 ();
 sg13g2_fill_2 FILLER_71_44 ();
 sg13g2_fill_2 FILLER_71_51 ();
 sg13g2_decap_8 FILLER_71_73 ();
 sg13g2_decap_8 FILLER_71_85 ();
 sg13g2_decap_8 FILLER_71_92 ();
 sg13g2_fill_2 FILLER_71_99 ();
 sg13g2_fill_1 FILLER_71_101 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_129 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_fill_1 FILLER_71_230 ();
 sg13g2_decap_8 FILLER_71_235 ();
 sg13g2_decap_8 FILLER_71_242 ();
 sg13g2_decap_4 FILLER_71_249 ();
 sg13g2_fill_1 FILLER_71_253 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_decap_4 FILLER_71_318 ();
 sg13g2_fill_2 FILLER_71_322 ();
 sg13g2_decap_4 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_332 ();
 sg13g2_decap_8 FILLER_71_347 ();
 sg13g2_fill_2 FILLER_71_354 ();
 sg13g2_fill_1 FILLER_71_356 ();
 sg13g2_fill_2 FILLER_71_372 ();
 sg13g2_fill_1 FILLER_71_387 ();
 sg13g2_fill_2 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_398 ();
 sg13g2_decap_8 FILLER_71_405 ();
 sg13g2_fill_1 FILLER_71_412 ();
 sg13g2_fill_2 FILLER_71_446 ();
 sg13g2_decap_8 FILLER_71_503 ();
 sg13g2_fill_2 FILLER_71_510 ();
 sg13g2_fill_1 FILLER_71_512 ();
 sg13g2_decap_4 FILLER_71_544 ();
 sg13g2_fill_2 FILLER_71_574 ();
 sg13g2_fill_2 FILLER_71_585 ();
 sg13g2_fill_2 FILLER_71_596 ();
 sg13g2_fill_1 FILLER_71_598 ();
 sg13g2_fill_2 FILLER_71_612 ();
 sg13g2_fill_1 FILLER_71_614 ();
 sg13g2_fill_2 FILLER_71_678 ();
 sg13g2_fill_2 FILLER_71_699 ();
 sg13g2_decap_8 FILLER_71_735 ();
 sg13g2_decap_4 FILLER_71_742 ();
 sg13g2_fill_1 FILLER_71_746 ();
 sg13g2_fill_1 FILLER_71_778 ();
 sg13g2_decap_8 FILLER_71_783 ();
 sg13g2_decap_4 FILLER_71_790 ();
 sg13g2_fill_2 FILLER_71_794 ();
 sg13g2_fill_2 FILLER_71_833 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_50 ();
 sg13g2_fill_2 FILLER_72_66 ();
 sg13g2_fill_1 FILLER_72_72 ();
 sg13g2_fill_2 FILLER_72_89 ();
 sg13g2_fill_2 FILLER_72_104 ();
 sg13g2_fill_1 FILLER_72_119 ();
 sg13g2_fill_2 FILLER_72_173 ();
 sg13g2_fill_2 FILLER_72_203 ();
 sg13g2_fill_2 FILLER_72_209 ();
 sg13g2_fill_1 FILLER_72_239 ();
 sg13g2_fill_1 FILLER_72_253 ();
 sg13g2_decap_8 FILLER_72_328 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_388 ();
 sg13g2_fill_1 FILLER_72_416 ();
 sg13g2_fill_2 FILLER_72_450 ();
 sg13g2_fill_1 FILLER_72_452 ();
 sg13g2_decap_4 FILLER_72_468 ();
 sg13g2_decap_8 FILLER_72_526 ();
 sg13g2_fill_2 FILLER_72_533 ();
 sg13g2_fill_1 FILLER_72_535 ();
 sg13g2_decap_4 FILLER_72_541 ();
 sg13g2_fill_1 FILLER_72_572 ();
 sg13g2_fill_1 FILLER_72_596 ();
 sg13g2_fill_2 FILLER_72_623 ();
 sg13g2_fill_1 FILLER_72_625 ();
 sg13g2_fill_2 FILLER_72_655 ();
 sg13g2_decap_4 FILLER_72_684 ();
 sg13g2_fill_1 FILLER_72_702 ();
 sg13g2_fill_1 FILLER_72_718 ();
 sg13g2_decap_4 FILLER_72_746 ();
 sg13g2_fill_1 FILLER_72_754 ();
 sg13g2_fill_1 FILLER_72_773 ();
 sg13g2_fill_2 FILLER_72_859 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_2 FILLER_73_30 ();
 sg13g2_decap_4 FILLER_73_119 ();
 sg13g2_fill_2 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_184 ();
 sg13g2_fill_2 FILLER_73_198 ();
 sg13g2_decap_4 FILLER_73_221 ();
 sg13g2_decap_4 FILLER_73_235 ();
 sg13g2_fill_2 FILLER_73_239 ();
 sg13g2_fill_1 FILLER_73_267 ();
 sg13g2_decap_4 FILLER_73_349 ();
 sg13g2_fill_2 FILLER_73_353 ();
 sg13g2_decap_8 FILLER_73_377 ();
 sg13g2_fill_2 FILLER_73_384 ();
 sg13g2_decap_4 FILLER_73_390 ();
 sg13g2_fill_2 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_414 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_fill_1 FILLER_73_464 ();
 sg13g2_decap_8 FILLER_73_470 ();
 sg13g2_fill_2 FILLER_73_550 ();
 sg13g2_fill_1 FILLER_73_552 ();
 sg13g2_decap_4 FILLER_73_558 ();
 sg13g2_fill_1 FILLER_73_562 ();
 sg13g2_fill_2 FILLER_73_567 ();
 sg13g2_fill_1 FILLER_73_584 ();
 sg13g2_fill_1 FILLER_73_595 ();
 sg13g2_fill_2 FILLER_73_670 ();
 sg13g2_fill_2 FILLER_73_729 ();
 sg13g2_fill_1 FILLER_73_731 ();
 sg13g2_fill_2 FILLER_73_741 ();
 sg13g2_fill_1 FILLER_73_743 ();
 sg13g2_fill_2 FILLER_73_771 ();
 sg13g2_fill_1 FILLER_73_773 ();
 sg13g2_fill_2 FILLER_73_823 ();
 sg13g2_fill_1 FILLER_73_848 ();
 sg13g2_fill_1 FILLER_74_22 ();
 sg13g2_fill_1 FILLER_74_47 ();
 sg13g2_fill_2 FILLER_74_62 ();
 sg13g2_fill_2 FILLER_74_100 ();
 sg13g2_fill_2 FILLER_74_151 ();
 sg13g2_fill_1 FILLER_74_162 ();
 sg13g2_fill_1 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_218 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_fill_1 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_309 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_fill_1 FILLER_74_340 ();
 sg13g2_fill_1 FILLER_74_417 ();
 sg13g2_decap_8 FILLER_74_449 ();
 sg13g2_fill_1 FILLER_74_456 ();
 sg13g2_fill_2 FILLER_74_475 ();
 sg13g2_fill_1 FILLER_74_504 ();
 sg13g2_fill_2 FILLER_74_529 ();
 sg13g2_fill_2 FILLER_74_585 ();
 sg13g2_decap_8 FILLER_74_617 ();
 sg13g2_fill_2 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_626 ();
 sg13g2_fill_2 FILLER_74_631 ();
 sg13g2_fill_1 FILLER_74_645 ();
 sg13g2_fill_2 FILLER_74_651 ();
 sg13g2_decap_8 FILLER_74_666 ();
 sg13g2_fill_2 FILLER_74_673 ();
 sg13g2_fill_2 FILLER_74_737 ();
 sg13g2_fill_1 FILLER_74_744 ();
 sg13g2_fill_2 FILLER_74_750 ();
 sg13g2_decap_4 FILLER_74_766 ();
 sg13g2_fill_1 FILLER_74_797 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_127 ();
 sg13g2_fill_2 FILLER_75_133 ();
 sg13g2_fill_2 FILLER_75_162 ();
 sg13g2_fill_1 FILLER_75_164 ();
 sg13g2_fill_2 FILLER_75_195 ();
 sg13g2_decap_4 FILLER_75_226 ();
 sg13g2_fill_1 FILLER_75_230 ();
 sg13g2_decap_8 FILLER_75_235 ();
 sg13g2_decap_8 FILLER_75_257 ();
 sg13g2_decap_4 FILLER_75_264 ();
 sg13g2_fill_2 FILLER_75_272 ();
 sg13g2_decap_4 FILLER_75_286 ();
 sg13g2_decap_8 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_319 ();
 sg13g2_decap_8 FILLER_75_326 ();
 sg13g2_decap_4 FILLER_75_333 ();
 sg13g2_fill_2 FILLER_75_337 ();
 sg13g2_fill_1 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_fill_1 FILLER_75_389 ();
 sg13g2_fill_2 FILLER_75_395 ();
 sg13g2_fill_1 FILLER_75_397 ();
 sg13g2_fill_1 FILLER_75_404 ();
 sg13g2_fill_1 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_436 ();
 sg13g2_fill_2 FILLER_75_442 ();
 sg13g2_fill_1 FILLER_75_444 ();
 sg13g2_decap_8 FILLER_75_458 ();
 sg13g2_decap_4 FILLER_75_465 ();
 sg13g2_fill_2 FILLER_75_479 ();
 sg13g2_fill_1 FILLER_75_481 ();
 sg13g2_fill_2 FILLER_75_490 ();
 sg13g2_fill_2 FILLER_75_529 ();
 sg13g2_fill_1 FILLER_75_531 ();
 sg13g2_fill_2 FILLER_75_556 ();
 sg13g2_fill_2 FILLER_75_597 ();
 sg13g2_fill_1 FILLER_75_599 ();
 sg13g2_decap_8 FILLER_75_613 ();
 sg13g2_fill_2 FILLER_75_620 ();
 sg13g2_fill_2 FILLER_75_658 ();
 sg13g2_fill_1 FILLER_75_660 ();
 sg13g2_fill_1 FILLER_75_688 ();
 sg13g2_fill_2 FILLER_75_694 ();
 sg13g2_fill_1 FILLER_75_702 ();
 sg13g2_fill_1 FILLER_75_708 ();
 sg13g2_fill_1 FILLER_75_782 ();
 sg13g2_fill_2 FILLER_75_800 ();
 sg13g2_fill_1 FILLER_75_802 ();
 sg13g2_fill_2 FILLER_75_817 ();
 sg13g2_fill_1 FILLER_75_819 ();
 sg13g2_fill_2 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_4 ();
 sg13g2_fill_2 FILLER_76_33 ();
 sg13g2_fill_2 FILLER_76_76 ();
 sg13g2_fill_1 FILLER_76_78 ();
 sg13g2_decap_8 FILLER_76_131 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_208 ();
 sg13g2_decap_4 FILLER_76_223 ();
 sg13g2_fill_1 FILLER_76_227 ();
 sg13g2_decap_8 FILLER_76_319 ();
 sg13g2_decap_4 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_382 ();
 sg13g2_fill_1 FILLER_76_384 ();
 sg13g2_fill_2 FILLER_76_413 ();
 sg13g2_fill_2 FILLER_76_454 ();
 sg13g2_decap_4 FILLER_76_477 ();
 sg13g2_fill_1 FILLER_76_481 ();
 sg13g2_decap_4 FILLER_76_486 ();
 sg13g2_fill_1 FILLER_76_490 ();
 sg13g2_fill_1 FILLER_76_498 ();
 sg13g2_fill_2 FILLER_76_504 ();
 sg13g2_fill_2 FILLER_76_533 ();
 sg13g2_fill_2 FILLER_76_562 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_fill_2 FILLER_76_647 ();
 sg13g2_fill_2 FILLER_76_664 ();
 sg13g2_decap_4 FILLER_76_670 ();
 sg13g2_fill_2 FILLER_76_711 ();
 sg13g2_fill_1 FILLER_76_713 ();
 sg13g2_fill_1 FILLER_76_732 ();
 sg13g2_fill_2 FILLER_76_738 ();
 sg13g2_decap_8 FILLER_76_758 ();
 sg13g2_decap_4 FILLER_76_765 ();
 sg13g2_fill_2 FILLER_76_769 ();
 sg13g2_fill_2 FILLER_76_798 ();
 sg13g2_fill_1 FILLER_76_800 ();
 sg13g2_fill_2 FILLER_76_819 ();
 sg13g2_fill_1 FILLER_76_821 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_50 ();
 sg13g2_fill_1 FILLER_77_65 ();
 sg13g2_fill_2 FILLER_77_101 ();
 sg13g2_fill_1 FILLER_77_134 ();
 sg13g2_decap_8 FILLER_77_144 ();
 sg13g2_fill_2 FILLER_77_218 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_fill_2 FILLER_77_279 ();
 sg13g2_fill_2 FILLER_77_294 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_348 ();
 sg13g2_fill_2 FILLER_77_358 ();
 sg13g2_fill_2 FILLER_77_415 ();
 sg13g2_fill_1 FILLER_77_417 ();
 sg13g2_fill_1 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_517 ();
 sg13g2_fill_1 FILLER_77_536 ();
 sg13g2_fill_2 FILLER_77_551 ();
 sg13g2_fill_1 FILLER_77_570 ();
 sg13g2_fill_2 FILLER_77_580 ();
 sg13g2_decap_4 FILLER_77_601 ();
 sg13g2_fill_1 FILLER_77_609 ();
 sg13g2_fill_2 FILLER_77_644 ();
 sg13g2_fill_2 FILLER_77_659 ();
 sg13g2_fill_1 FILLER_77_661 ();
 sg13g2_fill_2 FILLER_77_675 ();
 sg13g2_fill_2 FILLER_77_686 ();
 sg13g2_fill_1 FILLER_77_688 ();
 sg13g2_fill_2 FILLER_77_773 ();
 sg13g2_fill_1 FILLER_77_794 ();
 sg13g2_fill_2 FILLER_77_831 ();
 sg13g2_fill_1 FILLER_77_833 ();
 sg13g2_fill_1 FILLER_77_848 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_37 ();
 sg13g2_fill_1 FILLER_78_96 ();
 sg13g2_fill_1 FILLER_78_122 ();
 sg13g2_fill_2 FILLER_78_151 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_fill_2 FILLER_78_196 ();
 sg13g2_fill_2 FILLER_78_236 ();
 sg13g2_fill_2 FILLER_78_252 ();
 sg13g2_fill_1 FILLER_78_254 ();
 sg13g2_fill_2 FILLER_78_276 ();
 sg13g2_fill_1 FILLER_78_278 ();
 sg13g2_fill_2 FILLER_78_288 ();
 sg13g2_fill_1 FILLER_78_290 ();
 sg13g2_decap_8 FILLER_78_300 ();
 sg13g2_fill_2 FILLER_78_316 ();
 sg13g2_fill_1 FILLER_78_318 ();
 sg13g2_fill_2 FILLER_78_413 ();
 sg13g2_fill_2 FILLER_78_451 ();
 sg13g2_fill_1 FILLER_78_453 ();
 sg13g2_fill_2 FILLER_78_463 ();
 sg13g2_decap_4 FILLER_78_474 ();
 sg13g2_fill_1 FILLER_78_501 ();
 sg13g2_fill_1 FILLER_78_606 ();
 sg13g2_fill_2 FILLER_78_684 ();
 sg13g2_fill_1 FILLER_78_686 ();
 sg13g2_fill_2 FILLER_78_696 ();
 sg13g2_fill_1 FILLER_78_698 ();
 sg13g2_fill_2 FILLER_78_780 ();
 sg13g2_fill_1 FILLER_78_782 ();
 sg13g2_fill_1 FILLER_78_852 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_71 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_8 FILLER_79_139 ();
 sg13g2_decap_8 FILLER_79_146 ();
 sg13g2_decap_8 FILLER_79_153 ();
 sg13g2_decap_8 FILLER_79_160 ();
 sg13g2_fill_2 FILLER_79_167 ();
 sg13g2_fill_2 FILLER_79_205 ();
 sg13g2_decap_8 FILLER_79_211 ();
 sg13g2_fill_2 FILLER_79_218 ();
 sg13g2_fill_1 FILLER_79_220 ();
 sg13g2_decap_8 FILLER_79_276 ();
 sg13g2_fill_2 FILLER_79_342 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_fill_1 FILLER_79_425 ();
 sg13g2_decap_4 FILLER_79_439 ();
 sg13g2_fill_2 FILLER_79_555 ();
 sg13g2_fill_1 FILLER_79_602 ();
 sg13g2_fill_1 FILLER_79_626 ();
 sg13g2_fill_2 FILLER_79_640 ();
 sg13g2_fill_2 FILLER_79_691 ();
 sg13g2_fill_1 FILLER_79_834 ();
 sg13g2_fill_1 FILLER_80_52 ();
 sg13g2_fill_1 FILLER_80_90 ();
 sg13g2_fill_2 FILLER_80_105 ();
 sg13g2_fill_2 FILLER_80_125 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_199 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_fill_2 FILLER_80_216 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_fill_2 FILLER_80_241 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_decap_4 FILLER_80_291 ();
 sg13g2_fill_2 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_fill_1 FILLER_80_360 ();
 sg13g2_fill_2 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_477 ();
 sg13g2_fill_2 FILLER_80_484 ();
 sg13g2_fill_1 FILLER_80_566 ();
 sg13g2_fill_2 FILLER_80_632 ();
 sg13g2_fill_2 FILLER_80_712 ();
 sg13g2_fill_1 FILLER_80_731 ();
 sg13g2_fill_2 FILLER_80_736 ();
 sg13g2_fill_1 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_fill_2 FILLER_80_794 ();
 sg13g2_fill_1 FILLER_80_796 ();
 sg13g2_fill_1 FILLER_80_814 ();
 sg13g2_fill_1 FILLER_80_819 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[4] = net20;
 assign uo_out[5] = net21;
 assign uo_out[6] = net22;
 assign uo_out[7] = net23;
endmodule
