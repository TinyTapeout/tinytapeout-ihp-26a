module tt_um_cic_filter_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire \comb1[0] ;
 wire \comb1[10] ;
 wire \comb1[11] ;
 wire \comb1[12] ;
 wire \comb1[13] ;
 wire \comb1[14] ;
 wire \comb1[15] ;
 wire \comb1[1] ;
 wire \comb1[2] ;
 wire \comb1[3] ;
 wire \comb1[4] ;
 wire \comb1[5] ;
 wire \comb1[6] ;
 wire \comb1[7] ;
 wire \comb1[8] ;
 wire \comb1[9] ;
 wire \comb1_d[0] ;
 wire \comb1_d[10] ;
 wire \comb1_d[11] ;
 wire \comb1_d[12] ;
 wire \comb1_d[13] ;
 wire \comb1_d[14] ;
 wire \comb1_d[15] ;
 wire \comb1_d[1] ;
 wire \comb1_d[2] ;
 wire \comb1_d[3] ;
 wire \comb1_d[4] ;
 wire \comb1_d[5] ;
 wire \comb1_d[6] ;
 wire \comb1_d[7] ;
 wire \comb1_d[8] ;
 wire \comb1_d[9] ;
 wire \comb2[0] ;
 wire \comb2[10] ;
 wire \comb2[11] ;
 wire \comb2[12] ;
 wire \comb2[13] ;
 wire \comb2[14] ;
 wire \comb2[15] ;
 wire \comb2[1] ;
 wire \comb2[2] ;
 wire \comb2[3] ;
 wire \comb2[4] ;
 wire \comb2[5] ;
 wire \comb2[6] ;
 wire \comb2[7] ;
 wire \comb2[8] ;
 wire \comb2[9] ;
 wire \comb2_d[0] ;
 wire \comb2_d[10] ;
 wire \comb2_d[11] ;
 wire \comb2_d[12] ;
 wire \comb2_d[13] ;
 wire \comb2_d[14] ;
 wire \comb2_d[15] ;
 wire \comb2_d[1] ;
 wire \comb2_d[2] ;
 wire \comb2_d[3] ;
 wire \comb2_d[4] ;
 wire \comb2_d[5] ;
 wire \comb2_d[6] ;
 wire \comb2_d[7] ;
 wire \comb2_d[8] ;
 wire \comb2_d[9] ;
 wire \comb3_d[0] ;
 wire \comb3_d[10] ;
 wire \comb3_d[11] ;
 wire \comb3_d[12] ;
 wire \comb3_d[13] ;
 wire \comb3_d[14] ;
 wire \comb3_d[15] ;
 wire \comb3_d[1] ;
 wire \comb3_d[2] ;
 wire \comb3_d[3] ;
 wire \comb3_d[4] ;
 wire \comb3_d[5] ;
 wire \comb3_d[6] ;
 wire \comb3_d[7] ;
 wire \comb3_d[8] ;
 wire \comb3_d[9] ;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \int1[0] ;
 wire \int1[10] ;
 wire \int1[11] ;
 wire \int1[12] ;
 wire \int1[13] ;
 wire \int1[14] ;
 wire \int1[15] ;
 wire \int1[1] ;
 wire \int1[2] ;
 wire \int1[3] ;
 wire \int1[4] ;
 wire \int1[5] ;
 wire \int1[6] ;
 wire \int1[7] ;
 wire \int1[8] ;
 wire \int1[9] ;
 wire \int2[0] ;
 wire \int2[10] ;
 wire \int2[11] ;
 wire \int2[12] ;
 wire \int2[13] ;
 wire \int2[14] ;
 wire \int2[15] ;
 wire \int2[1] ;
 wire \int2[2] ;
 wire \int2[3] ;
 wire \int2[4] ;
 wire \int2[5] ;
 wire \int2[6] ;
 wire \int2[7] ;
 wire \int2[8] ;
 wire \int2[9] ;
 wire \int3[0] ;
 wire \int3[10] ;
 wire \int3[11] ;
 wire \int3[12] ;
 wire \int3[13] ;
 wire \int3[14] ;
 wire \int3[15] ;
 wire \int3[1] ;
 wire \int3[2] ;
 wire \int3[3] ;
 wire \int3[4] ;
 wire \int3[5] ;
 wire \int3[6] ;
 wire \int3[7] ;
 wire \int3[8] ;
 wire \int3[9] ;
 wire sample_en;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_0_clk;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;

 sg13g2_inv_1 _0566_ (.Y(_0000_),
    .A(net18));
 sg13g2_inv_1 _0567_ (.Y(_0142_),
    .A(net21));
 sg13g2_inv_1 _0568_ (.Y(_0143_),
    .A(net33));
 sg13g2_inv_1 _0569_ (.Y(_0144_),
    .A(net37));
 sg13g2_inv_1 _0570_ (.Y(_0145_),
    .A(net297));
 sg13g2_inv_1 _0571_ (.Y(_0146_),
    .A(net35));
 sg13g2_inv_1 _0572_ (.Y(_0147_),
    .A(\int3[4] ));
 sg13g2_inv_1 _0573_ (.Y(_0148_),
    .A(\int3[7] ));
 sg13g2_inv_1 _0574_ (.Y(_0149_),
    .A(\comb1_d[4] ));
 sg13g2_inv_1 _0575_ (.Y(_0150_),
    .A(\comb2[4] ));
 sg13g2_nand3_1 _0576_ (.B(net18),
    .C(net23),
    .A(\count[1] ),
    .Y(_0151_));
 sg13g2_nor2_1 _0577_ (.A(_0142_),
    .B(net24),
    .Y(_0152_));
 sg13g2_and2_1 _0578_ (.A(net19),
    .B(_0152_),
    .X(_0005_));
 sg13g2_xor2_1 _0579_ (.B(net18),
    .A(net25),
    .X(_0001_));
 sg13g2_a21o_1 _0580_ (.A2(net18),
    .A1(net25),
    .B1(net23),
    .X(_0153_));
 sg13g2_and2_1 _0581_ (.A(net24),
    .B(_0153_),
    .X(_0002_));
 sg13g2_xnor2_1 _0582_ (.Y(_0003_),
    .A(net21),
    .B(_0151_));
 sg13g2_xor2_1 _0583_ (.B(_0152_),
    .A(net19),
    .X(_0004_));
 sg13g2_nand2_1 _0584_ (.Y(_0154_),
    .A(net40),
    .B(net26));
 sg13g2_nand2_1 _0585_ (.Y(_0155_),
    .A(net302),
    .B(net260));
 sg13g2_nor2_1 _0586_ (.A(net302),
    .B(net260),
    .Y(_0156_));
 sg13g2_xor2_1 _0587_ (.B(net260),
    .A(\int2[1] ),
    .X(_0157_));
 sg13g2_xnor2_1 _0588_ (.Y(_0029_),
    .A(_0154_),
    .B(net261));
 sg13g2_and2_1 _0589_ (.A(net281),
    .B(net33),
    .X(_0158_));
 sg13g2_or2_1 _0590_ (.X(_0159_),
    .B(net33),
    .A(net281));
 sg13g2_nand2b_1 _0591_ (.Y(_0160_),
    .B(_0159_),
    .A_N(_0158_));
 sg13g2_o21ai_1 _0592_ (.B1(_0155_),
    .Y(_0161_),
    .A1(_0154_),
    .A2(_0156_));
 sg13g2_xnor2_1 _0593_ (.Y(_0030_),
    .A(_0160_),
    .B(_0161_));
 sg13g2_a21o_1 _0594_ (.A2(_0161_),
    .A1(_0159_),
    .B1(_0158_),
    .X(_0162_));
 sg13g2_xnor2_1 _0595_ (.Y(_0163_),
    .A(net285),
    .B(net46));
 sg13g2_nor2b_1 _0596_ (.A(_0163_),
    .B_N(_0162_),
    .Y(_0164_));
 sg13g2_xnor2_1 _0597_ (.Y(_0031_),
    .A(_0162_),
    .B(_0163_));
 sg13g2_a21o_2 _0598_ (.A2(net46),
    .A1(net285),
    .B1(_0164_),
    .X(_0165_));
 sg13g2_nand2_1 _0599_ (.Y(_0166_),
    .A(net268),
    .B(net284));
 sg13g2_xnor2_1 _0600_ (.Y(_0167_),
    .A(net268),
    .B(net284));
 sg13g2_nand2b_1 _0601_ (.Y(_0168_),
    .B(_0165_),
    .A_N(_0167_));
 sg13g2_xnor2_1 _0602_ (.Y(_0032_),
    .A(_0165_),
    .B(_0167_));
 sg13g2_nor2_1 _0603_ (.A(net290),
    .B(net42),
    .Y(_0169_));
 sg13g2_xnor2_1 _0604_ (.Y(_0170_),
    .A(net290),
    .B(net42));
 sg13g2_nand2_1 _0605_ (.Y(_0171_),
    .A(_0166_),
    .B(_0168_));
 sg13g2_a22oi_1 _0606_ (.Y(_0172_),
    .B1(net290),
    .B2(net42),
    .A2(net284),
    .A1(net268));
 sg13g2_xnor2_1 _0607_ (.Y(_0033_),
    .A(_0170_),
    .B(_0171_));
 sg13g2_xnor2_1 _0608_ (.Y(_0173_),
    .A(net275),
    .B(net37));
 sg13g2_a21oi_1 _0609_ (.A1(_0168_),
    .A2(_0172_),
    .Y(_0174_),
    .B1(_0169_));
 sg13g2_nor2b_1 _0610_ (.A(_0173_),
    .B_N(_0174_),
    .Y(_0175_));
 sg13g2_xnor2_1 _0611_ (.Y(_0034_),
    .A(_0173_),
    .B(_0174_));
 sg13g2_nor2_1 _0612_ (.A(\int2[7] ),
    .B(\int1[7] ),
    .Y(_0176_));
 sg13g2_xnor2_1 _0613_ (.Y(_0177_),
    .A(\int2[7] ),
    .B(net44));
 sg13g2_a21oi_1 _0614_ (.A1(net275),
    .A2(net37),
    .Y(_0178_),
    .B1(_0175_));
 sg13g2_xor2_1 _0615_ (.B(_0178_),
    .A(_0177_),
    .X(_0035_));
 sg13g2_nor4_1 _0616_ (.A(_0167_),
    .B(_0170_),
    .C(_0173_),
    .D(_0177_),
    .Y(_0179_));
 sg13g2_or4_1 _0617_ (.A(_0169_),
    .B(_0172_),
    .C(_0173_),
    .D(_0177_),
    .X(_0180_));
 sg13g2_a22oi_1 _0618_ (.Y(_0181_),
    .B1(\int2[7] ),
    .B2(\int1[7] ),
    .A2(\int1[6] ),
    .A1(\int2[6] ));
 sg13g2_o21ai_1 _0619_ (.B1(_0180_),
    .Y(_0182_),
    .A1(_0176_),
    .A2(_0181_));
 sg13g2_a21o_2 _0620_ (.A2(_0179_),
    .A1(_0165_),
    .B1(_0182_),
    .X(_0183_));
 sg13g2_nand2_1 _0621_ (.Y(_0184_),
    .A(net295),
    .B(net264));
 sg13g2_xnor2_1 _0622_ (.Y(_0185_),
    .A(net295),
    .B(net264));
 sg13g2_nor2b_1 _0623_ (.A(_0185_),
    .B_N(_0183_),
    .Y(_0186_));
 sg13g2_xnor2_1 _0624_ (.Y(_0036_),
    .A(_0183_),
    .B(_0185_));
 sg13g2_nand2_1 _0625_ (.Y(_0187_),
    .A(_0145_),
    .B(_0146_));
 sg13g2_xor2_1 _0626_ (.B(net35),
    .A(\int2[9] ),
    .X(_0188_));
 sg13g2_a21oi_1 _0627_ (.A1(\int2[8] ),
    .A2(net264),
    .Y(_0189_),
    .B1(_0186_));
 sg13g2_xnor2_1 _0628_ (.Y(_0037_),
    .A(_0188_),
    .B(net265));
 sg13g2_nand2_1 _0629_ (.Y(_0190_),
    .A(\int2[10] ),
    .B(net29));
 sg13g2_xnor2_1 _0630_ (.Y(_0191_),
    .A(net305),
    .B(net29));
 sg13g2_o21ai_1 _0631_ (.B1(_0184_),
    .Y(_0192_),
    .A1(_0145_),
    .A2(_0146_));
 sg13g2_o21ai_1 _0632_ (.B1(_0187_),
    .Y(_0193_),
    .A1(_0186_),
    .A2(_0192_));
 sg13g2_xor2_1 _0633_ (.B(_0193_),
    .A(_0191_),
    .X(_0023_));
 sg13g2_nor2_1 _0634_ (.A(\int2[11] ),
    .B(net313),
    .Y(_0194_));
 sg13g2_xor2_1 _0635_ (.B(net39),
    .A(net286),
    .X(_0195_));
 sg13g2_o21ai_1 _0636_ (.B1(_0190_),
    .Y(_0196_),
    .A1(_0191_),
    .A2(_0193_));
 sg13g2_xor2_1 _0637_ (.B(_0196_),
    .A(_0195_),
    .X(_0024_));
 sg13g2_nor2b_1 _0638_ (.A(_0191_),
    .B_N(_0195_),
    .Y(_0197_));
 sg13g2_nor2b_1 _0639_ (.A(_0185_),
    .B_N(_0197_),
    .Y(_0198_));
 sg13g2_and2_1 _0640_ (.A(_0188_),
    .B(_0198_),
    .X(_0199_));
 sg13g2_nor2_1 _0641_ (.A(_0190_),
    .B(_0194_),
    .Y(_0200_));
 sg13g2_a21oi_1 _0642_ (.A1(net286),
    .A2(net39),
    .Y(_0201_),
    .B1(_0200_));
 sg13g2_nand3_1 _0643_ (.B(_0192_),
    .C(_0197_),
    .A(_0187_),
    .Y(_0202_));
 sg13g2_nand2_1 _0644_ (.Y(_0203_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_a21o_2 _0645_ (.A2(_0199_),
    .A1(_0183_),
    .B1(_0203_),
    .X(_0204_));
 sg13g2_and2_1 _0646_ (.A(net271),
    .B(net41),
    .X(_0205_));
 sg13g2_or2_1 _0647_ (.X(_0206_),
    .B(net41),
    .A(net271));
 sg13g2_nand2b_1 _0648_ (.Y(_0207_),
    .B(_0206_),
    .A_N(_0205_));
 sg13g2_xnor2_1 _0649_ (.Y(_0025_),
    .A(_0204_),
    .B(_0207_));
 sg13g2_nand2_1 _0650_ (.Y(_0208_),
    .A(\int2[13] ),
    .B(net52));
 sg13g2_xor2_1 _0651_ (.B(net52),
    .A(net294),
    .X(_0209_));
 sg13g2_a21oi_1 _0652_ (.A1(_0204_),
    .A2(_0206_),
    .Y(_0210_),
    .B1(_0205_));
 sg13g2_xnor2_1 _0653_ (.Y(_0026_),
    .A(_0209_),
    .B(_0210_));
 sg13g2_and2_1 _0654_ (.A(\int2[14] ),
    .B(\int1[14] ),
    .X(_0211_));
 sg13g2_xor2_1 _0655_ (.B(net267),
    .A(net277),
    .X(_0212_));
 sg13g2_nor2b_1 _0656_ (.A(_0207_),
    .B_N(_0209_),
    .Y(_0213_));
 sg13g2_o21ai_1 _0657_ (.B1(_0205_),
    .Y(_0214_),
    .A1(\int2[13] ),
    .A2(net52));
 sg13g2_nand2_1 _0658_ (.Y(_0215_),
    .A(_0208_),
    .B(_0214_));
 sg13g2_a21o_1 _0659_ (.A2(_0213_),
    .A1(_0204_),
    .B1(_0215_),
    .X(_0216_));
 sg13g2_xor2_1 _0660_ (.B(_0216_),
    .A(_0212_),
    .X(_0027_));
 sg13g2_a21oi_1 _0661_ (.A1(_0212_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(_0211_));
 sg13g2_xor2_1 _0662_ (.B(net256),
    .A(net31),
    .X(_0218_));
 sg13g2_xnor2_1 _0663_ (.Y(_0028_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_xor2_1 _0664_ (.B(net26),
    .A(\int1[0] ),
    .X(_0022_));
 sg13g2_nand2_1 _0665_ (.Y(_0219_),
    .A(net28),
    .B(net26));
 sg13g2_nand2_1 _0666_ (.Y(_0220_),
    .A(\int2[1] ),
    .B(net262));
 sg13g2_nor2_1 _0667_ (.A(\int2[1] ),
    .B(net262),
    .Y(_0221_));
 sg13g2_xor2_1 _0668_ (.B(net262),
    .A(\int2[1] ),
    .X(_0222_));
 sg13g2_xnor2_1 _0669_ (.Y(_0045_),
    .A(_0219_),
    .B(net263));
 sg13g2_and2_1 _0670_ (.A(net281),
    .B(\int3[2] ),
    .X(_0223_));
 sg13g2_xor2_1 _0671_ (.B(\int3[2] ),
    .A(net281),
    .X(_0224_));
 sg13g2_o21ai_1 _0672_ (.B1(_0220_),
    .Y(_0225_),
    .A1(_0219_),
    .A2(_0221_));
 sg13g2_xor2_1 _0673_ (.B(_0225_),
    .A(net282),
    .X(_0046_));
 sg13g2_a21oi_1 _0674_ (.A1(net282),
    .A2(_0225_),
    .Y(_0226_),
    .B1(_0223_));
 sg13g2_nand2_1 _0675_ (.Y(_0227_),
    .A(net285),
    .B(net288));
 sg13g2_xnor2_1 _0676_ (.Y(_0228_),
    .A(net285),
    .B(net288));
 sg13g2_xor2_1 _0677_ (.B(_0228_),
    .A(_0226_),
    .X(_0047_));
 sg13g2_o21ai_1 _0678_ (.B1(_0227_),
    .Y(_0229_),
    .A1(_0226_),
    .A2(_0228_));
 sg13g2_xnor2_1 _0679_ (.Y(_0230_),
    .A(net268),
    .B(net312));
 sg13g2_nor2b_1 _0680_ (.A(_0230_),
    .B_N(_0229_),
    .Y(_0231_));
 sg13g2_xnor2_1 _0681_ (.Y(_0048_),
    .A(_0229_),
    .B(_0230_));
 sg13g2_nor2_1 _0682_ (.A(net290),
    .B(\int3[5] ),
    .Y(_0232_));
 sg13g2_xnor2_1 _0683_ (.Y(_0233_),
    .A(\int2[5] ),
    .B(\int3[5] ));
 sg13g2_a21oi_1 _0684_ (.A1(net268),
    .A2(\int3[4] ),
    .Y(_0234_),
    .B1(_0231_));
 sg13g2_xor2_1 _0685_ (.B(net269),
    .A(_0233_),
    .X(_0049_));
 sg13g2_and2_1 _0686_ (.A(net275),
    .B(\int3[6] ),
    .X(_0235_));
 sg13g2_xor2_1 _0687_ (.B(net303),
    .A(net275),
    .X(_0236_));
 sg13g2_nor2_1 _0688_ (.A(_0230_),
    .B(_0233_),
    .Y(_0237_));
 sg13g2_a22oi_1 _0689_ (.Y(_0238_),
    .B1(\int3[5] ),
    .B2(net290),
    .A2(\int3[4] ),
    .A1(net268));
 sg13g2_nor2_1 _0690_ (.A(_0232_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_a21o_2 _0691_ (.A2(_0237_),
    .A1(_0229_),
    .B1(_0239_),
    .X(_0240_));
 sg13g2_xor2_1 _0692_ (.B(_0240_),
    .A(_0236_),
    .X(_0050_));
 sg13g2_or2_1 _0693_ (.X(_0241_),
    .B(net291),
    .A(\int2[7] ));
 sg13g2_and2_1 _0694_ (.A(\int2[7] ),
    .B(net291),
    .X(_0242_));
 sg13g2_xor2_1 _0695_ (.B(net291),
    .A(\int2[7] ),
    .X(_0243_));
 sg13g2_a21oi_1 _0696_ (.A1(_0236_),
    .A2(_0240_),
    .Y(_0244_),
    .B1(_0235_));
 sg13g2_xnor2_1 _0697_ (.Y(_0051_),
    .A(net292),
    .B(_0244_));
 sg13g2_and2_1 _0698_ (.A(_0236_),
    .B(_0243_),
    .X(_0245_));
 sg13g2_a221oi_1 _0699_ (.B2(_0240_),
    .C1(_0242_),
    .B1(_0245_),
    .A1(_0235_),
    .Y(_0246_),
    .A2(_0241_));
 sg13g2_nand2_1 _0700_ (.Y(_0247_),
    .A(net295),
    .B(\int3[8] ));
 sg13g2_xor2_1 _0701_ (.B(net310),
    .A(net295),
    .X(_0248_));
 sg13g2_nand2b_1 _0702_ (.Y(_0249_),
    .B(_0248_),
    .A_N(_0246_));
 sg13g2_xnor2_1 _0703_ (.Y(_0052_),
    .A(_0246_),
    .B(_0248_));
 sg13g2_nor2_1 _0704_ (.A(net297),
    .B(\int3[9] ),
    .Y(_0250_));
 sg13g2_xor2_1 _0705_ (.B(\int3[9] ),
    .A(net297),
    .X(_0251_));
 sg13g2_and2_1 _0706_ (.A(_0247_),
    .B(_0249_),
    .X(_0252_));
 sg13g2_xnor2_1 _0707_ (.Y(_0053_),
    .A(net298),
    .B(_0252_));
 sg13g2_and2_1 _0708_ (.A(\int2[10] ),
    .B(\int3[10] ),
    .X(_0253_));
 sg13g2_xor2_1 _0709_ (.B(\int3[10] ),
    .A(net305),
    .X(_0254_));
 sg13g2_a22oi_1 _0710_ (.Y(_0255_),
    .B1(\int3[9] ),
    .B2(net297),
    .A2(\int3[8] ),
    .A1(net295));
 sg13g2_nor2_1 _0711_ (.A(_0250_),
    .B(_0255_),
    .Y(_0256_));
 sg13g2_a21oi_1 _0712_ (.A1(_0249_),
    .A2(_0255_),
    .Y(_0257_),
    .B1(_0250_));
 sg13g2_xor2_1 _0713_ (.B(_0257_),
    .A(net306),
    .X(_0039_));
 sg13g2_or2_1 _0714_ (.X(_0258_),
    .B(\int3[11] ),
    .A(\int2[11] ));
 sg13g2_and2_1 _0715_ (.A(\int2[11] ),
    .B(\int3[11] ),
    .X(_0259_));
 sg13g2_xor2_1 _0716_ (.B(net300),
    .A(net286),
    .X(_0260_));
 sg13g2_a21oi_1 _0717_ (.A1(_0254_),
    .A2(_0257_),
    .Y(_0261_),
    .B1(_0253_));
 sg13g2_xnor2_1 _0718_ (.Y(_0040_),
    .A(_0260_),
    .B(_0261_));
 sg13g2_and2_1 _0719_ (.A(_0254_),
    .B(_0260_),
    .X(_0262_));
 sg13g2_nand3_1 _0720_ (.B(_0251_),
    .C(_0262_),
    .A(_0248_),
    .Y(_0263_));
 sg13g2_a221oi_1 _0721_ (.B2(_0256_),
    .C1(_0259_),
    .B1(_0262_),
    .A1(_0253_),
    .Y(_0264_),
    .A2(_0258_));
 sg13g2_o21ai_1 _0722_ (.B1(_0264_),
    .Y(_0265_),
    .A1(_0246_),
    .A2(_0263_));
 sg13g2_xnor2_1 _0723_ (.Y(_0266_),
    .A(net271),
    .B(net308));
 sg13g2_nor2b_1 _0724_ (.A(_0266_),
    .B_N(_0265_),
    .Y(_0267_));
 sg13g2_xnor2_1 _0725_ (.Y(_0041_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_or2_1 _0726_ (.X(_0268_),
    .B(\int3[13] ),
    .A(\int2[13] ));
 sg13g2_xor2_1 _0727_ (.B(\int3[13] ),
    .A(\int2[13] ),
    .X(_0269_));
 sg13g2_a21oi_1 _0728_ (.A1(net271),
    .A2(\int3[12] ),
    .Y(_0270_),
    .B1(_0267_));
 sg13g2_xnor2_1 _0729_ (.Y(_0042_),
    .A(_0269_),
    .B(net272));
 sg13g2_nand2_1 _0730_ (.Y(_0271_),
    .A(\int2[14] ),
    .B(\int3[14] ));
 sg13g2_nor2_1 _0731_ (.A(\int2[14] ),
    .B(\int3[14] ),
    .Y(_0272_));
 sg13g2_xor2_1 _0732_ (.B(net279),
    .A(net277),
    .X(_0273_));
 sg13g2_nor2b_1 _0733_ (.A(_0266_),
    .B_N(_0269_),
    .Y(_0274_));
 sg13g2_and3_1 _0734_ (.X(_0275_),
    .A(net271),
    .B(\int3[12] ),
    .C(_0268_));
 sg13g2_a221oi_1 _0735_ (.B2(_0274_),
    .C1(_0275_),
    .B1(_0265_),
    .A1(\int2[13] ),
    .Y(_0276_),
    .A2(\int3[13] ));
 sg13g2_xnor2_1 _0736_ (.Y(_0043_),
    .A(_0273_),
    .B(_0276_));
 sg13g2_o21ai_1 _0737_ (.B1(_0271_),
    .Y(_0277_),
    .A1(_0272_),
    .A2(_0276_));
 sg13g2_xnor2_1 _0738_ (.Y(_0278_),
    .A(net256),
    .B(net258));
 sg13g2_xnor2_1 _0739_ (.Y(_0044_),
    .A(_0277_),
    .B(_0278_));
 sg13g2_xor2_1 _0740_ (.B(net26),
    .A(net28),
    .X(_0038_));
 sg13g2_nand3_1 _0741_ (.B(net40),
    .C(net1),
    .A(net260),
    .Y(_0279_));
 sg13g2_a21o_1 _0742_ (.A2(net1),
    .A1(net40),
    .B1(net260),
    .X(_0280_));
 sg13g2_and2_1 _0743_ (.A(_0279_),
    .B(_0280_),
    .X(_0013_));
 sg13g2_nor2_2 _0744_ (.A(_0143_),
    .B(_0279_),
    .Y(_0281_));
 sg13g2_xnor2_1 _0745_ (.Y(_0014_),
    .A(net33),
    .B(_0279_));
 sg13g2_xor2_1 _0746_ (.B(_0281_),
    .A(net46),
    .X(_0015_));
 sg13g2_nand3_1 _0747_ (.B(net284),
    .C(_0281_),
    .A(net46),
    .Y(_0282_));
 sg13g2_a21o_1 _0748_ (.A2(_0281_),
    .A1(net46),
    .B1(net284),
    .X(_0283_));
 sg13g2_and2_1 _0749_ (.A(_0282_),
    .B(_0283_),
    .X(_0016_));
 sg13g2_nand4_1 _0750_ (.B(\int1[4] ),
    .C(net42),
    .A(net274),
    .Y(_0284_),
    .D(_0281_));
 sg13g2_xnor2_1 _0751_ (.Y(_0017_),
    .A(net42),
    .B(_0282_));
 sg13g2_nor2_1 _0752_ (.A(_0144_),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_xnor2_1 _0753_ (.Y(_0018_),
    .A(net37),
    .B(_0284_));
 sg13g2_xor2_1 _0754_ (.B(_0285_),
    .A(net44),
    .X(_0019_));
 sg13g2_nand3_1 _0755_ (.B(net264),
    .C(_0285_),
    .A(net44),
    .Y(_0286_));
 sg13g2_a21o_1 _0756_ (.A2(_0285_),
    .A1(net44),
    .B1(net264),
    .X(_0287_));
 sg13g2_and2_1 _0757_ (.A(_0286_),
    .B(_0287_),
    .X(_0020_));
 sg13g2_nor2_1 _0758_ (.A(_0146_),
    .B(_0286_),
    .Y(_0288_));
 sg13g2_xnor2_1 _0759_ (.Y(_0021_),
    .A(net35),
    .B(_0286_));
 sg13g2_and2_1 _0760_ (.A(net29),
    .B(_0288_),
    .X(_0289_));
 sg13g2_xor2_1 _0761_ (.B(_0288_),
    .A(net29),
    .X(_0007_));
 sg13g2_xor2_1 _0762_ (.B(_0289_),
    .A(net39),
    .X(_0008_));
 sg13g2_and3_2 _0763_ (.X(_0290_),
    .A(net39),
    .B(net41),
    .C(_0289_));
 sg13g2_a21oi_1 _0764_ (.A1(net39),
    .A2(_0289_),
    .Y(_0291_),
    .B1(net41));
 sg13g2_nor2_1 _0765_ (.A(_0290_),
    .B(_0291_),
    .Y(_0009_));
 sg13g2_xor2_1 _0766_ (.B(_0290_),
    .A(net52),
    .X(_0010_));
 sg13g2_nand3_1 _0767_ (.B(net267),
    .C(_0290_),
    .A(net52),
    .Y(_0292_));
 sg13g2_a21o_1 _0768_ (.A2(_0290_),
    .A1(net52),
    .B1(net267),
    .X(_0293_));
 sg13g2_and2_1 _0769_ (.A(_0292_),
    .B(_0293_),
    .X(_0011_));
 sg13g2_xnor2_1 _0770_ (.Y(_0012_),
    .A(net31),
    .B(_0292_));
 sg13g2_xor2_1 _0771_ (.B(net1),
    .A(net40),
    .X(_0006_));
 sg13g2_mux2_1 _0772_ (.A0(net235),
    .A1(net28),
    .S(net109),
    .X(_0054_));
 sg13g2_mux2_1 _0773_ (.A0(net147),
    .A1(\int3[1] ),
    .S(net109),
    .X(_0055_));
 sg13g2_mux2_1 _0774_ (.A0(net204),
    .A1(\int3[2] ),
    .S(net109),
    .X(_0056_));
 sg13g2_mux2_1 _0775_ (.A0(net227),
    .A1(\int3[3] ),
    .S(net109),
    .X(_0057_));
 sg13g2_nor2_1 _0776_ (.A(net69),
    .B(net104),
    .Y(_0294_));
 sg13g2_a21oi_1 _0777_ (.A1(_0147_),
    .A2(net104),
    .Y(_0058_),
    .B1(_0294_));
 sg13g2_mux2_1 _0778_ (.A0(net176),
    .A1(\int3[5] ),
    .S(net104),
    .X(_0059_));
 sg13g2_mux2_1 _0779_ (.A0(net232),
    .A1(\int3[6] ),
    .S(net103),
    .X(_0060_));
 sg13g2_nor2_1 _0780_ (.A(net187),
    .B(net103),
    .Y(_0295_));
 sg13g2_a21oi_1 _0781_ (.A1(_0148_),
    .A2(net103),
    .Y(_0061_),
    .B1(_0295_));
 sg13g2_mux2_1 _0782_ (.A0(net225),
    .A1(\int3[8] ),
    .S(net98),
    .X(_0062_));
 sg13g2_mux2_1 _0783_ (.A0(net151),
    .A1(\int3[9] ),
    .S(net98),
    .X(_0063_));
 sg13g2_mux2_1 _0784_ (.A0(net223),
    .A1(\int3[10] ),
    .S(net94),
    .X(_0064_));
 sg13g2_mux2_1 _0785_ (.A0(net248),
    .A1(\int3[11] ),
    .S(net102),
    .X(_0065_));
 sg13g2_mux2_1 _0786_ (.A0(net241),
    .A1(\int3[12] ),
    .S(net94),
    .X(_0066_));
 sg13g2_mux2_1 _0787_ (.A0(net166),
    .A1(\int3[13] ),
    .S(net94),
    .X(_0067_));
 sg13g2_mux2_1 _0788_ (.A0(net162),
    .A1(\int3[14] ),
    .S(net94),
    .X(_0068_));
 sg13g2_mux2_1 _0789_ (.A0(net91),
    .A1(\int3[15] ),
    .S(net94),
    .X(_0069_));
 sg13g2_mux2_1 _0790_ (.A0(net208),
    .A1(\comb1[0] ),
    .S(net111),
    .X(_0070_));
 sg13g2_mux2_1 _0791_ (.A0(net222),
    .A1(net171),
    .S(net111),
    .X(_0071_));
 sg13g2_mux2_1 _0792_ (.A0(net218),
    .A1(net168),
    .S(net111),
    .X(_0072_));
 sg13g2_mux2_1 _0793_ (.A0(net251),
    .A1(net211),
    .S(net112),
    .X(_0073_));
 sg13g2_mux2_1 _0794_ (.A0(net234),
    .A1(net195),
    .S(net104),
    .X(_0074_));
 sg13g2_mux2_1 _0795_ (.A0(net82),
    .A1(net61),
    .S(net104),
    .X(_0075_));
 sg13g2_mux2_1 _0796_ (.A0(net219),
    .A1(net198),
    .S(net103),
    .X(_0076_));
 sg13g2_mux2_1 _0797_ (.A0(net65),
    .A1(\comb1[7] ),
    .S(net103),
    .X(_0077_));
 sg13g2_mux2_1 _0798_ (.A0(net200),
    .A1(\comb1[8] ),
    .S(net101),
    .X(_0078_));
 sg13g2_mux2_1 _0799_ (.A0(net93),
    .A1(\comb1[9] ),
    .S(net98),
    .X(_0079_));
 sg13g2_mux2_1 _0800_ (.A0(net202),
    .A1(net153),
    .S(net98),
    .X(_0080_));
 sg13g2_mux2_1 _0801_ (.A0(net252),
    .A1(\comb1[11] ),
    .S(net99),
    .X(_0081_));
 sg13g2_mux2_1 _0802_ (.A0(net203),
    .A1(net71),
    .S(net95),
    .X(_0082_));
 sg13g2_mux2_1 _0803_ (.A0(net149),
    .A1(\comb1[13] ),
    .S(net95),
    .X(_0083_));
 sg13g2_mux2_1 _0804_ (.A0(net181),
    .A1(net155),
    .S(net95),
    .X(_0084_));
 sg13g2_mux2_1 _0805_ (.A0(net89),
    .A1(\comb1[15] ),
    .S(net95),
    .X(_0085_));
 sg13g2_mux2_1 _0806_ (.A0(net59),
    .A1(\comb2[0] ),
    .S(net110),
    .X(_0086_));
 sg13g2_mux2_1 _0807_ (.A0(net67),
    .A1(\comb2[1] ),
    .S(net111),
    .X(_0087_));
 sg13g2_mux2_1 _0808_ (.A0(net178),
    .A1(net139),
    .S(net110),
    .X(_0088_));
 sg13g2_mux2_1 _0809_ (.A0(net250),
    .A1(net78),
    .S(net110),
    .X(_0089_));
 sg13g2_nor2_1 _0810_ (.A(net53),
    .B(net112),
    .Y(_0296_));
 sg13g2_a21oi_1 _0811_ (.A1(_0150_),
    .A2(net112),
    .Y(_0090_),
    .B1(net54));
 sg13g2_mux2_1 _0812_ (.A0(net164),
    .A1(\comb2[5] ),
    .S(net107),
    .X(_0091_));
 sg13g2_mux2_1 _0813_ (.A0(net85),
    .A1(\comb2[6] ),
    .S(net107),
    .X(_0092_));
 sg13g2_mux2_1 _0814_ (.A0(net143),
    .A1(\comb2[7] ),
    .S(net107),
    .X(_0093_));
 sg13g2_mux2_1 _0815_ (.A0(net197),
    .A1(net189),
    .S(net107),
    .X(_0094_));
 sg13g2_mux2_1 _0816_ (.A0(net74),
    .A1(\comb2[9] ),
    .S(net106),
    .X(_0095_));
 sg13g2_mux2_1 _0817_ (.A0(net182),
    .A1(net83),
    .S(net100),
    .X(_0096_));
 sg13g2_mux2_1 _0818_ (.A0(net179),
    .A1(\comb2[11] ),
    .S(net99),
    .X(_0097_));
 sg13g2_mux2_1 _0819_ (.A0(net240),
    .A1(net157),
    .S(net97),
    .X(_0098_));
 sg13g2_mux2_1 _0820_ (.A0(net160),
    .A1(\comb2[13] ),
    .S(net97),
    .X(_0099_));
 sg13g2_mux2_1 _0821_ (.A0(net210),
    .A1(net183),
    .S(net97),
    .X(_0100_));
 sg13g2_mux2_1 _0822_ (.A0(net87),
    .A1(\comb2[15] ),
    .S(net96),
    .X(_0101_));
 sg13g2_nand2b_1 _0823_ (.Y(_0297_),
    .B(\comb1_d[0] ),
    .A_N(net28));
 sg13g2_xor2_1 _0824_ (.B(net235),
    .A(net28),
    .X(_0298_));
 sg13g2_mux2_1 _0825_ (.A0(net247),
    .A1(_0298_),
    .S(net111),
    .X(_0102_));
 sg13g2_nor2_1 _0826_ (.A(net171),
    .B(net109),
    .Y(_0299_));
 sg13g2_nor2b_1 _0827_ (.A(net147),
    .B_N(\int3[1] ),
    .Y(_0300_));
 sg13g2_nand2b_1 _0828_ (.Y(_0301_),
    .B(net147),
    .A_N(\int3[1] ));
 sg13g2_nor2b_1 _0829_ (.A(_0300_),
    .B_N(_0301_),
    .Y(_0302_));
 sg13g2_xnor2_1 _0830_ (.Y(_0303_),
    .A(_0297_),
    .B(_0302_));
 sg13g2_a21oi_1 _0831_ (.A1(net109),
    .A2(_0303_),
    .Y(_0103_),
    .B1(net172));
 sg13g2_a21oi_1 _0832_ (.A1(_0297_),
    .A2(_0301_),
    .Y(_0304_),
    .B1(_0300_));
 sg13g2_nand2b_1 _0833_ (.Y(_0305_),
    .B(\int3[2] ),
    .A_N(net204));
 sg13g2_xor2_1 _0834_ (.B(\comb1_d[2] ),
    .A(\int3[2] ),
    .X(_0306_));
 sg13g2_xnor2_1 _0835_ (.Y(_0307_),
    .A(_0304_),
    .B(_0306_));
 sg13g2_nor2_1 _0836_ (.A(net168),
    .B(net113),
    .Y(_0308_));
 sg13g2_a21oi_1 _0837_ (.A1(net113),
    .A2(_0307_),
    .Y(_0104_),
    .B1(net169));
 sg13g2_nor2_1 _0838_ (.A(net211),
    .B(net109),
    .Y(_0309_));
 sg13g2_nand2b_1 _0839_ (.Y(_0310_),
    .B(\comb1_d[3] ),
    .A_N(\int3[3] ));
 sg13g2_o21ai_1 _0840_ (.B1(_0305_),
    .Y(_0311_),
    .A1(_0304_),
    .A2(_0306_));
 sg13g2_nor2b_1 _0841_ (.A(\comb1_d[3] ),
    .B_N(\int3[3] ),
    .Y(_0312_));
 sg13g2_xnor2_1 _0842_ (.Y(_0313_),
    .A(\int3[3] ),
    .B(\comb1_d[3] ));
 sg13g2_xnor2_1 _0843_ (.Y(_0314_),
    .A(_0311_),
    .B(_0313_));
 sg13g2_a21oi_1 _0844_ (.A1(net109),
    .A2(_0314_),
    .Y(_0105_),
    .B1(net212));
 sg13g2_xnor2_1 _0845_ (.Y(_0315_),
    .A(\int3[4] ),
    .B(net69));
 sg13g2_inv_1 _0846_ (.Y(_0316_),
    .A(_0315_));
 sg13g2_a21oi_2 _0847_ (.B1(_0312_),
    .Y(_0317_),
    .A2(_0311_),
    .A1(_0310_));
 sg13g2_or2_1 _0848_ (.X(_0318_),
    .B(_0317_),
    .A(_0316_));
 sg13g2_xnor2_1 _0849_ (.Y(_0319_),
    .A(_0316_),
    .B(_0317_));
 sg13g2_nor2_1 _0850_ (.A(net195),
    .B(net104),
    .Y(_0320_));
 sg13g2_a21oi_1 _0851_ (.A1(net104),
    .A2(_0319_),
    .Y(_0106_),
    .B1(_0320_));
 sg13g2_o21ai_1 _0852_ (.B1(_0318_),
    .Y(_0321_),
    .A1(_0147_),
    .A2(\comb1_d[4] ));
 sg13g2_nor2b_1 _0853_ (.A(\int3[5] ),
    .B_N(\comb1_d[5] ),
    .Y(_0322_));
 sg13g2_nor2b_1 _0854_ (.A(\comb1_d[5] ),
    .B_N(\int3[5] ),
    .Y(_0323_));
 sg13g2_nor2_1 _0855_ (.A(_0322_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_xnor2_1 _0856_ (.Y(_0325_),
    .A(_0321_),
    .B(_0324_));
 sg13g2_nor2_1 _0857_ (.A(net61),
    .B(net105),
    .Y(_0326_));
 sg13g2_a21oi_1 _0858_ (.A1(net104),
    .A2(_0325_),
    .Y(_0107_),
    .B1(_0326_));
 sg13g2_nor2_1 _0859_ (.A(net198),
    .B(net103),
    .Y(_0327_));
 sg13g2_nand2b_1 _0860_ (.Y(_0328_),
    .B(\int3[6] ),
    .A_N(net232));
 sg13g2_xor2_1 _0861_ (.B(\comb1_d[6] ),
    .A(\int3[6] ),
    .X(_0329_));
 sg13g2_a21oi_1 _0862_ (.A1(\int3[4] ),
    .A2(_0149_),
    .Y(_0330_),
    .B1(_0323_));
 sg13g2_nor2_1 _0863_ (.A(_0322_),
    .B(_0330_),
    .Y(_0331_));
 sg13g2_a21o_1 _0864_ (.A2(_0330_),
    .A1(_0318_),
    .B1(_0322_),
    .X(_0332_));
 sg13g2_xnor2_1 _0865_ (.Y(_0333_),
    .A(_0329_),
    .B(_0332_));
 sg13g2_a21oi_1 _0866_ (.A1(net103),
    .A2(_0333_),
    .Y(_0108_),
    .B1(_0327_));
 sg13g2_nand2_1 _0867_ (.Y(_0334_),
    .A(_0148_),
    .B(\comb1_d[7] ));
 sg13g2_xor2_1 _0868_ (.B(net187),
    .A(\int3[7] ),
    .X(_0335_));
 sg13g2_o21ai_1 _0869_ (.B1(_0328_),
    .Y(_0336_),
    .A1(_0329_),
    .A2(_0332_));
 sg13g2_xor2_1 _0870_ (.B(_0336_),
    .A(_0335_),
    .X(_0337_));
 sg13g2_nor2_1 _0871_ (.A(net245),
    .B(net103),
    .Y(_0338_));
 sg13g2_a21oi_1 _0872_ (.A1(net105),
    .A2(_0337_),
    .Y(_0109_),
    .B1(_0338_));
 sg13g2_nor2_1 _0873_ (.A(net236),
    .B(net101),
    .Y(_0339_));
 sg13g2_nor2_1 _0874_ (.A(_0329_),
    .B(_0335_),
    .Y(_0340_));
 sg13g2_nand3_1 _0875_ (.B(_0324_),
    .C(_0340_),
    .A(_0315_),
    .Y(_0341_));
 sg13g2_o21ai_1 _0876_ (.B1(_0328_),
    .Y(_0342_),
    .A1(_0148_),
    .A2(\comb1_d[7] ));
 sg13g2_a22oi_1 _0877_ (.Y(_0343_),
    .B1(_0342_),
    .B2(_0334_),
    .A2(_0340_),
    .A1(_0331_));
 sg13g2_o21ai_1 _0878_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0317_),
    .A2(_0341_));
 sg13g2_nor2b_1 _0879_ (.A(net225),
    .B_N(\int3[8] ),
    .Y(_0345_));
 sg13g2_xor2_1 _0880_ (.B(net225),
    .A(\int3[8] ),
    .X(_0346_));
 sg13g2_nand2b_1 _0881_ (.Y(_0347_),
    .B(_0344_),
    .A_N(_0346_));
 sg13g2_xor2_1 _0882_ (.B(_0346_),
    .A(_0344_),
    .X(_0348_));
 sg13g2_a21oi_1 _0883_ (.A1(net101),
    .A2(_0348_),
    .Y(_0110_),
    .B1(net237));
 sg13g2_nor2b_2 _0884_ (.A(\int3[9] ),
    .B_N(\comb1_d[9] ),
    .Y(_0349_));
 sg13g2_nor2b_1 _0885_ (.A(\comb1_d[9] ),
    .B_N(\int3[9] ),
    .Y(_0350_));
 sg13g2_nor2_1 _0886_ (.A(_0349_),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nor2b_1 _0887_ (.A(_0345_),
    .B_N(_0347_),
    .Y(_0352_));
 sg13g2_xnor2_1 _0888_ (.Y(_0353_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_mux2_1 _0889_ (.A0(net254),
    .A1(_0353_),
    .S(net98),
    .X(_0111_));
 sg13g2_nor2_1 _0890_ (.A(net153),
    .B(net98),
    .Y(_0354_));
 sg13g2_nor2b_1 _0891_ (.A(net223),
    .B_N(\int3[10] ),
    .Y(_0355_));
 sg13g2_nand2b_1 _0892_ (.Y(_0356_),
    .B(\int3[10] ),
    .A_N(\comb1_d[10] ));
 sg13g2_nand2b_1 _0893_ (.Y(_0357_),
    .B(net223),
    .A_N(\int3[10] ));
 sg13g2_nand2_1 _0894_ (.Y(_0358_),
    .A(_0356_),
    .B(_0357_));
 sg13g2_nor2_1 _0895_ (.A(_0345_),
    .B(_0350_),
    .Y(_0359_));
 sg13g2_nor2_1 _0896_ (.A(_0349_),
    .B(_0359_),
    .Y(_0360_));
 sg13g2_a21oi_1 _0897_ (.A1(_0347_),
    .A2(_0359_),
    .Y(_0361_),
    .B1(_0349_));
 sg13g2_xor2_1 _0898_ (.B(_0361_),
    .A(_0358_),
    .X(_0362_));
 sg13g2_a21oi_1 _0899_ (.A1(net98),
    .A2(_0362_),
    .Y(_0112_),
    .B1(_0354_));
 sg13g2_nand2b_1 _0900_ (.Y(_0363_),
    .B(\int3[11] ),
    .A_N(\comb1_d[11] ));
 sg13g2_nor2b_1 _0901_ (.A(\int3[11] ),
    .B_N(\comb1_d[11] ),
    .Y(_0364_));
 sg13g2_xnor2_1 _0902_ (.Y(_0365_),
    .A(net314),
    .B(net248));
 sg13g2_a21oi_1 _0903_ (.A1(_0357_),
    .A2(_0361_),
    .Y(_0366_),
    .B1(_0355_));
 sg13g2_xnor2_1 _0904_ (.Y(_0367_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_mux2_1 _0905_ (.A0(net255),
    .A1(_0367_),
    .S(net98),
    .X(_0113_));
 sg13g2_nor2_1 _0906_ (.A(net71),
    .B(net94),
    .Y(_0368_));
 sg13g2_nor2b_1 _0907_ (.A(_0358_),
    .B_N(_0365_),
    .Y(_0369_));
 sg13g2_inv_1 _0908_ (.Y(_0370_),
    .A(_0369_));
 sg13g2_nor4_1 _0909_ (.A(_0346_),
    .B(_0349_),
    .C(_0350_),
    .D(_0370_),
    .Y(_0371_));
 sg13g2_o21ai_1 _0910_ (.B1(_0363_),
    .Y(_0372_),
    .A1(_0356_),
    .A2(_0364_));
 sg13g2_a221oi_1 _0911_ (.B2(_0344_),
    .C1(_0372_),
    .B1(_0371_),
    .A1(_0360_),
    .Y(_0373_),
    .A2(_0369_));
 sg13g2_nor2b_1 _0912_ (.A(\comb1_d[12] ),
    .B_N(\int3[12] ),
    .Y(_0374_));
 sg13g2_xor2_1 _0913_ (.B(\comb1_d[12] ),
    .A(\int3[12] ),
    .X(_0375_));
 sg13g2_nor2_1 _0914_ (.A(_0373_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_xnor2_1 _0915_ (.Y(_0377_),
    .A(_0373_),
    .B(_0375_));
 sg13g2_a21oi_1 _0916_ (.A1(net94),
    .A2(_0377_),
    .Y(_0114_),
    .B1(net72));
 sg13g2_nor2b_1 _0917_ (.A(\comb1_d[13] ),
    .B_N(\int3[13] ),
    .Y(_0378_));
 sg13g2_nand2b_1 _0918_ (.Y(_0379_),
    .B(\comb1_d[13] ),
    .A_N(\int3[13] ));
 sg13g2_nor2b_1 _0919_ (.A(_0378_),
    .B_N(_0379_),
    .Y(_0380_));
 sg13g2_nor2_1 _0920_ (.A(_0374_),
    .B(_0376_),
    .Y(_0381_));
 sg13g2_xnor2_1 _0921_ (.Y(_0382_),
    .A(_0380_),
    .B(_0381_));
 sg13g2_mux2_1 _0922_ (.A0(net216),
    .A1(_0382_),
    .S(net94),
    .X(_0115_));
 sg13g2_nor2_1 _0923_ (.A(net155),
    .B(net95),
    .Y(_0383_));
 sg13g2_nor2b_1 _0924_ (.A(net162),
    .B_N(\int3[14] ),
    .Y(_0384_));
 sg13g2_nand2b_1 _0925_ (.Y(_0385_),
    .B(net162),
    .A_N(\int3[14] ));
 sg13g2_nor2b_1 _0926_ (.A(_0384_),
    .B_N(_0385_),
    .Y(_0386_));
 sg13g2_nand2b_1 _0927_ (.Y(_0387_),
    .B(_0380_),
    .A_N(_0375_));
 sg13g2_a21oi_1 _0928_ (.A1(_0374_),
    .A2(_0379_),
    .Y(_0388_),
    .B1(_0378_));
 sg13g2_o21ai_1 _0929_ (.B1(_0388_),
    .Y(_0389_),
    .A1(_0373_),
    .A2(_0387_));
 sg13g2_xnor2_1 _0930_ (.Y(_0390_),
    .A(_0386_),
    .B(_0389_));
 sg13g2_a21oi_1 _0931_ (.A1(net95),
    .A2(_0390_),
    .Y(_0116_),
    .B1(_0383_));
 sg13g2_a21oi_1 _0932_ (.A1(_0385_),
    .A2(_0389_),
    .Y(_0391_),
    .B1(_0384_));
 sg13g2_xor2_1 _0933_ (.B(net91),
    .A(\int3[15] ),
    .X(_0392_));
 sg13g2_xnor2_1 _0934_ (.Y(_0393_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_nor2_1 _0935_ (.A(net193),
    .B(net95),
    .Y(_0394_));
 sg13g2_a21oi_1 _0936_ (.A1(net95),
    .A2(_0393_),
    .Y(_0117_),
    .B1(_0394_));
 sg13g2_nand2b_1 _0937_ (.Y(_0395_),
    .B(\comb2_d[0] ),
    .A_N(\comb1[0] ));
 sg13g2_xor2_1 _0938_ (.B(\comb2_d[0] ),
    .A(\comb1[0] ),
    .X(_0396_));
 sg13g2_mux2_1 _0939_ (.A0(net185),
    .A1(_0396_),
    .S(net110),
    .X(_0118_));
 sg13g2_nor2_1 _0940_ (.A(net174),
    .B(net110),
    .Y(_0397_));
 sg13g2_nor2b_1 _0941_ (.A(\comb2_d[1] ),
    .B_N(\comb1[1] ),
    .Y(_0398_));
 sg13g2_xnor2_1 _0942_ (.Y(_0399_),
    .A(net171),
    .B(\comb2_d[1] ));
 sg13g2_xnor2_1 _0943_ (.Y(_0400_),
    .A(_0395_),
    .B(_0399_));
 sg13g2_a21oi_1 _0944_ (.A1(net111),
    .A2(_0400_),
    .Y(_0119_),
    .B1(_0397_));
 sg13g2_nor2_1 _0945_ (.A(net139),
    .B(net110),
    .Y(_0401_));
 sg13g2_a21o_2 _0946_ (.A2(_0399_),
    .A1(_0395_),
    .B1(_0398_),
    .X(_0402_));
 sg13g2_nor2b_1 _0947_ (.A(\comb2_d[2] ),
    .B_N(\comb1[2] ),
    .Y(_0403_));
 sg13g2_nand2b_1 _0948_ (.Y(_0404_),
    .B(\comb1[2] ),
    .A_N(\comb2_d[2] ));
 sg13g2_nand2b_1 _0949_ (.Y(_0405_),
    .B(\comb2_d[2] ),
    .A_N(\comb1[2] ));
 sg13g2_nand2_1 _0950_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_xor2_1 _0951_ (.B(_0406_),
    .A(_0402_),
    .X(_0407_));
 sg13g2_a21oi_1 _0952_ (.A1(net110),
    .A2(_0407_),
    .Y(_0120_),
    .B1(_0401_));
 sg13g2_nor2_1 _0953_ (.A(net78),
    .B(net110),
    .Y(_0408_));
 sg13g2_nand2b_1 _0954_ (.Y(_0409_),
    .B(\comb1[3] ),
    .A_N(\comb2_d[3] ));
 sg13g2_nor2b_1 _0955_ (.A(\comb1[3] ),
    .B_N(\comb2_d[3] ),
    .Y(_0410_));
 sg13g2_xor2_1 _0956_ (.B(\comb2_d[3] ),
    .A(\comb1[3] ),
    .X(_0411_));
 sg13g2_a21oi_1 _0957_ (.A1(_0402_),
    .A2(_0405_),
    .Y(_0412_),
    .B1(_0403_));
 sg13g2_xnor2_1 _0958_ (.Y(_0413_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_a21oi_1 _0959_ (.A1(net111),
    .A2(_0413_),
    .Y(_0121_),
    .B1(_0408_));
 sg13g2_nand2b_1 _0960_ (.Y(_0414_),
    .B(net195),
    .A_N(\comb2_d[4] ));
 sg13g2_xor2_1 _0961_ (.B(\comb2_d[4] ),
    .A(\comb1[4] ),
    .X(_0415_));
 sg13g2_o21ai_1 _0962_ (.B1(_0409_),
    .Y(_0416_),
    .A1(_0404_),
    .A2(_0410_));
 sg13g2_nor2_1 _0963_ (.A(_0406_),
    .B(_0411_),
    .Y(_0417_));
 sg13g2_a21oi_2 _0964_ (.B1(_0416_),
    .Y(_0418_),
    .A2(_0417_),
    .A1(_0402_));
 sg13g2_o21ai_1 _0965_ (.B1(_0409_),
    .Y(_0419_),
    .A1(_0410_),
    .A2(_0412_));
 sg13g2_xnor2_1 _0966_ (.Y(_0420_),
    .A(_0415_),
    .B(_0418_));
 sg13g2_nor2_1 _0967_ (.A(net56),
    .B(net112),
    .Y(_0421_));
 sg13g2_a21oi_1 _0968_ (.A1(net112),
    .A2(_0420_),
    .Y(_0122_),
    .B1(net57));
 sg13g2_nor2b_1 _0969_ (.A(\comb1[5] ),
    .B_N(\comb2_d[5] ),
    .Y(_0422_));
 sg13g2_nand2b_1 _0970_ (.Y(_0423_),
    .B(\comb1[5] ),
    .A_N(\comb2_d[5] ));
 sg13g2_nor2b_1 _0971_ (.A(_0422_),
    .B_N(_0423_),
    .Y(_0424_));
 sg13g2_o21ai_1 _0972_ (.B1(_0414_),
    .Y(_0425_),
    .A1(_0415_),
    .A2(_0418_));
 sg13g2_xor2_1 _0973_ (.B(_0425_),
    .A(_0424_),
    .X(_0426_));
 sg13g2_mux2_1 _0974_ (.A0(net239),
    .A1(_0426_),
    .S(net107),
    .X(_0123_));
 sg13g2_nor2_1 _0975_ (.A(net145),
    .B(net107),
    .Y(_0427_));
 sg13g2_nand2b_1 _0976_ (.Y(_0428_),
    .B(net198),
    .A_N(\comb2_d[6] ));
 sg13g2_xor2_1 _0977_ (.B(\comb2_d[6] ),
    .A(\comb1[6] ),
    .X(_0429_));
 sg13g2_o21ai_1 _0978_ (.B1(_0423_),
    .Y(_0430_),
    .A1(_0414_),
    .A2(_0422_));
 sg13g2_nor2b_1 _0979_ (.A(_0415_),
    .B_N(_0424_),
    .Y(_0431_));
 sg13g2_a21oi_1 _0980_ (.A1(_0419_),
    .A2(_0431_),
    .Y(_0432_),
    .B1(_0430_));
 sg13g2_xnor2_1 _0981_ (.Y(_0433_),
    .A(_0429_),
    .B(_0432_));
 sg13g2_a21oi_1 _0982_ (.A1(net108),
    .A2(_0433_),
    .Y(_0124_),
    .B1(_0427_));
 sg13g2_nor2b_1 _0983_ (.A(\comb1[7] ),
    .B_N(\comb2_d[7] ),
    .Y(_0434_));
 sg13g2_nand2b_1 _0984_ (.Y(_0435_),
    .B(\comb1[7] ),
    .A_N(\comb2_d[7] ));
 sg13g2_nor2b_1 _0985_ (.A(_0434_),
    .B_N(_0435_),
    .Y(_0436_));
 sg13g2_o21ai_1 _0986_ (.B1(_0428_),
    .Y(_0437_),
    .A1(_0429_),
    .A2(_0432_));
 sg13g2_xor2_1 _0987_ (.B(_0437_),
    .A(_0436_),
    .X(_0438_));
 sg13g2_mux2_1 _0988_ (.A0(net230),
    .A1(_0438_),
    .S(net108),
    .X(_0125_));
 sg13g2_nor2_1 _0989_ (.A(net189),
    .B(net106),
    .Y(_0439_));
 sg13g2_nor2b_1 _0990_ (.A(_0429_),
    .B_N(_0436_),
    .Y(_0440_));
 sg13g2_nand2_1 _0991_ (.Y(_0441_),
    .A(_0431_),
    .B(_0440_));
 sg13g2_o21ai_1 _0992_ (.B1(_0435_),
    .Y(_0442_),
    .A1(_0428_),
    .A2(_0434_));
 sg13g2_a21oi_1 _0993_ (.A1(_0430_),
    .A2(_0440_),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_o21ai_1 _0994_ (.B1(_0443_),
    .Y(_0444_),
    .A1(_0418_),
    .A2(_0441_));
 sg13g2_nand2b_1 _0995_ (.Y(_0445_),
    .B(\comb1[8] ),
    .A_N(\comb2_d[8] ));
 sg13g2_xor2_1 _0996_ (.B(\comb2_d[8] ),
    .A(\comb1[8] ),
    .X(_0446_));
 sg13g2_nand2b_1 _0997_ (.Y(_0447_),
    .B(_0444_),
    .A_N(_0446_));
 sg13g2_xor2_1 _0998_ (.B(_0446_),
    .A(_0444_),
    .X(_0448_));
 sg13g2_a21oi_1 _0999_ (.A1(net106),
    .A2(_0448_),
    .Y(_0126_),
    .B1(_0439_));
 sg13g2_nor2b_1 _1000_ (.A(\comb1[9] ),
    .B_N(\comb2_d[9] ),
    .Y(_0449_));
 sg13g2_nand2b_1 _1001_ (.Y(_0450_),
    .B(\comb1[9] ),
    .A_N(\comb2_d[9] ));
 sg13g2_nor2b_1 _1002_ (.A(_0449_),
    .B_N(_0450_),
    .Y(_0451_));
 sg13g2_nand2_1 _1003_ (.Y(_0452_),
    .A(_0445_),
    .B(_0447_));
 sg13g2_xor2_1 _1004_ (.B(_0452_),
    .A(_0451_),
    .X(_0453_));
 sg13g2_mux2_1 _1005_ (.A0(net206),
    .A1(_0453_),
    .S(net100),
    .X(_0127_));
 sg13g2_nor2_1 _1006_ (.A(net83),
    .B(net99),
    .Y(_0454_));
 sg13g2_nand2b_1 _1007_ (.Y(_0455_),
    .B(net153),
    .A_N(\comb2_d[10] ));
 sg13g2_xor2_1 _1008_ (.B(\comb2_d[10] ),
    .A(\comb1[10] ),
    .X(_0456_));
 sg13g2_o21ai_1 _1009_ (.B1(_0450_),
    .Y(_0457_),
    .A1(_0445_),
    .A2(_0449_));
 sg13g2_nor2b_1 _1010_ (.A(_0446_),
    .B_N(_0451_),
    .Y(_0458_));
 sg13g2_a21oi_1 _1011_ (.A1(_0444_),
    .A2(_0458_),
    .Y(_0459_),
    .B1(_0457_));
 sg13g2_xnor2_1 _1012_ (.Y(_0460_),
    .A(_0456_),
    .B(_0459_));
 sg13g2_a21oi_1 _1013_ (.A1(net99),
    .A2(_0460_),
    .Y(_0128_),
    .B1(_0454_));
 sg13g2_nand2b_1 _1014_ (.Y(_0461_),
    .B(\comb1[11] ),
    .A_N(\comb2_d[11] ));
 sg13g2_nor2b_1 _1015_ (.A(\comb1[11] ),
    .B_N(\comb2_d[11] ),
    .Y(_0462_));
 sg13g2_xnor2_1 _1016_ (.Y(_0463_),
    .A(\comb1[11] ),
    .B(\comb2_d[11] ));
 sg13g2_o21ai_1 _1017_ (.B1(_0455_),
    .Y(_0464_),
    .A1(_0456_),
    .A2(_0459_));
 sg13g2_xor2_1 _1018_ (.B(_0464_),
    .A(_0463_),
    .X(_0465_));
 sg13g2_mux2_1 _1019_ (.A0(net243),
    .A1(_0465_),
    .S(net99),
    .X(_0129_));
 sg13g2_nor2_1 _1020_ (.A(net157),
    .B(net97),
    .Y(_0466_));
 sg13g2_nor2b_1 _1021_ (.A(_0456_),
    .B_N(_0463_),
    .Y(_0467_));
 sg13g2_and2_1 _1022_ (.A(_0458_),
    .B(_0467_),
    .X(_0468_));
 sg13g2_o21ai_1 _1023_ (.B1(_0461_),
    .Y(_0469_),
    .A1(_0455_),
    .A2(_0462_));
 sg13g2_a221oi_1 _1024_ (.B2(_0444_),
    .C1(_0469_),
    .B1(_0468_),
    .A1(_0457_),
    .Y(_0470_),
    .A2(_0467_));
 sg13g2_nor2b_1 _1025_ (.A(net203),
    .B_N(\comb1[12] ),
    .Y(_0471_));
 sg13g2_xor2_1 _1026_ (.B(\comb2_d[12] ),
    .A(net71),
    .X(_0472_));
 sg13g2_nor2_1 _1027_ (.A(_0470_),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_xnor2_1 _1028_ (.Y(_0474_),
    .A(_0470_),
    .B(_0472_));
 sg13g2_a21oi_1 _1029_ (.A1(net97),
    .A2(_0474_),
    .Y(_0130_),
    .B1(net158));
 sg13g2_nor2b_1 _1030_ (.A(net149),
    .B_N(\comb1[13] ),
    .Y(_0475_));
 sg13g2_nand2b_1 _1031_ (.Y(_0476_),
    .B(\comb2_d[13] ),
    .A_N(\comb1[13] ));
 sg13g2_nor2b_1 _1032_ (.A(_0475_),
    .B_N(_0476_),
    .Y(_0477_));
 sg13g2_nor2_1 _1033_ (.A(_0471_),
    .B(_0473_),
    .Y(_0478_));
 sg13g2_xnor2_1 _1034_ (.Y(_0479_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_mux2_1 _1035_ (.A0(net220),
    .A1(_0479_),
    .S(net97),
    .X(_0131_));
 sg13g2_nor2_1 _1036_ (.A(net183),
    .B(net96),
    .Y(_0480_));
 sg13g2_nor2b_1 _1037_ (.A(net181),
    .B_N(\comb1[14] ),
    .Y(_0481_));
 sg13g2_nand2b_1 _1038_ (.Y(_0482_),
    .B(net181),
    .A_N(\comb1[14] ));
 sg13g2_nor2b_1 _1039_ (.A(_0481_),
    .B_N(_0482_),
    .Y(_0483_));
 sg13g2_nand2b_1 _1040_ (.Y(_0484_),
    .B(_0477_),
    .A_N(_0472_));
 sg13g2_a21oi_1 _1041_ (.A1(_0471_),
    .A2(_0476_),
    .Y(_0485_),
    .B1(_0475_));
 sg13g2_o21ai_1 _1042_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0470_),
    .A2(_0484_));
 sg13g2_xnor2_1 _1043_ (.Y(_0487_),
    .A(_0483_),
    .B(_0486_));
 sg13g2_a21oi_1 _1044_ (.A1(net96),
    .A2(_0487_),
    .Y(_0132_),
    .B1(_0480_));
 sg13g2_a21oi_1 _1045_ (.A1(_0482_),
    .A2(_0486_),
    .Y(_0488_),
    .B1(_0481_));
 sg13g2_xor2_1 _1046_ (.B(net89),
    .A(\comb1[15] ),
    .X(_0489_));
 sg13g2_xnor2_1 _1047_ (.Y(_0490_),
    .A(_0488_),
    .B(_0489_));
 sg13g2_nor2_1 _1048_ (.A(net141),
    .B(net96),
    .Y(_0491_));
 sg13g2_a21oi_1 _1049_ (.A1(net96),
    .A2(_0490_),
    .Y(_0133_),
    .B1(_0491_));
 sg13g2_nor2_1 _1050_ (.A(net106),
    .B(net76),
    .Y(_0492_));
 sg13g2_nor2b_1 _1051_ (.A(\comb3_d[2] ),
    .B_N(\comb2[2] ),
    .Y(_0493_));
 sg13g2_nor2b_1 _1052_ (.A(\comb3_d[3] ),
    .B_N(\comb2[3] ),
    .Y(_0494_));
 sg13g2_or2_1 _1053_ (.X(_0495_),
    .B(_0494_),
    .A(_0493_));
 sg13g2_nor2b_1 _1054_ (.A(\comb2[3] ),
    .B_N(\comb3_d[3] ),
    .Y(_0496_));
 sg13g2_nand2b_1 _1055_ (.Y(_0497_),
    .B(\comb3_d[3] ),
    .A_N(\comb2[3] ));
 sg13g2_nand2b_1 _1056_ (.Y(_0498_),
    .B(\comb2[1] ),
    .A_N(\comb3_d[1] ));
 sg13g2_nor2b_1 _1057_ (.A(\comb2[0] ),
    .B_N(\comb3_d[0] ),
    .Y(_0499_));
 sg13g2_nor2b_1 _1058_ (.A(\comb2[1] ),
    .B_N(\comb3_d[1] ),
    .Y(_0500_));
 sg13g2_o21ai_1 _1059_ (.B1(_0498_),
    .Y(_0501_),
    .A1(_0499_),
    .A2(_0500_));
 sg13g2_nor2b_1 _1060_ (.A(\comb2[2] ),
    .B_N(\comb3_d[2] ),
    .Y(_0502_));
 sg13g2_nor4_1 _1061_ (.A(_0493_),
    .B(_0494_),
    .C(_0496_),
    .D(_0502_),
    .Y(_0503_));
 sg13g2_a22oi_1 _1062_ (.Y(_0504_),
    .B1(_0501_),
    .B2(_0503_),
    .A2(_0497_),
    .A1(_0495_));
 sg13g2_nand2b_1 _1063_ (.Y(_0505_),
    .B(\comb2[6] ),
    .A_N(\comb3_d[6] ));
 sg13g2_nand2b_1 _1064_ (.Y(_0506_),
    .B(\comb2[7] ),
    .A_N(\comb3_d[7] ));
 sg13g2_nand2_1 _1065_ (.Y(_0507_),
    .A(_0505_),
    .B(_0506_));
 sg13g2_nand2b_1 _1066_ (.Y(_0508_),
    .B(\comb3_d[6] ),
    .A_N(\comb2[6] ));
 sg13g2_nand2b_1 _1067_ (.Y(_0509_),
    .B(\comb3_d[7] ),
    .A_N(\comb2[7] ));
 sg13g2_and4_1 _1068_ (.A(_0505_),
    .B(_0506_),
    .C(_0508_),
    .D(_0509_),
    .X(_0510_));
 sg13g2_nand2b_1 _1069_ (.Y(_0511_),
    .B(\comb2[4] ),
    .A_N(\comb3_d[4] ));
 sg13g2_nand2b_1 _1070_ (.Y(_0512_),
    .B(\comb2[5] ),
    .A_N(\comb3_d[5] ));
 sg13g2_nor2b_1 _1071_ (.A(\comb2[5] ),
    .B_N(\comb3_d[5] ),
    .Y(_0513_));
 sg13g2_a21oi_1 _1072_ (.A1(_0150_),
    .A2(\comb3_d[4] ),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_nand4_1 _1073_ (.B(_0511_),
    .C(_0512_),
    .A(_0510_),
    .Y(_0515_),
    .D(_0514_));
 sg13g2_nor2_1 _1074_ (.A(_0504_),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_a21oi_1 _1075_ (.A1(_0511_),
    .A2(_0512_),
    .Y(_0517_),
    .B1(_0513_));
 sg13g2_a22oi_1 _1076_ (.Y(_0518_),
    .B1(_0510_),
    .B2(_0517_),
    .A2(_0509_),
    .A1(_0507_));
 sg13g2_nor2b_1 _1077_ (.A(_0516_),
    .B_N(_0518_),
    .Y(_0519_));
 sg13g2_o21ai_1 _1078_ (.B1(_0518_),
    .Y(_0520_),
    .A1(_0504_),
    .A2(_0515_));
 sg13g2_nand2b_1 _1079_ (.Y(_0521_),
    .B(net189),
    .A_N(\comb3_d[8] ));
 sg13g2_xor2_1 _1080_ (.B(\comb3_d[8] ),
    .A(\comb2[8] ),
    .X(_0522_));
 sg13g2_xor2_1 _1081_ (.B(_0522_),
    .A(_0520_),
    .X(_0523_));
 sg13g2_a21oi_1 _1082_ (.A1(net106),
    .A2(_0523_),
    .Y(_0134_),
    .B1(_0492_));
 sg13g2_nor2b_1 _1083_ (.A(\comb2[9] ),
    .B_N(\comb3_d[9] ),
    .Y(_0524_));
 sg13g2_nand2b_1 _1084_ (.Y(_0525_),
    .B(\comb2[9] ),
    .A_N(\comb3_d[9] ));
 sg13g2_nor2b_1 _1085_ (.A(_0524_),
    .B_N(_0525_),
    .Y(_0526_));
 sg13g2_o21ai_1 _1086_ (.B1(_0521_),
    .Y(_0527_),
    .A1(_0519_),
    .A2(_0522_));
 sg13g2_xor2_1 _1087_ (.B(_0527_),
    .A(_0526_),
    .X(_0528_));
 sg13g2_mux2_1 _1088_ (.A0(net229),
    .A1(_0528_),
    .S(net107),
    .X(_0135_));
 sg13g2_nor2_1 _1089_ (.A(net106),
    .B(net48),
    .Y(_0529_));
 sg13g2_nor2b_1 _1090_ (.A(\comb3_d[10] ),
    .B_N(\comb2[10] ),
    .Y(_0530_));
 sg13g2_inv_1 _1091_ (.Y(_0531_),
    .A(_0530_));
 sg13g2_nand2b_1 _1092_ (.Y(_0532_),
    .B(\comb3_d[10] ),
    .A_N(\comb2[10] ));
 sg13g2_nand2_1 _1093_ (.Y(_0533_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_nor2b_1 _1094_ (.A(_0522_),
    .B_N(_0526_),
    .Y(_0534_));
 sg13g2_o21ai_1 _1095_ (.B1(_0525_),
    .Y(_0535_),
    .A1(_0521_),
    .A2(_0524_));
 sg13g2_a21oi_2 _1096_ (.B1(_0535_),
    .Y(_0536_),
    .A2(_0534_),
    .A1(_0520_));
 sg13g2_xnor2_1 _1097_ (.Y(_0537_),
    .A(_0533_),
    .B(_0536_));
 sg13g2_a21oi_1 _1098_ (.A1(net106),
    .A2(_0537_),
    .Y(_0136_),
    .B1(_0529_));
 sg13g2_nor2_1 _1099_ (.A(net106),
    .B(net50),
    .Y(_0538_));
 sg13g2_nor2b_1 _1100_ (.A(\comb3_d[11] ),
    .B_N(\comb2[11] ),
    .Y(_0539_));
 sg13g2_nand2b_1 _1101_ (.Y(_0540_),
    .B(\comb3_d[11] ),
    .A_N(\comb2[11] ));
 sg13g2_nor2b_1 _1102_ (.A(_0539_),
    .B_N(_0540_),
    .Y(_0541_));
 sg13g2_o21ai_1 _1103_ (.B1(_0531_),
    .Y(_0542_),
    .A1(_0533_),
    .A2(_0536_));
 sg13g2_xnor2_1 _1104_ (.Y(_0543_),
    .A(_0541_),
    .B(_0542_));
 sg13g2_a21oi_1 _1105_ (.A1(net100),
    .A2(_0543_),
    .Y(_0137_),
    .B1(_0538_));
 sg13g2_nor2_1 _1106_ (.A(net100),
    .B(net63),
    .Y(_0544_));
 sg13g2_a21oi_1 _1107_ (.A1(_0530_),
    .A2(_0540_),
    .Y(_0545_),
    .B1(_0539_));
 sg13g2_o21ai_1 _1108_ (.B1(_0540_),
    .Y(_0546_),
    .A1(_0532_),
    .A2(_0539_));
 sg13g2_a21oi_2 _1109_ (.B1(_0546_),
    .Y(_0547_),
    .A2(_0545_),
    .A1(_0536_));
 sg13g2_nor2b_1 _1110_ (.A(\comb3_d[12] ),
    .B_N(\comb2[12] ),
    .Y(_0548_));
 sg13g2_xnor2_1 _1111_ (.Y(_0549_),
    .A(\comb2[12] ),
    .B(\comb3_d[12] ));
 sg13g2_xnor2_1 _1112_ (.Y(_0550_),
    .A(_0547_),
    .B(_0549_));
 sg13g2_a21oi_1 _1113_ (.A1(net100),
    .A2(_0550_),
    .Y(_0138_),
    .B1(_0544_));
 sg13g2_nor2b_1 _1114_ (.A(\comb3_d[13] ),
    .B_N(\comb2[13] ),
    .Y(_0551_));
 sg13g2_nand2b_1 _1115_ (.Y(_0552_),
    .B(\comb3_d[13] ),
    .A_N(\comb2[13] ));
 sg13g2_nor2b_1 _1116_ (.A(_0551_),
    .B_N(_0552_),
    .Y(_0553_));
 sg13g2_a21oi_1 _1117_ (.A1(_0547_),
    .A2(_0549_),
    .Y(_0554_),
    .B1(_0548_));
 sg13g2_xnor2_1 _1118_ (.Y(_0555_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_mux2_1 _1119_ (.A0(net214),
    .A1(_0555_),
    .S(net100),
    .X(_0139_));
 sg13g2_nor2_1 _1120_ (.A(net100),
    .B(net80),
    .Y(_0556_));
 sg13g2_nand2b_1 _1121_ (.Y(_0557_),
    .B(net183),
    .A_N(\comb3_d[14] ));
 sg13g2_xor2_1 _1122_ (.B(\comb3_d[14] ),
    .A(\comb2[14] ),
    .X(_0558_));
 sg13g2_and2_1 _1123_ (.A(_0549_),
    .B(_0553_),
    .X(_0559_));
 sg13g2_a221oi_1 _1124_ (.B2(_0547_),
    .C1(_0551_),
    .B1(_0559_),
    .A1(_0548_),
    .Y(_0560_),
    .A2(_0552_));
 sg13g2_xnor2_1 _1125_ (.Y(_0561_),
    .A(_0558_),
    .B(_0560_));
 sg13g2_a21oi_1 _1126_ (.A1(net99),
    .A2(_0561_),
    .Y(_0140_),
    .B1(_0556_));
 sg13g2_o21ai_1 _1127_ (.B1(_0557_),
    .Y(_0562_),
    .A1(_0558_),
    .A2(_0560_));
 sg13g2_xnor2_1 _1128_ (.Y(_0563_),
    .A(net141),
    .B(net87));
 sg13g2_nor2_1 _1129_ (.A(net99),
    .B(net191),
    .Y(_0564_));
 sg13g2_xnor2_1 _1130_ (.Y(_0565_),
    .A(_0562_),
    .B(_0563_));
 sg13g2_a21oi_1 _1131_ (.A1(net99),
    .A2(_0565_),
    .Y(_0141_),
    .B1(_0564_));
 sg13g2_dfrbpq_1 _1132_ (.RESET_B(net135),
    .D(_0054_),
    .Q(\comb1_d[0] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1133_ (.RESET_B(net129),
    .D(net148),
    .Q(\comb1_d[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1134_ (.RESET_B(net129),
    .D(net205),
    .Q(\comb1_d[2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1135_ (.RESET_B(net129),
    .D(net228),
    .Q(\comb1_d[3] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1136_ (.RESET_B(net127),
    .D(net70),
    .Q(\comb1_d[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1137_ (.RESET_B(net125),
    .D(net177),
    .Q(\comb1_d[5] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1138_ (.RESET_B(net137),
    .D(net233),
    .Q(\comb1_d[6] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1139_ (.RESET_B(net127),
    .D(net188),
    .Q(\comb1_d[7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1140_ (.RESET_B(net119),
    .D(net226),
    .Q(\comb1_d[8] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1141_ (.RESET_B(net119),
    .D(net152),
    .Q(\comb1_d[9] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1142_ (.RESET_B(net119),
    .D(net224),
    .Q(\comb1_d[10] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1143_ (.RESET_B(net117),
    .D(net249),
    .Q(\comb1_d[11] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1144_ (.RESET_B(net116),
    .D(net242),
    .Q(\comb1_d[12] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1145_ (.RESET_B(net116),
    .D(net167),
    .Q(\comb1_d[13] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1146_ (.RESET_B(net116),
    .D(net163),
    .Q(\comb1_d[14] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1147_ (.RESET_B(net116),
    .D(net92),
    .Q(\comb1_d[15] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1148_ (.RESET_B(net133),
    .D(net209),
    .Q(\comb2_d[0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1149_ (.RESET_B(net135),
    .D(_0071_),
    .Q(\comb2_d[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1150_ (.RESET_B(net135),
    .D(_0072_),
    .Q(\comb2_d[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1151_ (.RESET_B(net135),
    .D(_0073_),
    .Q(\comb2_d[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1152_ (.RESET_B(net132),
    .D(_0074_),
    .Q(\comb2_d[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1153_ (.RESET_B(net132),
    .D(_0075_),
    .Q(\comb2_d[5] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1154_ (.RESET_B(net132),
    .D(_0076_),
    .Q(\comb2_d[6] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1155_ (.RESET_B(net132),
    .D(net66),
    .Q(\comb2_d[7] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1156_ (.RESET_B(net123),
    .D(net201),
    .Q(\comb2_d[8] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1157_ (.RESET_B(net123),
    .D(net138),
    .Q(\comb2_d[9] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1158_ (.RESET_B(net123),
    .D(_0080_),
    .Q(\comb2_d[10] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1159_ (.RESET_B(net123),
    .D(net253),
    .Q(\comb2_d[11] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1160_ (.RESET_B(net121),
    .D(_0082_),
    .Q(\comb2_d[12] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1161_ (.RESET_B(net121),
    .D(net150),
    .Q(\comb2_d[13] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1162_ (.RESET_B(net120),
    .D(_0084_),
    .Q(\comb2_d[14] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1163_ (.RESET_B(net120),
    .D(net90),
    .Q(\comb2_d[15] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1164_ (.RESET_B(net133),
    .D(net60),
    .Q(\comb3_d[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1165_ (.RESET_B(net133),
    .D(net68),
    .Q(\comb3_d[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1166_ (.RESET_B(net133),
    .D(_0088_),
    .Q(\comb3_d[2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1167_ (.RESET_B(net134),
    .D(_0089_),
    .Q(\comb3_d[3] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1168_ (.RESET_B(net132),
    .D(net55),
    .Q(\comb3_d[4] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1169_ (.RESET_B(net134),
    .D(net165),
    .Q(\comb3_d[5] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1170_ (.RESET_B(net131),
    .D(net86),
    .Q(\comb3_d[6] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1171_ (.RESET_B(net136),
    .D(net144),
    .Q(\comb3_d[7] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1172_ (.RESET_B(net131),
    .D(_0094_),
    .Q(\comb3_d[8] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1173_ (.RESET_B(net131),
    .D(net75),
    .Q(\comb3_d[9] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1174_ (.RESET_B(net122),
    .D(_0096_),
    .Q(\comb3_d[10] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1175_ (.RESET_B(net122),
    .D(net180),
    .Q(\comb3_d[11] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1176_ (.RESET_B(net120),
    .D(_0098_),
    .Q(\comb3_d[12] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1177_ (.RESET_B(net120),
    .D(net161),
    .Q(\comb3_d[13] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1178_ (.RESET_B(net121),
    .D(_0100_),
    .Q(\comb3_d[14] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1179_ (.RESET_B(net120),
    .D(net88),
    .Q(\comb3_d[15] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1180_ (.RESET_B(net135),
    .D(_0102_),
    .Q(\comb1[0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1181_ (.RESET_B(net135),
    .D(net173),
    .Q(\comb1[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1182_ (.RESET_B(net135),
    .D(net170),
    .Q(\comb1[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1183_ (.RESET_B(net135),
    .D(net213),
    .Q(\comb1[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1184_ (.RESET_B(net127),
    .D(net196),
    .Q(\comb1[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1185_ (.RESET_B(net127),
    .D(net62),
    .Q(\comb1[5] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1186_ (.RESET_B(net127),
    .D(net199),
    .Q(\comb1[6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1187_ (.RESET_B(net127),
    .D(net246),
    .Q(\comb1[7] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1188_ (.RESET_B(net123),
    .D(net238),
    .Q(\comb1[8] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1189_ (.RESET_B(net123),
    .D(_0111_),
    .Q(\comb1[9] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1190_ (.RESET_B(net123),
    .D(net154),
    .Q(\comb1[10] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1191_ (.RESET_B(net123),
    .D(_0113_),
    .Q(\comb1[11] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1192_ (.RESET_B(net121),
    .D(net73),
    .Q(\comb1[12] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1193_ (.RESET_B(net121),
    .D(net217),
    .Q(\comb1[13] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1194_ (.RESET_B(net121),
    .D(net156),
    .Q(\comb1[14] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1195_ (.RESET_B(net121),
    .D(net194),
    .Q(\comb1[15] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1196_ (.RESET_B(net133),
    .D(net186),
    .Q(\comb2[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1197_ (.RESET_B(net133),
    .D(net175),
    .Q(\comb2[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1198_ (.RESET_B(net133),
    .D(net140),
    .Q(\comb2[2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1199_ (.RESET_B(net133),
    .D(net79),
    .Q(\comb2[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1200_ (.RESET_B(net136),
    .D(net58),
    .Q(\comb2[4] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1201_ (.RESET_B(net134),
    .D(_0123_),
    .Q(\comb2[5] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1202_ (.RESET_B(net132),
    .D(net146),
    .Q(\comb2[6] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1203_ (.RESET_B(net132),
    .D(net231),
    .Q(\comb2[7] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1204_ (.RESET_B(net131),
    .D(net190),
    .Q(\comb2[8] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1205_ (.RESET_B(net131),
    .D(net207),
    .Q(\comb2[9] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1206_ (.RESET_B(net122),
    .D(net84),
    .Q(\comb2[10] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1207_ (.RESET_B(net122),
    .D(net244),
    .Q(\comb2[11] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1208_ (.RESET_B(net120),
    .D(net159),
    .Q(\comb2[12] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1209_ (.RESET_B(net124),
    .D(net221),
    .Q(\comb2[13] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1210_ (.RESET_B(net120),
    .D(net184),
    .Q(\comb2[14] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1211_ (.RESET_B(net120),
    .D(net142),
    .Q(\comb2[15] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1212_ (.RESET_B(net128),
    .D(_0000_),
    .Q(\count[0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1213_ (.RESET_B(net128),
    .D(_0001_),
    .Q(\count[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1214_ (.RESET_B(net128),
    .D(_0002_),
    .Q(\count[2] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1215_ (.RESET_B(net130),
    .D(net22),
    .Q(\count[3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1216_ (.RESET_B(net130),
    .D(net20),
    .Q(\count[4] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1217_ (.RESET_B(net128),
    .D(_0005_),
    .Q(sample_en),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1218_ (.RESET_B(net129),
    .D(_0006_),
    .Q(\int1[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1219_ (.RESET_B(net130),
    .D(_0013_),
    .Q(\int1[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1220_ (.RESET_B(net128),
    .D(net34),
    .Q(\int1[2] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1221_ (.RESET_B(net125),
    .D(net47),
    .Q(\int1[3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1222_ (.RESET_B(net125),
    .D(_0016_),
    .Q(\int1[4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1223_ (.RESET_B(net126),
    .D(net43),
    .Q(\int1[5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1224_ (.RESET_B(net125),
    .D(net38),
    .Q(\int1[6] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1225_ (.RESET_B(net118),
    .D(net45),
    .Q(\int1[7] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1226_ (.RESET_B(net118),
    .D(_0020_),
    .Q(\int1[8] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1227_ (.RESET_B(net118),
    .D(net36),
    .Q(\int1[9] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1228_ (.RESET_B(net115),
    .D(net30),
    .Q(\int1[10] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1229_ (.RESET_B(net115),
    .D(_0008_),
    .Q(\int1[11] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1230_ (.RESET_B(net114),
    .D(_0009_),
    .Q(\int1[12] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1231_ (.RESET_B(net114),
    .D(_0010_),
    .Q(\int1[13] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1232_ (.RESET_B(net114),
    .D(_0011_),
    .Q(\int1[14] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1233_ (.RESET_B(net114),
    .D(net32),
    .Q(\int1[15] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1234_ (.RESET_B(net129),
    .D(net27),
    .Q(\int2[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1235_ (.RESET_B(net129),
    .D(_0029_),
    .Q(\int2[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1236_ (.RESET_B(net128),
    .D(_0030_),
    .Q(\int2[2] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1237_ (.RESET_B(net128),
    .D(_0031_),
    .Q(\int2[3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1238_ (.RESET_B(net126),
    .D(_0032_),
    .Q(\int2[4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1239_ (.RESET_B(net126),
    .D(_0033_),
    .Q(\int2[5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1240_ (.RESET_B(net125),
    .D(_0034_),
    .Q(\int2[6] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1241_ (.RESET_B(net125),
    .D(net276),
    .Q(\int2[7] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1242_ (.RESET_B(net118),
    .D(net296),
    .Q(\int2[8] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1243_ (.RESET_B(net118),
    .D(net266),
    .Q(\int2[9] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1244_ (.RESET_B(net115),
    .D(_0023_),
    .Q(\int2[10] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1245_ (.RESET_B(net115),
    .D(net287),
    .Q(\int2[11] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1246_ (.RESET_B(net114),
    .D(_0025_),
    .Q(\int2[12] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _1247_ (.RESET_B(net114),
    .D(_0026_),
    .Q(\int2[13] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1248_ (.RESET_B(net114),
    .D(net278),
    .Q(\int2[14] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1249_ (.RESET_B(net114),
    .D(net257),
    .Q(\int2[15] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1250_ (.RESET_B(net131),
    .D(net77),
    .Q(uo_out[0]),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1251_ (.RESET_B(net131),
    .D(_0135_),
    .Q(uo_out[1]),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1252_ (.RESET_B(net131),
    .D(net49),
    .Q(uo_out[2]),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1253_ (.RESET_B(net122),
    .D(net51),
    .Q(uo_out[3]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1254_ (.RESET_B(net122),
    .D(net64),
    .Q(uo_out[4]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1255_ (.RESET_B(net124),
    .D(net215),
    .Q(uo_out[5]),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1256_ (.RESET_B(net122),
    .D(net81),
    .Q(uo_out[6]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1257_ (.RESET_B(net122),
    .D(net192),
    .Q(uo_out[7]),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1258_ (.RESET_B(net129),
    .D(_0038_),
    .Q(\int3[0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1259_ (.RESET_B(net129),
    .D(_0045_),
    .Q(\int3[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1260_ (.RESET_B(net130),
    .D(net283),
    .Q(\int3[2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1261_ (.RESET_B(net128),
    .D(net289),
    .Q(\int3[3] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1262_ (.RESET_B(net126),
    .D(_0048_),
    .Q(\int3[4] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1263_ (.RESET_B(net126),
    .D(net270),
    .Q(\int3[5] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1264_ (.RESET_B(net125),
    .D(net304),
    .Q(\int3[6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1265_ (.RESET_B(net125),
    .D(net293),
    .Q(\int3[7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1266_ (.RESET_B(net118),
    .D(net311),
    .Q(\int3[8] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1267_ (.RESET_B(net118),
    .D(net299),
    .Q(\int3[9] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1268_ (.RESET_B(net118),
    .D(net307),
    .Q(\int3[10] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1269_ (.RESET_B(net115),
    .D(net301),
    .Q(\int3[11] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1270_ (.RESET_B(net116),
    .D(net309),
    .Q(\int3[12] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _1271_ (.RESET_B(net116),
    .D(net273),
    .Q(\int3[13] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _1272_ (.RESET_B(net116),
    .D(net280),
    .Q(\int3[14] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1273_ (.RESET_B(net116),
    .D(net259),
    .Q(\int3[15] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_tielo tt_um_cic_filter_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_cic_filter_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_cic_filter_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_cic_filter_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_cic_filter_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_cic_filter_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_cic_filter_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_cic_filter_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_cic_filter_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_cic_filter_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_cic_filter_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_cic_filter_demo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_cic_filter_demo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_cic_filter_demo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_cic_filter_demo_17 (.L_LO(net17));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 fanout94 (.A(net102),
    .X(net94));
 sg13g2_buf_8 fanout95 (.A(net97),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(net102),
    .X(net97));
 sg13g2_buf_8 fanout98 (.A(net101),
    .X(net98));
 sg13g2_buf_8 fanout99 (.A(net101),
    .X(net99));
 sg13g2_buf_8 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_8 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_8 fanout102 (.A(sample_en),
    .X(net102));
 sg13g2_buf_8 fanout103 (.A(net105),
    .X(net103));
 sg13g2_buf_8 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net108),
    .X(net105));
 sg13g2_buf_8 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_8 fanout107 (.A(net108),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(sample_en),
    .X(net108));
 sg13g2_buf_8 fanout109 (.A(net113),
    .X(net109));
 sg13g2_buf_8 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_8 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_8 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(sample_en),
    .X(net113));
 sg13g2_buf_8 fanout114 (.A(net117),
    .X(net114));
 sg13g2_buf_8 fanout115 (.A(net117),
    .X(net115));
 sg13g2_buf_8 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_8 fanout117 (.A(net119),
    .X(net117));
 sg13g2_buf_8 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(rst_n),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net124),
    .X(net121));
 sg13g2_buf_8 fanout122 (.A(net124),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(rst_n),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net127),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(net137),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(net130),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(net137),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(net136),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(rst_n),
    .X(net137));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_cic_filter_demo_2 (.L_LO(net2));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\count[0] ),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold2 (.A(\count[4] ),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0004_),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold4 (.A(\count[3] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0003_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold6 (.A(\count[2] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0151_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold8 (.A(\count[1] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold9 (.A(\int2[0] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0022_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold11 (.A(\int3[0] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold12 (.A(\int1[10] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0007_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold14 (.A(\int1[15] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0012_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold16 (.A(\int1[2] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0014_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold18 (.A(\int1[9] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0021_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold20 (.A(\int1[6] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0018_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold22 (.A(\int1[11] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold23 (.A(\int1[0] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold24 (.A(\int1[12] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold25 (.A(\int1[5] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0017_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold27 (.A(\int1[7] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0019_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold29 (.A(\int1[3] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0015_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold31 (.A(uo_out[2]),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0136_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold33 (.A(uo_out[3]),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0137_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold35 (.A(\int1[13] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold36 (.A(\comb3_d[4] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0296_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0090_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold39 (.A(\comb2[4] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0421_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0122_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold42 (.A(\comb3_d[0] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0086_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold44 (.A(\comb1[5] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0107_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold46 (.A(uo_out[4]),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0138_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold48 (.A(\comb2_d[7] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0077_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold50 (.A(\comb3_d[1] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0087_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold52 (.A(\comb1_d[4] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0058_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold54 (.A(\comb1[12] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0368_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0114_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold57 (.A(\comb3_d[9] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0095_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold59 (.A(uo_out[0]),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0134_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold61 (.A(\comb2[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0121_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold63 (.A(uo_out[6]),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0140_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold65 (.A(\comb2_d[5] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold66 (.A(\comb2[10] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0128_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold68 (.A(\comb3_d[6] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0092_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold70 (.A(\comb3_d[15] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0101_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold72 (.A(\comb2_d[15] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0085_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold74 (.A(\comb1_d[15] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0069_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold76 (.A(\comb2_d[9] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0079_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold78 (.A(\comb2[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0120_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold80 (.A(\comb2[15] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0133_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold82 (.A(\comb3_d[7] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0093_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold84 (.A(\comb2[6] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0124_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold86 (.A(\comb1_d[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0055_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold88 (.A(\comb2_d[13] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0083_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold90 (.A(\comb1_d[9] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0063_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold92 (.A(\comb1[10] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0112_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold94 (.A(\comb1[14] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0116_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold96 (.A(\comb2[12] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0466_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0130_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold99 (.A(\comb3_d[13] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0099_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold101 (.A(\comb1_d[14] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0068_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold103 (.A(\comb3_d[5] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0091_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold105 (.A(\comb1_d[13] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0067_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold107 (.A(\comb1[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0308_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0104_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold110 (.A(\comb1[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0299_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0103_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold113 (.A(\comb2[1] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0119_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold115 (.A(\comb1_d[5] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0059_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold117 (.A(\comb3_d[2] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold118 (.A(\comb3_d[11] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0097_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold120 (.A(\comb2_d[14] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold121 (.A(\comb3_d[10] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold122 (.A(\comb2[14] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0132_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold124 (.A(\comb2[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0118_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold126 (.A(\comb1_d[7] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0061_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold128 (.A(\comb2[8] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0126_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold130 (.A(uo_out[7]),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0141_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold132 (.A(\comb1[15] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0117_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold134 (.A(\comb1[4] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0106_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold136 (.A(\comb3_d[8] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold137 (.A(\comb1[6] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0108_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold139 (.A(\comb2_d[8] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0078_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold141 (.A(\comb2_d[10] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold142 (.A(\comb2_d[12] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold143 (.A(\comb1_d[2] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0056_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold145 (.A(\comb2[9] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0127_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold147 (.A(\comb2_d[0] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0070_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold149 (.A(\comb3_d[14] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold150 (.A(\comb1[3] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0309_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0105_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold153 (.A(uo_out[5]),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0139_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold155 (.A(\comb1[13] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0115_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold157 (.A(\comb2_d[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold158 (.A(\comb2_d[6] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold159 (.A(\comb2[13] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0131_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold161 (.A(\comb2_d[1] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold162 (.A(\comb1_d[10] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0064_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold164 (.A(\comb1_d[8] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0062_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold166 (.A(\comb1_d[3] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0057_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold168 (.A(uo_out[1]),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold169 (.A(\comb2[7] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0125_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold171 (.A(\comb1_d[6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0060_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold173 (.A(\comb2_d[4] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold174 (.A(\comb1_d[0] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold175 (.A(\comb1[8] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0339_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0110_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold178 (.A(\comb2[5] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold179 (.A(\comb3_d[12] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold180 (.A(\comb1_d[12] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0066_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold182 (.A(\comb2[11] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0129_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold184 (.A(\comb1[7] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0109_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold186 (.A(\comb1[0] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold187 (.A(\comb1_d[11] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0065_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold189 (.A(\comb3_d[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold190 (.A(\comb2_d[3] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold191 (.A(\comb2_d[11] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0081_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold193 (.A(\comb1[9] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold194 (.A(\comb1[11] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold195 (.A(\int2[15] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0028_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold197 (.A(\int3[15] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0044_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold199 (.A(\int1[1] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0157_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold201 (.A(\int3[1] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0222_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold203 (.A(\int1[8] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0189_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0037_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold206 (.A(\int1[14] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold207 (.A(\int2[4] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0234_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0049_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold210 (.A(\int2[12] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0270_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0042_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold213 (.A(\int1[3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold214 (.A(\int2[6] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0035_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold216 (.A(\int2[14] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0027_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold218 (.A(\int3[14] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0043_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold220 (.A(\int2[2] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0224_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0046_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold223 (.A(\int1[4] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold224 (.A(\int2[3] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold225 (.A(\int2[11] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0024_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold227 (.A(\int3[3] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0047_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold229 (.A(\int2[5] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold230 (.A(\int3[7] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0243_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0051_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold233 (.A(\int2[13] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold234 (.A(\int2[8] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0036_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold236 (.A(\int2[9] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0251_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0053_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold239 (.A(\int3[11] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0040_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold241 (.A(\int2[1] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold242 (.A(\int3[6] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0050_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold244 (.A(\int2[10] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0254_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0039_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold247 (.A(\int3[12] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0041_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold249 (.A(\int3[8] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0052_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold251 (.A(\int3[4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold252 (.A(\int1[11] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold253 (.A(\int3[11] ),
    .X(net314));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_84 ();
 sg13g2_fill_1 FILLER_7_86 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_132 ();
 sg13g2_decap_8 FILLER_7_139 ();
 sg13g2_decap_8 FILLER_7_146 ();
 sg13g2_fill_1 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_fill_2 FILLER_7_166 ();
 sg13g2_decap_8 FILLER_7_171 ();
 sg13g2_decap_8 FILLER_7_178 ();
 sg13g2_decap_4 FILLER_7_185 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_decap_8 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_4 FILLER_7_304 ();
 sg13g2_fill_2 FILLER_7_308 ();
 sg13g2_fill_2 FILLER_7_346 ();
 sg13g2_fill_1 FILLER_7_348 ();
 sg13g2_fill_1 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_57 ();
 sg13g2_decap_8 FILLER_8_64 ();
 sg13g2_decap_8 FILLER_8_71 ();
 sg13g2_decap_4 FILLER_8_78 ();
 sg13g2_decap_8 FILLER_8_104 ();
 sg13g2_decap_4 FILLER_8_111 ();
 sg13g2_fill_1 FILLER_8_115 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_decap_4 FILLER_8_178 ();
 sg13g2_fill_2 FILLER_8_182 ();
 sg13g2_decap_4 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_decap_4 FILLER_8_254 ();
 sg13g2_fill_1 FILLER_8_258 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_4 FILLER_8_281 ();
 sg13g2_fill_1 FILLER_8_285 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_fill_2 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_fill_2 FILLER_9_53 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_fill_2 FILLER_9_61 ();
 sg13g2_fill_1 FILLER_9_73 ();
 sg13g2_fill_1 FILLER_9_164 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_239 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_4 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_29 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_fill_1 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_52 ();
 sg13g2_fill_1 FILLER_10_58 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_decap_4 FILLER_10_244 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_304 ();
 sg13g2_fill_2 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_75 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_367 ();
 sg13g2_fill_1 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_fill_2 FILLER_12_90 ();
 sg13g2_fill_2 FILLER_12_114 ();
 sg13g2_fill_1 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_2 FILLER_12_170 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_decap_4 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_281 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_185 ();
 sg13g2_decap_8 FILLER_13_192 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_fill_2 FILLER_13_228 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_decap_4 FILLER_13_300 ();
 sg13g2_fill_2 FILLER_13_375 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_22 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_decap_4 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_372 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_54 ();
 sg13g2_fill_2 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_89 ();
 sg13g2_fill_2 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_4 FILLER_15_287 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_15_399 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_40 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_2 FILLER_16_82 ();
 sg13g2_fill_1 FILLER_16_134 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_4 FILLER_16_293 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_decap_4 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_fill_1 FILLER_17_83 ();
 sg13g2_fill_1 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_decap_4 FILLER_17_181 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_decap_4 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_1 FILLER_18_45 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_decap_4 FILLER_18_117 ();
 sg13g2_decap_8 FILLER_18_170 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_decap_4 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_304 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_decap_8 FILLER_19_44 ();
 sg13g2_decap_4 FILLER_19_51 ();
 sg13g2_decap_8 FILLER_19_97 ();
 sg13g2_fill_2 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_106 ();
 sg13g2_decap_4 FILLER_19_120 ();
 sg13g2_decap_4 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_177 ();
 sg13g2_decap_8 FILLER_19_184 ();
 sg13g2_decap_4 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_decap_4 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_370 ();
 sg13g2_fill_2 FILLER_19_391 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_decap_8 FILLER_20_93 ();
 sg13g2_fill_2 FILLER_20_100 ();
 sg13g2_decap_4 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_142 ();
 sg13g2_decap_4 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_decap_4 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_9 ();
 sg13g2_fill_1 FILLER_21_29 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_87 ();
 sg13g2_decap_8 FILLER_21_94 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_fill_2 FILLER_21_191 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_decap_4 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_9 ();
 sg13g2_decap_4 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_54 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_decap_8 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_4 FILLER_22_196 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_decap_8 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_4 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_94 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_202 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_71 ();
 sg13g2_fill_1 FILLER_25_82 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_decap_4 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_303 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_359 ();
 sg13g2_decap_4 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_decap_4 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_123 ();
 sg13g2_decap_4 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_34 ();
 sg13g2_decap_4 FILLER_29_40 ();
 sg13g2_fill_1 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_decap_4 FILLER_29_118 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_decap_4 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_381 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_decap_4 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_31_44 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_decap_4 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_decap_4 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_9 ();
 sg13g2_fill_1 FILLER_32_13 ();
 sg13g2_fill_2 FILLER_32_24 ();
 sg13g2_fill_1 FILLER_32_26 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_decap_4 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_decap_4 FILLER_32_297 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_2 FILLER_32_367 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_38 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_decap_4 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_243 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_fill_2 FILLER_34_57 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_52 ();
 sg13g2_fill_2 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_2 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_58 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_decap_4 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_2 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_201 ();
 sg13g2_fill_2 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_379 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_18 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_97 ();
 sg13g2_fill_1 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_380 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule
